// Reading file 'cantest.asc'..

module chip (input io_13_31_1, output io_4_31_0, input io_16_0_0, input io_19_0_1, output io_19_31_1);

reg n1 = 0;
// (0, 0, 'glb_netwk_0')
// (1, 2, 'lutff_global/s_r')
// (1, 3, 'lutff_global/s_r')
// (1, 6, 'lutff_global/s_r')
// (1, 8, 'lutff_global/s_r')
// (1, 9, 'lutff_global/s_r')
// (1, 10, 'lutff_global/s_r')
// (1, 11, 'lutff_global/s_r')
// (1, 12, 'lutff_global/s_r')
// (1, 13, 'lutff_global/s_r')
// (1, 14, 'lutff_global/s_r')
// (1, 15, 'lutff_global/s_r')
// (1, 16, 'lutff_global/s_r')
// (1, 17, 'lutff_global/s_r')
// (1, 19, 'lutff_global/s_r')
// (1, 20, 'lutff_global/s_r')
// (1, 21, 'lutff_global/s_r')
// (2, 1, 'lutff_global/s_r')
// (2, 2, 'lutff_global/s_r')
// (2, 3, 'lutff_global/s_r')
// (2, 6, 'lutff_global/s_r')
// (2, 7, 'lutff_global/s_r')
// (2, 8, 'lutff_global/s_r')
// (2, 9, 'lutff_global/s_r')
// (2, 10, 'lutff_global/s_r')
// (2, 11, 'lutff_global/s_r')
// (2, 12, 'lutff_global/s_r')
// (2, 13, 'lutff_global/s_r')
// (2, 14, 'lutff_global/s_r')
// (2, 15, 'lutff_global/s_r')
// (2, 16, 'lutff_global/s_r')
// (2, 17, 'lutff_global/s_r')
// (2, 18, 'lutff_global/s_r')
// (2, 19, 'lutff_global/s_r')
// (2, 20, 'lutff_global/s_r')
// (2, 21, 'lutff_global/s_r')
// (3, 1, 'lutff_global/s_r')
// (3, 2, 'lutff_global/s_r')
// (3, 3, 'lutff_global/s_r')
// (3, 4, 'lutff_global/s_r')
// (3, 5, 'lutff_global/s_r')
// (3, 6, 'lutff_global/s_r')
// (3, 7, 'lutff_global/s_r')
// (3, 8, 'lutff_global/s_r')
// (3, 9, 'lutff_global/s_r')
// (3, 10, 'lutff_global/s_r')
// (3, 11, 'lutff_global/s_r')
// (3, 12, 'lutff_global/s_r')
// (3, 14, 'lutff_global/s_r')
// (3, 15, 'lutff_global/s_r')
// (3, 16, 'lutff_global/s_r')
// (3, 17, 'lutff_global/s_r')
// (3, 18, 'lutff_global/s_r')
// (3, 20, 'lutff_global/s_r')
// (3, 21, 'lutff_global/s_r')
// (4, 1, 'lutff_global/s_r')
// (4, 2, 'lutff_global/s_r')
// (4, 3, 'lutff_global/s_r')
// (4, 4, 'lutff_global/s_r')
// (4, 5, 'lutff_global/s_r')
// (4, 6, 'lutff_global/s_r')
// (4, 7, 'lutff_global/s_r')
// (4, 10, 'lutff_global/s_r')
// (4, 11, 'lutff_global/s_r')
// (4, 12, 'lutff_global/s_r')
// (4, 14, 'lutff_global/s_r')
// (4, 15, 'lutff_global/s_r')
// (4, 16, 'lutff_global/s_r')
// (4, 17, 'lutff_global/s_r')
// (4, 20, 'lutff_global/s_r')
// (5, 1, 'lutff_global/s_r')
// (5, 2, 'lutff_global/s_r')
// (5, 3, 'lutff_global/s_r')
// (5, 4, 'lutff_global/s_r')
// (5, 5, 'lutff_global/s_r')
// (5, 7, 'lutff_global/s_r')
// (5, 11, 'lutff_global/s_r')
// (5, 14, 'lutff_global/s_r')
// (5, 15, 'lutff_global/s_r')
// (5, 16, 'lutff_global/s_r')
// (5, 17, 'lutff_global/s_r')
// (5, 18, 'lutff_global/s_r')
// (5, 19, 'lutff_global/s_r')
// (5, 20, 'lutff_global/s_r')
// (7, 1, 'lutff_global/s_r')
// (7, 2, 'lutff_global/s_r')
// (7, 3, 'lutff_global/s_r')
// (7, 4, 'lutff_global/s_r')
// (7, 8, 'lutff_global/s_r')
// (7, 9, 'lutff_global/s_r')
// (7, 12, 'lutff_global/s_r')
// (7, 14, 'lutff_global/s_r')
// (7, 17, 'lutff_global/s_r')
// (7, 21, 'lutff_global/s_r')
// (8, 1, 'lutff_global/s_r')
// (8, 2, 'lutff_global/s_r')
// (8, 3, 'lutff_global/s_r')
// (8, 4, 'lutff_global/s_r')
// (8, 5, 'lutff_global/s_r')
// (8, 8, 'lutff_global/s_r')
// (8, 9, 'lutff_global/s_r')
// (8, 12, 'lutff_global/s_r')
// (8, 13, 'lutff_global/s_r')
// (8, 14, 'lutff_global/s_r')
// (8, 20, 'lutff_global/s_r')
// (8, 21, 'lutff_global/s_r')
// (9, 1, 'lutff_global/s_r')
// (9, 3, 'lutff_global/s_r')
// (9, 4, 'lutff_global/s_r')
// (9, 5, 'lutff_global/s_r')
// (9, 7, 'lutff_global/s_r')
// (9, 12, 'lutff_global/s_r')
// (9, 14, 'lutff_global/s_r')
// (9, 21, 'lutff_global/s_r')
// (10, 1, 'lutff_global/s_r')
// (10, 2, 'lutff_global/s_r')
// (10, 3, 'lutff_global/s_r')
// (10, 4, 'lutff_global/s_r')
// (10, 5, 'lutff_global/s_r')
// (10, 12, 'lutff_global/s_r')
// (10, 17, 'lutff_global/s_r')
// (10, 19, 'lutff_global/s_r')
// (10, 20, 'lutff_global/s_r')
// (10, 21, 'lutff_global/s_r')
// (11, 2, 'lutff_global/s_r')
// (11, 3, 'lutff_global/s_r')
// (11, 4, 'lutff_global/s_r')
// (11, 5, 'lutff_global/s_r')
// (11, 6, 'lutff_global/s_r')
// (11, 12, 'lutff_global/s_r')
// (11, 13, 'lutff_global/s_r')
// (11, 14, 'lutff_global/s_r')
// (11, 15, 'lutff_global/s_r')
// (11, 17, 'lutff_global/s_r')
// (11, 19, 'lutff_global/s_r')
// (11, 20, 'lutff_global/s_r')
// (11, 21, 'lutff_global/s_r')
// (11, 30, 'lutff_global/s_r')
// (12, 5, 'lutff_global/s_r')
// (12, 7, 'lutff_global/s_r')
// (12, 8, 'lutff_global/s_r')
// (12, 9, 'lutff_global/s_r')
// (12, 10, 'lutff_global/s_r')
// (12, 11, 'lutff_global/s_r')
// (12, 14, 'lutff_global/s_r')
// (12, 15, 'lutff_global/s_r')
// (12, 17, 'lutff_global/s_r')
// (12, 18, 'lutff_global/s_r')
// (12, 19, 'lutff_global/s_r')
// (12, 20, 'lutff_global/s_r')
// (12, 21, 'lutff_global/s_r')
// (12, 22, 'lutff_global/s_r')
// (12, 23, 'lutff_global/s_r')
// (13, 0, 'fabout')
// (13, 0, 'local_g1_0')
// (13, 0, 'span12_vert_8')
// (13, 1, 'sp12_v_b_8')
// (13, 2, 'lutff_global/s_r')
// (13, 2, 'sp12_v_b_7')
// (13, 3, 'sp12_v_b_4')
// (13, 4, 'lutff_global/s_r')
// (13, 4, 'sp12_v_b_3')
// (13, 5, 'lutff_global/s_r')
// (13, 5, 'sp12_h_r_0')
// (13, 5, 'sp12_v_b_0')
// (13, 6, 'lutff_global/s_r')
// (13, 8, 'lutff_global/s_r')
// (13, 9, 'lutff_global/s_r')
// (13, 10, 'lutff_global/s_r')
// (13, 11, 'lutff_global/s_r')
// (13, 12, 'lutff_global/s_r')
// (13, 14, 'lutff_global/s_r')
// (13, 18, 'lutff_global/s_r')
// (13, 19, 'lutff_global/s_r')
// (13, 21, 'lutff_global/s_r')
// (13, 22, 'lutff_global/s_r')
// (13, 23, 'lutff_global/s_r')
// (14, 1, 'lutff_global/s_r')
// (14, 2, 'lutff_global/s_r')
// (14, 3, 'lutff_global/s_r')
// (14, 4, 'lutff_global/s_r')
// (14, 5, 'lutff_global/s_r')
// (14, 5, 'sp12_h_r_3')
// (14, 6, 'lutff_global/s_r')
// (14, 7, 'lutff_global/s_r')
// (14, 10, 'lutff_global/s_r')
// (14, 11, 'lutff_global/s_r')
// (14, 13, 'lutff_global/s_r')
// (14, 13, 'sp4_r_v_b_44')
// (14, 14, 'sp4_r_v_b_33')
// (14, 15, 'local_g3_4')
// (14, 15, 'lutff_4/in_1')
// (14, 15, 'sp4_r_v_b_20')
// (14, 16, 'lutff_global/s_r')
// (14, 16, 'sp4_r_v_b_9')
// (14, 18, 'lutff_global/s_r')
// (14, 19, 'lutff_global/s_r')
// (14, 21, 'lutff_global/s_r')
// (15, 2, 'lutff_global/s_r')
// (15, 3, 'lutff_global/s_r')
// (15, 4, 'lutff_global/s_r')
// (15, 5, 'lutff_global/s_r')
// (15, 5, 'sp12_h_r_4')
// (15, 12, 'lutff_global/s_r')
// (15, 12, 'sp4_h_r_9')
// (15, 12, 'sp4_r_v_b_47')
// (15, 12, 'sp4_v_t_44')
// (15, 13, 'lutff_global/s_r')
// (15, 13, 'sp4_r_v_b_34')
// (15, 13, 'sp4_v_b_44')
// (15, 14, 'sp4_r_v_b_23')
// (15, 14, 'sp4_v_b_33')
// (15, 15, 'lutff_global/s_r')
// (15, 15, 'sp4_r_v_b_10')
// (15, 15, 'sp4_v_b_20')
// (15, 16, 'lutff_global/s_r')
// (15, 16, 'sp4_h_r_8')
// (15, 16, 'sp4_v_b_9')
// (15, 17, 'lutff_global/s_r')
// (15, 20, 'lutff_global/s_r')
// (15, 21, 'lutff_global/s_r')
// (16, 1, 'lutff_global/s_r')
// (16, 2, 'lutff_global/s_r')
// (16, 3, 'lutff_global/s_r')
// (16, 5, 'lutff_global/s_r')
// (16, 5, 'sp12_h_r_7')
// (16, 6, 'lutff_global/s_r')
// (16, 11, 'sp4_h_r_10')
// (16, 11, 'sp4_v_t_47')
// (16, 12, 'sp4_h_r_20')
// (16, 12, 'sp4_v_b_47')
// (16, 13, 'lutff_global/s_r')
// (16, 13, 'sp4_v_b_34')
// (16, 14, 'local_g1_7')
// (16, 14, 'lutff_1/in_1')
// (16, 14, 'sp4_v_b_23')
// (16, 15, 'sp4_h_r_8')
// (16, 15, 'sp4_v_b_10')
// (16, 16, 'local_g0_5')
// (16, 16, 'lutff_1/in_0')
// (16, 16, 'lutff_3/in_2')
// (16, 16, 'sp4_h_r_21')
// (16, 17, 'lutff_global/s_r')
// (16, 18, 'lutff_global/s_r')
// (16, 19, 'lutff_global/s_r')
// (17, 5, 'sp12_h_r_8')
// (17, 11, 'lutff_global/s_r')
// (17, 11, 'sp4_h_r_23')
// (17, 12, 'sp4_h_r_33')
// (17, 13, 'lutff_global/s_r')
// (17, 14, 'lutff_global/s_r')
// (17, 15, 'local_g0_5')
// (17, 15, 'lutff_2/in_3')
// (17, 15, 'lutff_7/in_2')
// (17, 15, 'sp4_h_r_21')
// (17, 16, 'sp4_h_r_32')
// (17, 18, 'lutff_global/s_r')
// (17, 20, 'lutff_global/s_r')
// (18, 5, 'sp12_h_r_11')
// (18, 6, 'lutff_global/s_r')
// (18, 11, 'sp4_h_r_34')
// (18, 12, 'sp4_h_r_44')
// (18, 12, 'sp4_r_v_b_36')
// (18, 13, 'sp4_r_v_b_25')
// (18, 13, 'sp4_r_v_b_38')
// (18, 14, 'local_g2_4')
// (18, 14, 'lutff_0/in_2')
// (18, 14, 'lutff_3/in_3')
// (18, 14, 'sp4_r_v_b_12')
// (18, 14, 'sp4_r_v_b_27')
// (18, 15, 'sp4_h_r_32')
// (18, 15, 'sp4_r_v_b_1')
// (18, 15, 'sp4_r_v_b_14')
// (18, 16, 'sp4_h_r_45')
// (18, 16, 'sp4_r_v_b_3')
// (19, 5, 'sp12_h_r_12')
// (19, 6, 'sp4_h_r_1')
// (19, 8, 'sp4_h_r_2')
// (19, 8, 'sp4_r_v_b_40')
// (19, 9, 'sp4_r_v_b_29')
// (19, 10, 'sp4_r_v_b_16')
// (19, 11, 'sp4_h_r_47')
// (19, 11, 'sp4_h_r_7')
// (19, 11, 'sp4_r_v_b_5')
// (19, 11, 'sp4_v_t_36')
// (19, 12, 'sp4_h_l_44')
// (19, 12, 'sp4_h_r_9')
// (19, 12, 'sp4_r_v_b_45')
// (19, 12, 'sp4_v_b_36')
// (19, 12, 'sp4_v_t_38')
// (19, 13, 'sp4_r_v_b_32')
// (19, 13, 'sp4_v_b_25')
// (19, 13, 'sp4_v_b_38')
// (19, 14, 'sp4_r_v_b_21')
// (19, 14, 'sp4_v_b_12')
// (19, 14, 'sp4_v_b_27')
// (19, 15, 'sp4_h_r_45')
// (19, 15, 'sp4_r_v_b_8')
// (19, 15, 'sp4_v_b_1')
// (19, 15, 'sp4_v_b_14')
// (19, 16, 'sp4_h_l_45')
// (19, 16, 'sp4_v_b_3')
// (20, 4, 'lutff_global/s_r')
// (20, 5, 'sp12_h_r_15')
// (20, 6, 'local_g0_4')
// (20, 6, 'lutff_7/in_1')
// (20, 6, 'lutff_global/s_r')
// (20, 6, 'sp4_h_r_12')
// (20, 7, 'sp4_h_r_5')
// (20, 7, 'sp4_v_t_40')
// (20, 8, 'local_g1_7')
// (20, 8, 'lutff_5/in_3')
// (20, 8, 'sp4_h_r_15')
// (20, 8, 'sp4_v_b_40')
// (20, 9, 'sp4_v_b_29')
// (20, 10, 'sp4_v_b_16')
// (20, 11, 'sp4_h_l_47')
// (20, 11, 'sp4_h_r_18')
// (20, 11, 'sp4_v_b_5')
// (20, 11, 'sp4_v_t_45')
// (20, 12, 'sp4_h_r_20')
// (20, 12, 'sp4_v_b_45')
// (20, 13, 'sp4_v_b_32')
// (20, 14, 'sp4_v_b_21')
// (20, 15, 'sp4_h_l_45')
// (20, 15, 'sp4_v_b_8')
// (21, 5, 'sp12_h_r_16')
// (21, 6, 'sp4_h_r_25')
// (21, 7, 'lutff_global/s_r')
// (21, 7, 'sp4_h_r_16')
// (21, 8, 'lutff_global/s_r')
// (21, 8, 'sp4_h_r_26')
// (21, 11, 'sp4_h_r_31')
// (21, 12, 'sp4_h_r_33')
// (22, 3, 'sp4_r_v_b_36')
// (22, 4, 'neigh_op_tnr_6')
// (22, 4, 'sp4_r_v_b_25')
// (22, 4, 'sp4_r_v_b_41')
// (22, 5, 'neigh_op_rgt_6')
// (22, 5, 'sp12_h_r_19')
// (22, 5, 'sp4_r_v_b_12')
// (22, 5, 'sp4_r_v_b_28')
// (22, 5, 'sp4_r_v_b_44')
// (22, 6, 'neigh_op_bnr_6')
// (22, 6, 'sp4_h_r_36')
// (22, 6, 'sp4_r_v_b_1')
// (22, 6, 'sp4_r_v_b_17')
// (22, 6, 'sp4_r_v_b_33')
// (22, 7, 'local_g1_4')
// (22, 7, 'lutff_5/in_2')
// (22, 7, 'lutff_global/s_r')
// (22, 7, 'sp4_h_r_29')
// (22, 7, 'sp4_r_v_b_20')
// (22, 7, 'sp4_r_v_b_4')
// (22, 8, 'local_g2_1')
// (22, 8, 'lutff_1/in_2')
// (22, 8, 'lutff_2/in_1')
// (22, 8, 'lutff_6/in_1')
// (22, 8, 'sp4_h_r_39')
// (22, 8, 'sp4_r_v_b_42')
// (22, 8, 'sp4_r_v_b_9')
// (22, 9, 'sp4_r_v_b_31')
// (22, 9, 'sp4_r_v_b_44')
// (22, 10, 'sp4_r_v_b_18')
// (22, 10, 'sp4_r_v_b_33')
// (22, 11, 'sp4_h_r_42')
// (22, 11, 'sp4_r_v_b_20')
// (22, 11, 'sp4_r_v_b_7')
// (22, 12, 'sp4_h_r_44')
// (22, 12, 'sp4_r_v_b_9')
// (23, 2, 'sp4_v_t_36')
// (23, 3, 'sp4_v_b_36')
// (23, 3, 'sp4_v_t_41')
// (23, 4, 'neigh_op_top_6')
// (23, 4, 'sp4_r_v_b_40')
// (23, 4, 'sp4_v_b_25')
// (23, 4, 'sp4_v_b_41')
// (23, 4, 'sp4_v_t_44')
// (23, 5, 'lutff_6/out')
// (23, 5, 'sp12_h_r_20')
// (23, 5, 'sp4_r_v_b_29')
// (23, 5, 'sp4_v_b_12')
// (23, 5, 'sp4_v_b_28')
// (23, 5, 'sp4_v_b_44')
// (23, 6, 'neigh_op_bot_6')
// (23, 6, 'sp4_h_l_36')
// (23, 6, 'sp4_r_v_b_16')
// (23, 6, 'sp4_v_b_1')
// (23, 6, 'sp4_v_b_17')
// (23, 6, 'sp4_v_b_33')
// (23, 7, 'local_g1_5')
// (23, 7, 'lutff_2/in_2')
// (23, 7, 'lutff_global/s_r')
// (23, 7, 'sp4_h_r_40')
// (23, 7, 'sp4_r_v_b_5')
// (23, 7, 'sp4_v_b_20')
// (23, 7, 'sp4_v_b_4')
// (23, 7, 'sp4_v_t_42')
// (23, 8, 'sp4_h_l_39')
// (23, 8, 'sp4_v_b_42')
// (23, 8, 'sp4_v_b_9')
// (23, 8, 'sp4_v_t_44')
// (23, 9, 'sp4_v_b_31')
// (23, 9, 'sp4_v_b_44')
// (23, 10, 'sp4_v_b_18')
// (23, 10, 'sp4_v_b_33')
// (23, 11, 'sp4_h_l_42')
// (23, 11, 'sp4_v_b_20')
// (23, 11, 'sp4_v_b_7')
// (23, 12, 'sp4_h_l_44')
// (23, 12, 'sp4_v_b_9')
// (24, 3, 'sp4_v_t_40')
// (24, 4, 'neigh_op_tnl_6')
// (24, 4, 'sp4_v_b_40')
// (24, 5, 'neigh_op_lft_6')
// (24, 5, 'sp12_h_r_23')
// (24, 5, 'sp4_v_b_29')
// (24, 6, 'neigh_op_bnl_6')
// (24, 6, 'sp4_v_b_16')
// (24, 7, 'sp4_h_l_40')
// (24, 7, 'sp4_v_b_5')
// (25, 5, 'sp12_h_l_23')

wire io_13_31_1;
// (0, 0, 'glb_netwk_1')
// (1, 2, 'lutff_global/clk')
// (1, 3, 'lutff_global/clk')
// (1, 4, 'lutff_global/clk')
// (1, 5, 'lutff_global/clk')
// (1, 6, 'lutff_global/clk')
// (1, 8, 'lutff_global/clk')
// (1, 9, 'lutff_global/clk')
// (1, 10, 'lutff_global/clk')
// (1, 11, 'lutff_global/clk')
// (1, 12, 'lutff_global/clk')
// (1, 13, 'lutff_global/clk')
// (1, 14, 'lutff_global/clk')
// (1, 15, 'lutff_global/clk')
// (1, 16, 'lutff_global/clk')
// (1, 17, 'lutff_global/clk')
// (1, 19, 'lutff_global/clk')
// (1, 20, 'lutff_global/clk')
// (1, 21, 'lutff_global/clk')
// (2, 1, 'lutff_global/clk')
// (2, 2, 'lutff_global/clk')
// (2, 3, 'lutff_global/clk')
// (2, 4, 'lutff_global/clk')
// (2, 5, 'lutff_global/clk')
// (2, 6, 'lutff_global/clk')
// (2, 7, 'lutff_global/clk')
// (2, 8, 'lutff_global/clk')
// (2, 9, 'lutff_global/clk')
// (2, 10, 'lutff_global/clk')
// (2, 11, 'lutff_global/clk')
// (2, 12, 'lutff_global/clk')
// (2, 13, 'lutff_global/clk')
// (2, 14, 'lutff_global/clk')
// (2, 15, 'lutff_global/clk')
// (2, 16, 'lutff_global/clk')
// (2, 17, 'lutff_global/clk')
// (2, 18, 'lutff_global/clk')
// (2, 19, 'lutff_global/clk')
// (2, 20, 'lutff_global/clk')
// (2, 21, 'lutff_global/clk')
// (3, 1, 'lutff_global/clk')
// (3, 2, 'lutff_global/clk')
// (3, 3, 'lutff_global/clk')
// (3, 4, 'lutff_global/clk')
// (3, 5, 'lutff_global/clk')
// (3, 6, 'lutff_global/clk')
// (3, 7, 'lutff_global/clk')
// (3, 8, 'lutff_global/clk')
// (3, 9, 'lutff_global/clk')
// (3, 10, 'lutff_global/clk')
// (3, 11, 'lutff_global/clk')
// (3, 12, 'lutff_global/clk')
// (3, 14, 'lutff_global/clk')
// (3, 15, 'lutff_global/clk')
// (3, 16, 'lutff_global/clk')
// (3, 17, 'lutff_global/clk')
// (3, 18, 'lutff_global/clk')
// (3, 20, 'lutff_global/clk')
// (3, 21, 'lutff_global/clk')
// (4, 1, 'lutff_global/clk')
// (4, 2, 'lutff_global/clk')
// (4, 3, 'lutff_global/clk')
// (4, 4, 'lutff_global/clk')
// (4, 5, 'lutff_global/clk')
// (4, 6, 'lutff_global/clk')
// (4, 7, 'lutff_global/clk')
// (4, 8, 'lutff_global/clk')
// (4, 9, 'lutff_global/clk')
// (4, 10, 'lutff_global/clk')
// (4, 11, 'lutff_global/clk')
// (4, 12, 'lutff_global/clk')
// (4, 14, 'lutff_global/clk')
// (4, 15, 'lutff_global/clk')
// (4, 16, 'lutff_global/clk')
// (4, 17, 'lutff_global/clk')
// (4, 20, 'lutff_global/clk')
// (5, 1, 'lutff_global/clk')
// (5, 2, 'lutff_global/clk')
// (5, 3, 'lutff_global/clk')
// (5, 4, 'lutff_global/clk')
// (5, 5, 'lutff_global/clk')
// (5, 6, 'lutff_global/clk')
// (5, 7, 'lutff_global/clk')
// (5, 8, 'lutff_global/clk')
// (5, 9, 'lutff_global/clk')
// (5, 10, 'lutff_global/clk')
// (5, 11, 'lutff_global/clk')
// (5, 12, 'lutff_global/clk')
// (5, 13, 'lutff_global/clk')
// (5, 14, 'lutff_global/clk')
// (5, 15, 'lutff_global/clk')
// (5, 16, 'lutff_global/clk')
// (5, 17, 'lutff_global/clk')
// (5, 18, 'lutff_global/clk')
// (5, 19, 'lutff_global/clk')
// (5, 20, 'lutff_global/clk')
// (7, 1, 'lutff_global/clk')
// (7, 2, 'lutff_global/clk')
// (7, 3, 'lutff_global/clk')
// (7, 4, 'lutff_global/clk')
// (7, 5, 'lutff_global/clk')
// (7, 6, 'lutff_global/clk')
// (7, 7, 'lutff_global/clk')
// (7, 8, 'lutff_global/clk')
// (7, 9, 'lutff_global/clk')
// (7, 10, 'lutff_global/clk')
// (7, 11, 'lutff_global/clk')
// (7, 12, 'lutff_global/clk')
// (7, 13, 'lutff_global/clk')
// (7, 14, 'lutff_global/clk')
// (7, 17, 'lutff_global/clk')
// (7, 21, 'lutff_global/clk')
// (8, 1, 'lutff_global/clk')
// (8, 2, 'lutff_global/clk')
// (8, 3, 'lutff_global/clk')
// (8, 4, 'lutff_global/clk')
// (8, 5, 'lutff_global/clk')
// (8, 8, 'lutff_global/clk')
// (8, 9, 'lutff_global/clk')
// (8, 10, 'lutff_global/clk')
// (8, 11, 'lutff_global/clk')
// (8, 12, 'lutff_global/clk')
// (8, 13, 'lutff_global/clk')
// (8, 14, 'lutff_global/clk')
// (8, 20, 'lutff_global/clk')
// (8, 21, 'lutff_global/clk')
// (8, 22, 'lutff_global/clk')
// (9, 1, 'lutff_global/clk')
// (9, 3, 'lutff_global/clk')
// (9, 4, 'lutff_global/clk')
// (9, 5, 'lutff_global/clk')
// (9, 6, 'lutff_global/clk')
// (9, 7, 'lutff_global/clk')
// (9, 8, 'lutff_global/clk')
// (9, 9, 'lutff_global/clk')
// (9, 10, 'lutff_global/clk')
// (9, 11, 'lutff_global/clk')
// (9, 12, 'lutff_global/clk')
// (9, 13, 'lutff_global/clk')
// (9, 14, 'lutff_global/clk')
// (9, 15, 'lutff_global/clk')
// (9, 17, 'lutff_global/clk')
// (9, 21, 'lutff_global/clk')
// (10, 1, 'lutff_global/clk')
// (10, 2, 'lutff_global/clk')
// (10, 3, 'lutff_global/clk')
// (10, 4, 'lutff_global/clk')
// (10, 5, 'lutff_global/clk')
// (10, 6, 'lutff_global/clk')
// (10, 7, 'lutff_global/clk')
// (10, 8, 'lutff_global/clk')
// (10, 9, 'lutff_global/clk')
// (10, 10, 'lutff_global/clk')
// (10, 11, 'lutff_global/clk')
// (10, 12, 'lutff_global/clk')
// (10, 13, 'lutff_global/clk')
// (10, 14, 'lutff_global/clk')
// (10, 15, 'lutff_global/clk')
// (10, 16, 'lutff_global/clk')
// (10, 17, 'lutff_global/clk')
// (10, 19, 'lutff_global/clk')
// (10, 20, 'lutff_global/clk')
// (10, 21, 'lutff_global/clk')
// (11, 2, 'lutff_global/clk')
// (11, 3, 'lutff_global/clk')
// (11, 4, 'lutff_global/clk')
// (11, 5, 'lutff_global/clk')
// (11, 6, 'lutff_global/clk')
// (11, 7, 'lutff_global/clk')
// (11, 8, 'lutff_global/clk')
// (11, 9, 'lutff_global/clk')
// (11, 10, 'lutff_global/clk')
// (11, 11, 'lutff_global/clk')
// (11, 12, 'lutff_global/clk')
// (11, 13, 'lutff_global/clk')
// (11, 14, 'lutff_global/clk')
// (11, 15, 'lutff_global/clk')
// (11, 16, 'lutff_global/clk')
// (11, 17, 'lutff_global/clk')
// (11, 18, 'lutff_global/clk')
// (11, 19, 'lutff_global/clk')
// (11, 20, 'lutff_global/clk')
// (11, 21, 'lutff_global/clk')
// (11, 30, 'lutff_global/clk')
// (12, 5, 'lutff_global/clk')
// (12, 7, 'lutff_global/clk')
// (12, 8, 'lutff_global/clk')
// (12, 9, 'lutff_global/clk')
// (12, 10, 'lutff_global/clk')
// (12, 11, 'lutff_global/clk')
// (12, 12, 'lutff_global/clk')
// (12, 13, 'lutff_global/clk')
// (12, 14, 'lutff_global/clk')
// (12, 15, 'lutff_global/clk')
// (12, 16, 'lutff_global/clk')
// (12, 17, 'lutff_global/clk')
// (12, 18, 'lutff_global/clk')
// (12, 19, 'lutff_global/clk')
// (12, 20, 'lutff_global/clk')
// (12, 21, 'lutff_global/clk')
// (12, 22, 'lutff_global/clk')
// (12, 23, 'lutff_global/clk')
// (12, 30, 'neigh_op_tnr_2')
// (12, 30, 'neigh_op_tnr_6')
// (12, 31, 'span4_horz_r_2')
// (13, 2, 'lutff_global/clk')
// (13, 4, 'lutff_global/clk')
// (13, 5, 'lutff_global/clk')
// (13, 6, 'lutff_global/clk')
// (13, 7, 'lutff_global/clk')
// (13, 8, 'lutff_global/clk')
// (13, 9, 'lutff_global/clk')
// (13, 10, 'lutff_global/clk')
// (13, 11, 'lutff_global/clk')
// (13, 12, 'lutff_global/clk')
// (13, 13, 'lutff_global/clk')
// (13, 14, 'lutff_global/clk')
// (13, 15, 'lutff_global/clk')
// (13, 16, 'lutff_global/clk')
// (13, 18, 'lutff_global/clk')
// (13, 19, 'lutff_global/clk')
// (13, 20, 'lutff_global/clk')
// (13, 21, 'lutff_global/clk')
// (13, 22, 'lutff_global/clk')
// (13, 23, 'lutff_global/clk')
// (13, 30, 'neigh_op_top_2')
// (13, 30, 'neigh_op_top_6')
// (13, 31, 'fabout')
// (13, 31, 'io_1/D_IN_0')
// (13, 31, 'io_1/PAD')
// (13, 31, 'local_g1_6')
// (13, 31, 'span4_horz_r_6')
// (14, 1, 'lutff_global/clk')
// (14, 2, 'lutff_global/clk')
// (14, 3, 'lutff_global/clk')
// (14, 4, 'lutff_global/clk')
// (14, 5, 'lutff_global/clk')
// (14, 6, 'lutff_global/clk')
// (14, 7, 'lutff_global/clk')
// (14, 8, 'lutff_global/clk')
// (14, 9, 'lutff_global/clk')
// (14, 10, 'lutff_global/clk')
// (14, 11, 'lutff_global/clk')
// (14, 13, 'lutff_global/clk')
// (14, 16, 'lutff_global/clk')
// (14, 17, 'lutff_global/clk')
// (14, 18, 'lutff_global/clk')
// (14, 19, 'lutff_global/clk')
// (14, 20, 'lutff_global/clk')
// (14, 21, 'lutff_global/clk')
// (14, 30, 'neigh_op_tnl_2')
// (14, 30, 'neigh_op_tnl_6')
// (14, 31, 'span4_horz_r_10')
// (15, 2, 'lutff_global/clk')
// (15, 3, 'lutff_global/clk')
// (15, 4, 'lutff_global/clk')
// (15, 5, 'lutff_global/clk')
// (15, 6, 'lutff_global/clk')
// (15, 7, 'lutff_global/clk')
// (15, 8, 'lutff_global/clk')
// (15, 9, 'lutff_global/clk')
// (15, 10, 'lutff_global/clk')
// (15, 11, 'lutff_global/clk')
// (15, 12, 'lutff_global/clk')
// (15, 13, 'lutff_global/clk')
// (15, 14, 'lutff_global/clk')
// (15, 15, 'lutff_global/clk')
// (15, 16, 'lutff_global/clk')
// (15, 17, 'lutff_global/clk')
// (15, 19, 'lutff_global/clk')
// (15, 20, 'lutff_global/clk')
// (15, 21, 'lutff_global/clk')
// (15, 22, 'lutff_global/clk')
// (15, 23, 'lutff_global/clk')
// (15, 31, 'span4_horz_r_14')
// (16, 1, 'lutff_global/clk')
// (16, 2, 'lutff_global/clk')
// (16, 3, 'lutff_global/clk')
// (16, 4, 'lutff_global/clk')
// (16, 5, 'lutff_global/clk')
// (16, 6, 'lutff_global/clk')
// (16, 7, 'lutff_global/clk')
// (16, 8, 'lutff_global/clk')
// (16, 9, 'lutff_global/clk')
// (16, 10, 'lutff_global/clk')
// (16, 11, 'lutff_global/clk')
// (16, 12, 'lutff_global/clk')
// (16, 13, 'lutff_global/clk')
// (16, 14, 'lutff_global/clk')
// (16, 15, 'lutff_global/clk')
// (16, 16, 'lutff_global/clk')
// (16, 17, 'lutff_global/clk')
// (16, 18, 'lutff_global/clk')
// (16, 19, 'lutff_global/clk')
// (16, 20, 'lutff_global/clk')
// (16, 21, 'lutff_global/clk')
// (16, 22, 'lutff_global/clk')
// (16, 23, 'lutff_global/clk')
// (16, 24, 'lutff_global/clk')
// (16, 31, 'span4_horz_l_14')
// (17, 1, 'lutff_global/clk')
// (17, 2, 'lutff_global/clk')
// (17, 3, 'lutff_global/clk')
// (17, 4, 'lutff_global/clk')
// (17, 5, 'lutff_global/clk')
// (17, 7, 'lutff_global/clk')
// (17, 8, 'lutff_global/clk')
// (17, 9, 'lutff_global/clk')
// (17, 10, 'lutff_global/clk')
// (17, 11, 'lutff_global/clk')
// (17, 12, 'lutff_global/clk')
// (17, 13, 'lutff_global/clk')
// (17, 14, 'lutff_global/clk')
// (17, 15, 'lutff_global/clk')
// (17, 16, 'lutff_global/clk')
// (17, 17, 'lutff_global/clk')
// (17, 18, 'lutff_global/clk')
// (17, 20, 'lutff_global/clk')
// (17, 21, 'lutff_global/clk')
// (17, 22, 'lutff_global/clk')
// (17, 23, 'lutff_global/clk')
// (17, 24, 'lutff_global/clk')
// (18, 2, 'lutff_global/clk')
// (18, 3, 'lutff_global/clk')
// (18, 4, 'lutff_global/clk')
// (18, 5, 'lutff_global/clk')
// (18, 6, 'lutff_global/clk')
// (18, 7, 'lutff_global/clk')
// (18, 8, 'lutff_global/clk')
// (18, 9, 'lutff_global/clk')
// (18, 10, 'lutff_global/clk')
// (18, 11, 'lutff_global/clk')
// (18, 12, 'lutff_global/clk')
// (18, 13, 'lutff_global/clk')
// (18, 14, 'lutff_global/clk')
// (18, 15, 'lutff_global/clk')
// (18, 16, 'lutff_global/clk')
// (18, 17, 'lutff_global/clk')
// (18, 18, 'lutff_global/clk')
// (18, 19, 'lutff_global/clk')
// (18, 20, 'lutff_global/clk')
// (18, 21, 'lutff_global/clk')
// (18, 22, 'lutff_global/clk')
// (18, 23, 'lutff_global/clk')
// (18, 24, 'lutff_global/clk')
// (19, 5, 'ram/RCLK')
// (19, 6, 'ram/WCLK')
// (19, 7, 'ram/RCLK')
// (19, 8, 'ram/WCLK')
// (19, 9, 'ram/RCLK')
// (19, 10, 'ram/WCLK')
// (19, 11, 'ram/RCLK')
// (19, 12, 'ram/WCLK')
// (19, 13, 'ram/RCLK')
// (19, 14, 'ram/WCLK')
// (19, 15, 'ram/RCLK')
// (19, 16, 'ram/WCLK')
// (20, 1, 'lutff_global/clk')
// (20, 2, 'lutff_global/clk')
// (20, 3, 'lutff_global/clk')
// (20, 4, 'lutff_global/clk')
// (20, 5, 'lutff_global/clk')
// (20, 6, 'lutff_global/clk')
// (20, 8, 'lutff_global/clk')
// (20, 9, 'lutff_global/clk')
// (20, 10, 'lutff_global/clk')
// (20, 11, 'lutff_global/clk')
// (20, 12, 'lutff_global/clk')
// (20, 13, 'lutff_global/clk')
// (20, 14, 'lutff_global/clk')
// (20, 15, 'lutff_global/clk')
// (20, 16, 'lutff_global/clk')
// (20, 17, 'lutff_global/clk')
// (20, 18, 'lutff_global/clk')
// (20, 19, 'lutff_global/clk')
// (20, 20, 'lutff_global/clk')
// (20, 21, 'lutff_global/clk')
// (20, 22, 'lutff_global/clk')
// (20, 23, 'lutff_global/clk')
// (21, 1, 'lutff_global/clk')
// (21, 2, 'lutff_global/clk')
// (21, 3, 'lutff_global/clk')
// (21, 4, 'lutff_global/clk')
// (21, 5, 'lutff_global/clk')
// (21, 6, 'lutff_global/clk')
// (21, 7, 'lutff_global/clk')
// (21, 8, 'lutff_global/clk')
// (21, 9, 'lutff_global/clk')
// (21, 10, 'lutff_global/clk')
// (21, 11, 'lutff_global/clk')
// (21, 12, 'lutff_global/clk')
// (21, 13, 'lutff_global/clk')
// (21, 14, 'lutff_global/clk')
// (21, 15, 'lutff_global/clk')
// (21, 16, 'lutff_global/clk')
// (21, 17, 'lutff_global/clk')
// (21, 18, 'lutff_global/clk')
// (21, 19, 'lutff_global/clk')
// (21, 20, 'lutff_global/clk')
// (21, 21, 'lutff_global/clk')
// (21, 22, 'lutff_global/clk')
// (21, 23, 'lutff_global/clk')
// (21, 24, 'lutff_global/clk')
// (22, 2, 'lutff_global/clk')
// (22, 3, 'lutff_global/clk')
// (22, 5, 'lutff_global/clk')
// (22, 6, 'lutff_global/clk')
// (22, 7, 'lutff_global/clk')
// (22, 8, 'lutff_global/clk')
// (22, 9, 'lutff_global/clk')
// (22, 10, 'lutff_global/clk')
// (22, 11, 'lutff_global/clk')
// (22, 12, 'lutff_global/clk')
// (22, 13, 'lutff_global/clk')
// (22, 14, 'lutff_global/clk')
// (22, 15, 'lutff_global/clk')
// (22, 16, 'lutff_global/clk')
// (22, 17, 'lutff_global/clk')
// (22, 18, 'lutff_global/clk')
// (22, 19, 'lutff_global/clk')
// (22, 20, 'lutff_global/clk')
// (22, 21, 'lutff_global/clk')
// (22, 22, 'lutff_global/clk')
// (22, 23, 'lutff_global/clk')
// (23, 2, 'lutff_global/clk')
// (23, 3, 'lutff_global/clk')
// (23, 5, 'lutff_global/clk')
// (23, 6, 'lutff_global/clk')
// (23, 7, 'lutff_global/clk')
// (23, 8, 'lutff_global/clk')
// (23, 11, 'lutff_global/clk')
// (23, 12, 'lutff_global/clk')
// (23, 13, 'lutff_global/clk')
// (23, 14, 'lutff_global/clk')
// (23, 15, 'lutff_global/clk')
// (23, 16, 'lutff_global/clk')
// (23, 17, 'lutff_global/clk')
// (23, 18, 'lutff_global/clk')
// (23, 19, 'lutff_global/clk')
// (23, 20, 'lutff_global/clk')
// (23, 21, 'lutff_global/clk')
// (23, 22, 'lutff_global/clk')
// (24, 3, 'lutff_global/clk')
// (24, 13, 'lutff_global/clk')
// (24, 14, 'lutff_global/clk')
// (24, 15, 'lutff_global/clk')
// (24, 16, 'lutff_global/clk')
// (24, 17, 'lutff_global/clk')
// (24, 18, 'lutff_global/clk')
// (24, 19, 'lutff_global/clk')
// (24, 20, 'lutff_global/clk')
// (24, 21, 'lutff_global/clk')

wire n3;
// (0, 0, 'glb_netwk_2')
// (17, 12, 'lutff_global/s_r')
// (17, 18, 'neigh_op_tnr_3')
// (17, 19, 'neigh_op_rgt_3')
// (17, 20, 'neigh_op_bnr_3')
// (18, 11, 'lutff_global/s_r')
// (18, 12, 'lutff_global/s_r')
// (18, 13, 'lutff_global/s_r')
// (18, 14, 'lutff_global/s_r')
// (18, 18, 'neigh_op_top_3')
// (18, 19, 'lutff_3/out')
// (18, 19, 'sp4_r_v_b_39')
// (18, 20, 'neigh_op_bot_3')
// (18, 20, 'sp4_r_v_b_26')
// (18, 21, 'sp4_r_v_b_15')
// (18, 22, 'sp4_r_v_b_2')
// (18, 23, 'sp4_r_v_b_39')
// (18, 24, 'sp4_r_v_b_26')
// (18, 25, 'sp4_r_v_b_15')
// (18, 26, 'sp4_r_v_b_2')
// (18, 27, 'sp4_r_v_b_39')
// (18, 28, 'sp4_r_v_b_26')
// (18, 29, 'sp4_r_v_b_15')
// (18, 30, 'sp4_r_v_b_2')
// (19, 18, 'neigh_op_tnl_3')
// (19, 18, 'sp4_v_t_39')
// (19, 19, 'neigh_op_lft_3')
// (19, 19, 'sp4_v_b_39')
// (19, 20, 'neigh_op_bnl_3')
// (19, 20, 'sp4_v_b_26')
// (19, 21, 'sp4_v_b_15')
// (19, 22, 'sp4_v_b_2')
// (19, 22, 'sp4_v_t_39')
// (19, 23, 'sp4_v_b_39')
// (19, 24, 'sp4_v_b_26')
// (19, 25, 'sp4_v_b_15')
// (19, 26, 'sp4_v_b_2')
// (19, 26, 'sp4_v_t_39')
// (19, 27, 'sp4_v_b_39')
// (19, 28, 'sp4_v_b_26')
// (19, 29, 'sp4_v_b_15')
// (19, 30, 'sp4_v_b_2')
// (19, 30, 'sp4_v_t_40')
// (19, 31, 'fabout')
// (19, 31, 'local_g1_0')
// (19, 31, 'span4_vert_40')
// (20, 11, 'lutff_global/s_r')
// (20, 14, 'lutff_global/s_r')
// (21, 10, 'lutff_global/s_r')
// (22, 12, 'lutff_global/s_r')

wire n4;
// (0, 0, 'glb_netwk_3')
// (4, 8, 'lutff_global/cen')
// (4, 9, 'lutff_global/cen')
// (4, 12, 'sp4_r_v_b_42')
// (4, 13, 'sp4_r_v_b_31')
// (4, 14, 'sp4_r_v_b_18')
// (4, 15, 'sp4_r_v_b_7')
// (5, 6, 'lutff_global/cen')
// (5, 8, 'lutff_global/cen')
// (5, 9, 'lutff_global/cen')
// (5, 10, 'lutff_global/cen')
// (5, 11, 'sp4_v_t_42')
// (5, 12, 'lutff_global/cen')
// (5, 12, 'sp4_v_b_42')
// (5, 13, 'lutff_global/cen')
// (5, 13, 'sp4_v_b_31')
// (5, 14, 'local_g1_2')
// (5, 14, 'lutff_7/in_2')
// (5, 14, 'sp4_v_b_18')
// (5, 15, 'sp4_h_r_7')
// (5, 15, 'sp4_v_b_7')
// (5, 16, 'sp4_r_v_b_45')
// (5, 17, 'sp4_r_v_b_32')
// (5, 18, 'sp4_r_v_b_21')
// (5, 19, 'sp4_r_v_b_8')
// (5, 20, 'sp4_r_v_b_41')
// (5, 21, 'sp4_r_v_b_28')
// (5, 22, 'sp4_r_v_b_17')
// (5, 23, 'sp4_r_v_b_4')
// (5, 24, 'sp4_r_v_b_37')
// (5, 25, 'sp4_r_v_b_24')
// (5, 26, 'sp4_r_v_b_13')
// (5, 27, 'sp4_r_v_b_0')
// (5, 28, 'sp4_r_v_b_38')
// (5, 29, 'sp4_r_v_b_27')
// (5, 30, 'sp4_r_v_b_14')
// (6, 15, 'sp4_h_r_18')
// (6, 15, 'sp4_h_r_2')
// (6, 15, 'sp4_v_t_45')
// (6, 16, 'sp4_v_b_45')
// (6, 17, 'sp4_v_b_32')
// (6, 18, 'sp4_v_b_21')
// (6, 19, 'sp4_v_b_8')
// (6, 19, 'sp4_v_t_41')
// (6, 20, 'sp4_v_b_41')
// (6, 21, 'sp4_v_b_28')
// (6, 22, 'sp4_v_b_17')
// (6, 23, 'sp4_v_b_4')
// (6, 23, 'sp4_v_t_37')
// (6, 24, 'sp4_v_b_37')
// (6, 25, 'sp4_v_b_24')
// (6, 26, 'sp4_v_b_13')
// (6, 27, 'sp4_v_b_0')
// (6, 27, 'sp4_v_t_38')
// (6, 28, 'sp4_v_b_38')
// (6, 29, 'sp4_v_b_27')
// (6, 30, 'sp4_v_b_14')
// (6, 31, 'fabout')
// (6, 31, 'local_g0_3')
// (6, 31, 'span4_vert_3')
// (7, 5, 'lutff_global/cen')
// (7, 6, 'lutff_global/cen')
// (7, 7, 'lutff_global/cen')
// (7, 10, 'lutff_global/cen')
// (7, 11, 'lutff_global/cen')
// (7, 12, 'sp4_r_v_b_43')
// (7, 13, 'lutff_global/cen')
// (7, 13, 'sp4_r_v_b_30')
// (7, 14, 'local_g3_3')
// (7, 14, 'lutff_1/in_3')
// (7, 14, 'sp4_r_v_b_19')
// (7, 15, 'sp4_h_r_15')
// (7, 15, 'sp4_h_r_31')
// (7, 15, 'sp4_r_v_b_6')
// (8, 10, 'lutff_global/cen')
// (8, 11, 'lutff_global/cen')
// (8, 11, 'sp4_v_t_43')
// (8, 12, 'sp4_v_b_43')
// (8, 13, 'sp4_v_b_30')
// (8, 14, 'sp4_v_b_19')
// (8, 15, 'sp4_h_r_26')
// (8, 15, 'sp4_h_r_42')
// (8, 15, 'sp4_h_r_6')
// (8, 15, 'sp4_v_b_6')
// (9, 6, 'lutff_global/cen')
// (9, 8, 'lutff_global/cen')
// (9, 9, 'lutff_global/cen')
// (9, 10, 'lutff_global/cen')
// (9, 11, 'lutff_global/cen')
// (9, 13, 'lutff_global/cen')
// (9, 15, 'lutff_global/cen')
// (9, 15, 'sp4_h_l_42')
// (9, 15, 'sp4_h_r_19')
// (9, 15, 'sp4_h_r_39')
// (9, 15, 'sp4_h_r_7')
// (10, 6, 'lutff_global/cen')
// (10, 7, 'lutff_global/cen')
// (10, 8, 'lutff_global/cen')
// (10, 9, 'lutff_global/cen')
// (10, 10, 'lutff_global/cen')
// (10, 11, 'lutff_global/cen')
// (10, 13, 'lutff_global/cen')
// (10, 14, 'lutff_global/cen')
// (10, 15, 'lutff_global/cen')
// (10, 15, 'sp4_h_l_39')
// (10, 15, 'sp4_h_r_18')
// (10, 15, 'sp4_h_r_2')
// (10, 15, 'sp4_h_r_30')
// (10, 16, 'lutff_global/cen')
// (11, 7, 'lutff_global/cen')
// (11, 8, 'lutff_global/cen')
// (11, 9, 'lutff_global/cen')
// (11, 10, 'lutff_global/cen')
// (11, 11, 'lutff_global/cen')
// (11, 14, 'local_g2_5')
// (11, 14, 'lutff_5/in_2')
// (11, 14, 'neigh_op_tnr_5')
// (11, 15, 'neigh_op_rgt_5')
// (11, 15, 'sp4_h_r_15')
// (11, 15, 'sp4_h_r_31')
// (11, 15, 'sp4_h_r_43')
// (11, 16, 'lutff_global/cen')
// (11, 16, 'neigh_op_bnr_5')
// (12, 12, 'lutff_global/cen')
// (12, 13, 'lutff_global/cen')
// (12, 14, 'neigh_op_top_5')
// (12, 15, 'lutff_5/out')
// (12, 15, 'sp4_h_l_43')
// (12, 15, 'sp4_h_r_10')
// (12, 15, 'sp4_h_r_26')
// (12, 15, 'sp4_h_r_42')
// (12, 16, 'lutff_global/cen')
// (12, 16, 'neigh_op_bot_5')
// (13, 7, 'lutff_global/cen')
// (13, 14, 'neigh_op_tnl_5')
// (13, 15, 'neigh_op_lft_5')
// (13, 15, 'sp4_h_l_42')
// (13, 15, 'sp4_h_r_23')
// (13, 15, 'sp4_h_r_39')
// (13, 16, 'neigh_op_bnl_5')
// (14, 15, 'sp4_h_l_39')
// (14, 15, 'sp4_h_r_34')
// (15, 15, 'sp4_h_r_47')
// (16, 15, 'sp4_h_l_47')

reg n5 = 0;
// (0, 0, 'glb_netwk_4')
// (1, 12, 'glb2local_3')
// (1, 12, 'local_g0_7')
// (1, 12, 'lutff_3/in_2')
// (1, 13, 'glb2local_2')
// (1, 13, 'local_g0_6')
// (1, 13, 'lutff_6/in_0')
// (1, 15, 'glb2local_1')
// (1, 15, 'local_g0_5')
// (1, 15, 'lutff_2/in_3')
// (1, 15, 'lutff_3/in_0')
// (2, 10, 'glb2local_0')
// (2, 10, 'local_g0_4')
// (2, 10, 'lutff_7/in_1')
// (2, 13, 'glb2local_2')
// (2, 13, 'local_g0_6')
// (2, 13, 'lutff_4/in_0')
// (2, 14, 'glb2local_0')
// (2, 14, 'local_g0_4')
// (2, 14, 'lutff_1/in_1')
// (2, 14, 'lutff_4/in_2')
// (2, 15, 'glb2local_1')
// (2, 15, 'local_g0_5')
// (2, 15, 'lutff_1/in_0')
// (3, 3, 'glb2local_0')
// (3, 3, 'local_g0_4')
// (3, 3, 'lutff_3/in_1')
// (3, 5, 'glb2local_3')
// (3, 5, 'local_g0_7')
// (3, 5, 'lutff_0/in_3')
// (3, 12, 'glb2local_1')
// (3, 12, 'local_g0_5')
// (3, 12, 'lutff_4/in_3')
// (3, 21, 'glb2local_0')
// (3, 21, 'local_g0_4')
// (3, 21, 'lutff_4/in_0')
// (3, 21, 'lutff_5/in_1')
// (3, 21, 'lutff_7/in_3')
// (4, 9, 'glb2local_0')
// (4, 9, 'local_g0_4')
// (4, 9, 'lutff_3/in_1')
// (4, 15, 'glb2local_2')
// (4, 15, 'local_g0_6')
// (4, 15, 'lutff_2/in_2')
// (5, 1, 'glb2local_1')
// (5, 1, 'local_g0_5')
// (5, 1, 'lutff_3/in_2')
// (5, 6, 'glb2local_2')
// (5, 6, 'glb2local_3')
// (5, 6, 'local_g0_6')
// (5, 6, 'local_g0_7')
// (5, 6, 'lutff_3/in_2')
// (5, 6, 'lutff_5/in_3')
// (5, 6, 'lutff_6/in_2')
// (5, 8, 'glb2local_2')
// (5, 8, 'glb2local_3')
// (5, 8, 'local_g0_6')
// (5, 8, 'local_g0_7')
// (5, 8, 'lutff_1/in_2')
// (5, 8, 'lutff_2/in_1')
// (5, 8, 'lutff_4/in_1')
// (5, 8, 'lutff_7/in_3')
// (5, 9, 'glb2local_2')
// (5, 9, 'local_g0_6')
// (5, 9, 'lutff_0/in_2')
// (5, 9, 'lutff_1/in_3')
// (5, 9, 'lutff_2/in_0')
// (5, 9, 'lutff_3/in_1')
// (5, 9, 'lutff_5/in_1')
// (5, 10, 'glb2local_0')
// (5, 10, 'local_g0_4')
// (5, 10, 'lutff_0/in_0')
// (5, 10, 'lutff_1/in_3')
// (5, 10, 'lutff_2/in_0')
// (5, 17, 'glb2local_0')
// (5, 17, 'local_g0_4')
// (5, 17, 'lutff_1/in_1')
// (7, 1, 'glb2local_0')
// (7, 1, 'local_g0_4')
// (7, 1, 'lutff_5/in_3')
// (7, 1, 'lutff_6/in_0')
// (7, 3, 'glb2local_2')
// (7, 3, 'local_g0_6')
// (7, 3, 'lutff_1/in_1')
// (7, 3, 'lutff_7/in_1')
// (7, 4, 'glb2local_1')
// (7, 4, 'local_g0_5')
// (7, 4, 'lutff_1/in_0')
// (7, 4, 'lutff_2/in_3')
// (7, 4, 'lutff_6/in_3')
// (7, 5, 'glb2local_0')
// (7, 5, 'glb2local_3')
// (7, 5, 'local_g0_4')
// (7, 5, 'local_g0_7')
// (7, 5, 'lutff_0/in_3')
// (7, 5, 'lutff_2/in_2')
// (7, 5, 'lutff_3/in_0')
// (7, 5, 'lutff_4/in_2')
// (7, 5, 'lutff_6/in_1')
// (7, 6, 'glb2local_2')
// (7, 6, 'local_g0_6')
// (7, 6, 'lutff_4/in_2')
// (7, 6, 'lutff_7/in_3')
// (7, 7, 'glb2local_2')
// (7, 7, 'local_g0_6')
// (7, 7, 'lutff_3/in_1')
// (7, 10, 'glb2local_0')
// (7, 10, 'local_g0_4')
// (7, 10, 'lutff_1/in_3')
// (7, 17, 'glb2local_3')
// (7, 17, 'local_g0_7')
// (7, 17, 'lutff_1/in_0')
// (7, 17, 'lutff_2/in_3')
// (7, 17, 'lutff_4/in_1')
// (7, 17, 'lutff_5/in_0')
// (7, 21, 'glb2local_2')
// (7, 21, 'local_g0_6')
// (7, 21, 'lutff_5/in_3')
// (8, 2, 'glb2local_0')
// (8, 2, 'local_g0_4')
// (8, 2, 'lutff_7/in_1')
// (8, 3, 'glb2local_0')
// (8, 3, 'local_g0_4')
// (8, 3, 'lutff_2/in_2')
// (8, 3, 'lutff_7/in_3')
// (8, 4, 'glb2local_1')
// (8, 4, 'local_g0_5')
// (8, 4, 'lutff_1/in_0')
// (8, 5, 'glb2local_1')
// (8, 5, 'local_g0_5')
// (8, 5, 'lutff_4/in_3')
// (8, 5, 'lutff_7/in_0')
// (9, 2, 'glb2local_2')
// (9, 2, 'local_g0_6')
// (9, 2, 'lutff_4/in_0')
// (9, 5, 'glb2local_2')
// (9, 5, 'local_g0_6')
// (9, 5, 'lutff_0/in_2')
// (9, 5, 'lutff_4/in_2')
// (9, 5, 'lutff_5/in_3')
// (9, 6, 'glb2local_3')
// (9, 6, 'local_g0_7')
// (9, 6, 'lutff_1/in_2')
// (9, 8, 'glb2local_3')
// (9, 8, 'local_g0_7')
// (9, 8, 'lutff_1/in_2')
// (9, 8, 'lutff_3/in_0')
// (9, 8, 'lutff_4/in_1')
// (9, 8, 'lutff_6/in_3')
// (9, 11, 'glb2local_3')
// (9, 11, 'local_g0_7')
// (9, 11, 'lutff_6/in_3')
// (10, 2, 'glb2local_2')
// (10, 2, 'local_g0_6')
// (10, 2, 'lutff_0/in_0')
// (10, 2, 'lutff_3/in_1')
// (10, 2, 'lutff_4/in_2')
// (10, 3, 'glb2local_1')
// (10, 3, 'local_g0_5')
// (10, 3, 'lutff_2/in_3')
// (10, 3, 'lutff_6/in_3')
// (10, 3, 'lutff_7/in_0')
// (10, 4, 'glb2local_3')
// (10, 4, 'local_g0_7')
// (10, 4, 'lutff_0/in_1')
// (10, 4, 'lutff_1/in_2')
// (10, 4, 'lutff_2/in_3')
// (10, 4, 'lutff_3/in_2')
// (10, 5, 'glb2local_0')
// (10, 5, 'local_g0_4')
// (10, 5, 'lutff_5/in_1')
// (10, 6, 'glb2local_3')
// (10, 6, 'local_g0_7')
// (10, 6, 'lutff_4/in_1')
// (10, 7, 'glb2local_2')
// (10, 7, 'local_g0_6')
// (10, 7, 'lutff_0/in_0')
// (10, 7, 'lutff_1/in_1')
// (10, 7, 'lutff_5/in_3')
// (10, 7, 'lutff_6/in_2')
// (10, 8, 'glb2local_0')
// (10, 8, 'local_g0_4')
// (10, 8, 'lutff_2/in_0')
// (10, 8, 'lutff_4/in_2')
// (10, 9, 'glb2local_0')
// (10, 9, 'local_g0_4')
// (10, 9, 'lutff_0/in_2')
// (10, 9, 'lutff_4/in_2')
// (10, 9, 'lutff_6/in_0')
// (10, 13, 'glb2local_3')
// (10, 13, 'local_g0_7')
// (10, 13, 'lutff_4/in_1')
// (10, 19, 'glb2local_1')
// (10, 19, 'local_g0_5')
// (10, 19, 'lutff_4/in_1')
// (10, 20, 'glb2local_3')
// (10, 20, 'local_g0_7')
// (10, 20, 'lutff_5/in_2')
// (10, 29, 'neigh_op_tnr_0')
// (10, 30, 'neigh_op_rgt_0')
// (10, 31, 'logic_op_bnr_0')
// (11, 2, 'glb2local_1')
// (11, 2, 'local_g0_5')
// (11, 2, 'lutff_2/in_3')
// (11, 3, 'glb2local_3')
// (11, 3, 'local_g0_7')
// (11, 3, 'lutff_2/in_1')
// (11, 3, 'lutff_5/in_2')
// (11, 3, 'lutff_6/in_3')
// (11, 4, 'glb2local_0')
// (11, 4, 'local_g0_4')
// (11, 4, 'lutff_5/in_1')
// (11, 6, 'glb2local_3')
// (11, 6, 'local_g0_7')
// (11, 6, 'lutff_1/in_0')
// (11, 7, 'glb2local_2')
// (11, 7, 'local_g0_6')
// (11, 7, 'lutff_4/in_0')
// (11, 8, 'glb2local_0')
// (11, 8, 'glb2local_3')
// (11, 8, 'local_g0_4')
// (11, 8, 'local_g0_7')
// (11, 8, 'lutff_2/in_3')
// (11, 8, 'lutff_3/in_1')
// (11, 8, 'lutff_4/in_2')
// (11, 8, 'lutff_5/in_0')
// (11, 8, 'lutff_6/in_1')
// (11, 8, 'lutff_7/in_0')
// (11, 9, 'glb2local_1')
// (11, 9, 'glb2local_2')
// (11, 9, 'local_g0_5')
// (11, 9, 'local_g0_6')
// (11, 9, 'lutff_1/in_2')
// (11, 9, 'lutff_4/in_0')
// (11, 9, 'lutff_5/in_0')
// (11, 15, 'glb2local_2')
// (11, 15, 'local_g0_6')
// (11, 15, 'lutff_3/in_1')
// (11, 19, 'glb2local_1')
// (11, 19, 'local_g0_5')
// (11, 19, 'lutff_4/in_3')
// (11, 19, 'lutff_5/in_2')
// (11, 20, 'glb2local_2')
// (11, 20, 'local_g0_6')
// (11, 20, 'lutff_3/in_3')
// (11, 20, 'lutff_4/in_2')
// (11, 20, 'lutff_6/in_2')
// (11, 21, 'glb2local_3')
// (11, 21, 'local_g0_7')
// (11, 21, 'lutff_4/in_3')
// (11, 21, 'lutff_5/in_2')
// (11, 29, 'neigh_op_top_0')
// (11, 30, 'glb2local_2')
// (11, 30, 'local_g0_6')
// (11, 30, 'lutff_0/in_0')
// (11, 30, 'lutff_0/out')
// (11, 31, 'logic_op_bot_0')
// (12, 2, 'glb2local_3')
// (12, 2, 'local_g0_7')
// (12, 2, 'lutff_3/in_0')
// (12, 11, 'glb2local_1')
// (12, 11, 'local_g0_5')
// (12, 11, 'lutff_3/in_0')
// (12, 14, 'glb2local_1')
// (12, 14, 'local_g0_5')
// (12, 14, 'lutff_7/in_2')
// (12, 16, 'glb2local_2')
// (12, 16, 'local_g0_6')
// (12, 16, 'lutff_2/in_2')
// (12, 17, 'glb2local_1')
// (12, 17, 'local_g0_5')
// (12, 17, 'lutff_1/in_2')
// (12, 18, 'glb2local_3')
// (12, 18, 'local_g0_7')
// (12, 18, 'lutff_2/in_3')
// (12, 19, 'glb2local_2')
// (12, 19, 'local_g0_6')
// (12, 19, 'lutff_1/in_3')
// (12, 19, 'lutff_3/in_1')
// (12, 19, 'lutff_7/in_1')
// (12, 20, 'glb2local_2')
// (12, 20, 'local_g0_6')
// (12, 20, 'lutff_1/in_1')
// (12, 20, 'lutff_4/in_0')
// (12, 20, 'lutff_7/in_3')
// (12, 22, 'glb2local_3')
// (12, 22, 'local_g0_7')
// (12, 22, 'lutff_7/in_2')
// (12, 23, 'glb2local_2')
// (12, 23, 'local_g0_6')
// (12, 23, 'lutff_4/in_2')
// (12, 29, 'neigh_op_tnl_0')
// (12, 30, 'neigh_op_lft_0')
// (12, 31, 'fabout')
// (12, 31, 'local_g1_0')
// (12, 31, 'logic_op_bnl_0')
// (13, 18, 'glb2local_0')
// (13, 18, 'local_g0_4')
// (13, 18, 'lutff_0/in_0')
// (13, 18, 'lutff_2/in_0')
// (13, 18, 'lutff_6/in_0')
// (13, 18, 'lutff_7/in_3')
// (13, 19, 'glb2local_2')
// (13, 19, 'local_g0_6')
// (13, 19, 'lutff_7/in_1')
// (13, 21, 'glb2local_1')
// (13, 21, 'local_g0_5')
// (13, 21, 'lutff_1/in_2')
// (13, 21, 'lutff_2/in_1')
// (13, 21, 'lutff_3/in_2')
// (13, 21, 'lutff_6/in_1')
// (13, 22, 'glb2local_3')
// (13, 22, 'local_g0_7')
// (13, 22, 'lutff_2/in_1')
// (13, 22, 'lutff_3/in_0')
// (13, 22, 'lutff_4/in_1')
// (13, 22, 'lutff_5/in_0')
// (13, 22, 'lutff_6/in_1')
// (13, 23, 'glb2local_1')
// (13, 23, 'local_g0_5')
// (13, 23, 'lutff_7/in_2')
// (14, 1, 'glb2local_3')
// (14, 1, 'local_g0_7')
// (14, 1, 'lutff_0/in_1')
// (14, 16, 'glb2local_1')
// (14, 16, 'local_g0_5')
// (14, 16, 'lutff_1/in_0')
// (14, 16, 'lutff_7/in_2')
// (14, 17, 'glb2local_0')
// (14, 17, 'local_g0_4')
// (14, 17, 'lutff_5/in_3')
// (14, 21, 'glb2local_0')
// (14, 21, 'local_g0_4')
// (14, 21, 'lutff_1/in_1')
// (14, 21, 'lutff_5/in_3')
// (15, 17, 'glb2local_2')
// (15, 17, 'local_g0_6')
// (15, 17, 'lutff_0/in_0')
// (15, 20, 'glb2local_2')
// (15, 20, 'local_g0_6')
// (15, 20, 'lutff_0/in_0')
// (15, 20, 'lutff_2/in_0')
// (15, 20, 'lutff_6/in_0')
// (17, 20, 'glb2local_3')
// (17, 20, 'local_g0_7')
// (17, 20, 'lutff_4/in_3')

reg n6 = 0;
// (0, 0, 'glb_netwk_5')
// (1, 4, 'glb2local_0')
// (1, 4, 'glb2local_1')
// (1, 4, 'local_g0_4')
// (1, 4, 'local_g0_5')
// (1, 4, 'lutff_4/in_1')
// (1, 4, 'lutff_5/in_1')
// (1, 5, 'glb2local_3')
// (1, 5, 'local_g0_7')
// (1, 5, 'lutff_6/in_1')
// (2, 1, 'glb2local_3')
// (2, 1, 'local_g0_7')
// (2, 1, 'lutff_6/in_1')
// (2, 2, 'glb2local_3')
// (2, 2, 'local_g0_7')
// (2, 2, 'lutff_0/in_1')
// (2, 2, 'lutff_5/in_0')
// (2, 4, 'glb2local_2')
// (2, 4, 'local_g0_6')
// (2, 4, 'lutff_7/in_3')
// (2, 5, 'glb2local_0')
// (2, 5, 'glb2local_3')
// (2, 5, 'local_g0_4')
// (2, 5, 'local_g0_7')
// (2, 5, 'lutff_3/in_3')
// (2, 5, 'lutff_5/in_0')
// (2, 5, 'lutff_7/in_3')
// (2, 6, 'glb2local_0')
// (2, 6, 'local_g0_4')
// (2, 6, 'lutff_0/in_2')
// (2, 7, 'glb2local_3')
// (2, 7, 'local_g0_7')
// (2, 7, 'lutff_1/in_2')
// (2, 7, 'lutff_2/in_1')
// (3, 1, 'glb2local_2')
// (3, 1, 'local_g0_6')
// (3, 1, 'lutff_0/in_0')
// (3, 1, 'lutff_2/in_2')
// (3, 2, 'glb2local_2')
// (3, 2, 'local_g0_6')
// (3, 2, 'lutff_2/in_2')
// (3, 2, 'lutff_4/in_0')
// (3, 4, 'glb2local_0')
// (3, 4, 'glb2local_1')
// (3, 4, 'local_g0_4')
// (3, 4, 'local_g0_5')
// (3, 4, 'lutff_5/in_3')
// (3, 4, 'lutff_7/in_2')
// (3, 5, 'glb2local_1')
// (3, 5, 'local_g0_5')
// (3, 5, 'lutff_1/in_2')
// (3, 5, 'lutff_6/in_3')
// (3, 6, 'glb2local_2')
// (3, 6, 'local_g0_6')
// (3, 6, 'lutff_1/in_3')
// (3, 6, 'lutff_7/in_3')
// (3, 7, 'glb2local_2')
// (3, 7, 'local_g0_6')
// (3, 7, 'lutff_4/in_0')
// (4, 1, 'glb2local_1')
// (4, 1, 'local_g0_5')
// (4, 1, 'lutff_2/in_1')
// (4, 1, 'lutff_3/in_2')
// (4, 1, 'lutff_6/in_3')
// (4, 2, 'glb2local_0')
// (4, 2, 'glb2local_1')
// (4, 2, 'local_g0_4')
// (4, 2, 'local_g0_5')
// (4, 2, 'lutff_3/in_1')
// (4, 2, 'lutff_4/in_1')
// (4, 3, 'glb2local_1')
// (4, 3, 'local_g0_5')
// (4, 3, 'lutff_1/in_0')
// (4, 3, 'lutff_7/in_0')
// (4, 3, 'neigh_op_tnr_5')
// (4, 4, 'glb2local_1')
// (4, 4, 'local_g0_5')
// (4, 4, 'lutff_1/in_2')
// (4, 4, 'lutff_3/in_2')
// (4, 4, 'neigh_op_rgt_5')
// (4, 4, 'sp4_r_v_b_42')
// (4, 5, 'glb2local_1')
// (4, 5, 'local_g0_5')
// (4, 5, 'lutff_3/in_2')
// (4, 5, 'lutff_5/in_2')
// (4, 5, 'lutff_6/in_3')
// (4, 5, 'neigh_op_bnr_5')
// (4, 5, 'sp4_r_v_b_31')
// (4, 6, 'glb2local_3')
// (4, 6, 'local_g0_7')
// (4, 6, 'lutff_0/in_1')
// (4, 6, 'sp4_r_v_b_18')
// (4, 7, 'glb2local_0')
// (4, 7, 'glb2local_3')
// (4, 7, 'local_g0_4')
// (4, 7, 'local_g0_7')
// (4, 7, 'lutff_1/in_3')
// (4, 7, 'lutff_3/in_0')
// (4, 7, 'lutff_7/in_1')
// (4, 7, 'sp4_r_v_b_7')
// (5, 1, 'glb2local_0')
// (5, 1, 'local_g0_4')
// (5, 1, 'lutff_0/in_2')
// (5, 1, 'lutff_7/in_3')
// (5, 2, 'glb2local_1')
// (5, 2, 'local_g0_5')
// (5, 2, 'lutff_0/in_1')
// (5, 3, 'glb2local_0')
// (5, 3, 'local_g0_4')
// (5, 3, 'lutff_4/in_2')
// (5, 3, 'lutff_5/in_3')
// (5, 3, 'lutff_7/in_3')
// (5, 3, 'neigh_op_top_5')
// (5, 3, 'sp4_h_r_7')
// (5, 3, 'sp4_v_t_42')
// (5, 4, 'glb2local_0')
// (5, 4, 'local_g0_4')
// (5, 4, 'lutff_1/in_3')
// (5, 4, 'lutff_3/in_3')
// (5, 4, 'lutff_4/in_0')
// (5, 4, 'lutff_5/in_1')
// (5, 4, 'lutff_5/out')
// (5, 4, 'lutff_6/in_2')
// (5, 4, 'lutff_7/in_1')
// (5, 4, 'sp4_v_b_42')
// (5, 5, 'glb2local_0')
// (5, 5, 'glb2local_1')
// (5, 5, 'local_g0_4')
// (5, 5, 'local_g0_5')
// (5, 5, 'lutff_0/in_3')
// (5, 5, 'lutff_1/in_0')
// (5, 5, 'lutff_5/in_1')
// (5, 5, 'neigh_op_bot_5')
// (5, 5, 'sp4_v_b_31')
// (5, 6, 'glb2local_1')
// (5, 6, 'local_g0_5')
// (5, 6, 'lutff_4/in_3')
// (5, 6, 'lutff_7/in_2')
// (5, 6, 'sp4_v_b_18')
// (5, 7, 'glb2local_0')
// (5, 7, 'local_g0_4')
// (5, 7, 'lutff_5/in_1')
// (5, 7, 'lutff_6/in_2')
// (5, 7, 'sp4_v_b_7')
// (6, 3, 'neigh_op_tnl_5')
// (6, 3, 'sp4_h_r_18')
// (6, 4, 'neigh_op_lft_5')
// (6, 5, 'neigh_op_bnl_5')
// (7, 1, 'glb2local_1')
// (7, 1, 'glb2local_2')
// (7, 1, 'local_g0_5')
// (7, 1, 'local_g0_6')
// (7, 1, 'lutff_1/in_1')
// (7, 1, 'lutff_2/in_3')
// (7, 3, 'sp4_h_r_31')
// (8, 1, 'glb2local_2')
// (8, 1, 'local_g0_6')
// (8, 1, 'lutff_1/in_1')
// (8, 1, 'lutff_6/in_0')
// (8, 1, 'sp4_r_v_b_25')
// (8, 2, 'glb2local_2')
// (8, 2, 'local_g0_6')
// (8, 2, 'lutff_5/in_1')
// (8, 2, 'sp4_r_v_b_12')
// (8, 3, 'sp4_h_r_42')
// (8, 3, 'sp4_r_v_b_1')
// (9, 0, 'span4_horz_r_0')
// (9, 0, 'span4_vert_25')
// (9, 1, 'glb2local_0')
// (9, 1, 'glb2local_3')
// (9, 1, 'local_g0_4')
// (9, 1, 'local_g0_7')
// (9, 1, 'lutff_1/in_2')
// (9, 1, 'lutff_4/in_2')
// (9, 1, 'sp4_v_b_25')
// (9, 2, 'glb2local_3')
// (9, 2, 'local_g0_7')
// (9, 2, 'lutff_3/in_2')
// (9, 2, 'lutff_5/in_2')
// (9, 2, 'lutff_6/in_3')
// (9, 2, 'sp4_v_b_12')
// (9, 3, 'glb2local_1')
// (9, 3, 'local_g0_5')
// (9, 3, 'lutff_5/in_0')
// (9, 3, 'sp4_h_l_42')
// (9, 3, 'sp4_v_b_1')
// (9, 4, 'glb2local_0')
// (9, 4, 'glb2local_3')
// (9, 4, 'local_g0_4')
// (9, 4, 'local_g0_7')
// (9, 4, 'lutff_5/in_3')
// (9, 4, 'lutff_7/in_2')
// (10, 0, 'span4_horz_r_4')
// (10, 1, 'glb2local_0')
// (10, 1, 'glb2local_1')
// (10, 1, 'local_g0_4')
// (10, 1, 'local_g0_5')
// (10, 1, 'lutff_0/in_1')
// (10, 1, 'lutff_4/in_3')
// (10, 1, 'lutff_6/in_2')
// (10, 2, 'glb2local_0')
// (10, 2, 'glb2local_1')
// (10, 2, 'local_g0_4')
// (10, 2, 'local_g0_5')
// (10, 2, 'lutff_1/in_2')
// (10, 2, 'lutff_2/in_1')
// (10, 2, 'lutff_6/in_2')
// (10, 3, 'glb2local_3')
// (10, 3, 'local_g0_7')
// (10, 3, 'lutff_1/in_0')
// (10, 3, 'lutff_4/in_1')
// (10, 4, 'glb2local_1')
// (10, 4, 'local_g0_5')
// (10, 4, 'lutff_4/in_3')
// (11, 0, 'span4_horz_r_8')
// (11, 2, 'glb2local_3')
// (11, 2, 'local_g0_7')
// (11, 2, 'lutff_3/in_0')
// (12, 0, 'fabout')
// (12, 0, 'local_g1_4')
// (12, 0, 'span4_horz_r_12')
// (13, 0, 'span4_horz_l_12')

reg n7 = 0;
// (0, 0, 'glb_netwk_6')
// (5, 0, 'span4_horz_r_3')
// (6, 0, 'fabout')
// (6, 0, 'local_g0_7')
// (6, 0, 'span4_horz_r_7')
// (7, 0, 'span4_horz_r_11')
// (8, 0, 'span4_horz_r_15')
// (8, 1, 'sp4_r_v_b_19')
// (8, 2, 'sp4_r_v_b_6')
// (9, 0, 'span4_horz_l_15')
// (9, 0, 'span4_vert_19')
// (9, 1, 'sp4_v_b_19')
// (9, 2, 'sp4_h_r_6')
// (9, 2, 'sp4_v_b_6')
// (10, 2, 'sp4_h_r_19')
// (11, 2, 'sp4_h_r_30')
// (12, 2, 'sp4_h_r_43')
// (13, 2, 'sp4_h_l_43')
// (13, 2, 'sp4_h_r_6')
// (14, 2, 'sp4_h_r_19')
// (15, 2, 'sp4_h_r_30')
// (16, 2, 'sp4_h_r_43')
// (17, 2, 'sp4_h_l_43')
// (17, 2, 'sp4_h_r_10')
// (18, 2, 'sp4_h_r_23')
// (19, 2, 'sp4_h_r_34')
// (19, 3, 'sp4_r_v_b_42')
// (19, 4, 'sp4_r_v_b_31')
// (19, 5, 'sp4_r_v_b_18')
// (19, 6, 'sp4_r_v_b_7')
// (20, 1, 'neigh_op_tnr_1')
// (20, 1, 'sp4_r_v_b_47')
// (20, 2, 'neigh_op_rgt_1')
// (20, 2, 'sp4_h_r_47')
// (20, 2, 'sp4_h_r_7')
// (20, 2, 'sp4_r_v_b_34')
// (20, 2, 'sp4_v_t_42')
// (20, 3, 'neigh_op_bnr_1')
// (20, 3, 'sp4_r_v_b_23')
// (20, 3, 'sp4_v_b_42')
// (20, 4, 'local_g2_2')
// (20, 4, 'lutff_4/in_0')
// (20, 4, 'lutff_5/in_3')
// (20, 4, 'sp4_r_v_b_10')
// (20, 4, 'sp4_v_b_31')
// (20, 5, 'local_g0_2')
// (20, 5, 'lutff_7/in_3')
// (20, 5, 'sp4_v_b_18')
// (20, 6, 'sp4_v_b_7')
// (21, 0, 'span4_vert_47')
// (21, 1, 'neigh_op_top_1')
// (21, 1, 'sp4_r_v_b_14')
// (21, 1, 'sp4_r_v_b_46')
// (21, 1, 'sp4_v_b_47')
// (21, 2, 'lutff_1/out')
// (21, 2, 'sp4_h_l_47')
// (21, 2, 'sp4_h_r_18')
// (21, 2, 'sp4_h_r_2')
// (21, 2, 'sp4_r_v_b_3')
// (21, 2, 'sp4_r_v_b_35')
// (21, 2, 'sp4_v_b_34')
// (21, 3, 'lutff_global/s_r')
// (21, 3, 'neigh_op_bot_1')
// (21, 3, 'sp4_r_v_b_22')
// (21, 3, 'sp4_r_v_b_46')
// (21, 3, 'sp4_v_b_23')
// (21, 4, 'lutff_global/s_r')
// (21, 4, 'sp4_r_v_b_11')
// (21, 4, 'sp4_r_v_b_35')
// (21, 4, 'sp4_v_b_10')
// (21, 5, 'lutff_global/s_r')
// (21, 5, 'sp4_r_v_b_22')
// (21, 6, 'sp4_r_v_b_11')
// (22, 0, 'span4_vert_14')
// (22, 0, 'span4_vert_46')
// (22, 1, 'neigh_op_tnl_1')
// (22, 1, 'sp4_v_b_14')
// (22, 1, 'sp4_v_b_46')
// (22, 2, 'neigh_op_lft_1')
// (22, 2, 'sp4_h_r_15')
// (22, 2, 'sp4_h_r_31')
// (22, 2, 'sp4_v_b_3')
// (22, 2, 'sp4_v_b_35')
// (22, 2, 'sp4_v_t_46')
// (22, 3, 'neigh_op_bnl_1')
// (22, 3, 'sp4_v_b_22')
// (22, 3, 'sp4_v_b_46')
// (22, 4, 'local_g0_3')
// (22, 4, 'lutff_3/in_2')
// (22, 4, 'sp4_v_b_11')
// (22, 4, 'sp4_v_b_35')
// (22, 5, 'local_g0_6')
// (22, 5, 'local_g1_6')
// (22, 5, 'lutff_2/in_2')
// (22, 5, 'lutff_7/in_2')
// (22, 5, 'sp4_v_b_22')
// (22, 6, 'sp4_v_b_11')
// (23, 2, 'sp4_h_r_26')
// (23, 2, 'sp4_h_r_42')
// (24, 2, 'sp4_h_l_42')
// (24, 2, 'sp4_h_r_39')
// (24, 3, 'lutff_global/s_r')
// (25, 2, 'sp4_h_l_39')

wire n8;
// (0, 0, 'glb_netwk_7')
// (0, 8, 'sp12_h_r_4')
// (1, 8, 'glb2local_0')
// (1, 8, 'local_g0_4')
// (1, 8, 'local_g0_7')
// (1, 8, 'lutff_3/in_2')
// (1, 8, 'lutff_6/in_2')
// (1, 8, 'sp12_h_r_7')
// (1, 9, 'sp4_r_v_b_36')
// (1, 10, 'sp4_r_v_b_25')
// (1, 11, 'sp4_r_v_b_12')
// (1, 12, 'sp4_r_v_b_1')
// (2, 8, 'sp12_h_r_8')
// (2, 8, 'sp4_v_t_36')
// (2, 9, 'local_g2_4')
// (2, 9, 'lutff_2/in_2')
// (2, 9, 'sp4_v_b_36')
// (2, 10, 'sp4_v_b_25')
// (2, 11, 'sp4_v_b_12')
// (2, 12, 'sp4_h_r_8')
// (2, 12, 'sp4_v_b_1')
// (3, 8, 'sp12_h_r_11')
// (3, 12, 'sp4_h_r_21')
// (3, 13, 'glb2local_0')
// (3, 13, 'local_g0_4')
// (3, 13, 'lutff_2/in_2')
// (3, 17, 'sp4_r_v_b_45')
// (3, 18, 'sp4_h_r_6')
// (3, 18, 'sp4_r_v_b_32')
// (3, 19, 'sp4_r_v_b_21')
// (3, 20, 'sp4_r_v_b_8')
// (3, 21, 'sp4_h_r_6')
// (4, 8, 'glb2local_0')
// (4, 8, 'glb2local_3')
// (4, 8, 'local_g0_4')
// (4, 8, 'local_g0_7')
// (4, 8, 'lutff_1/in_2')
// (4, 8, 'lutff_2/in_0')
// (4, 8, 'sp12_h_r_12')
// (4, 12, 'sp4_h_r_32')
// (4, 13, 'glb2local_1')
// (4, 13, 'glb2local_2')
// (4, 13, 'local_g0_5')
// (4, 13, 'local_g0_6')
// (4, 13, 'lutff_1/in_1')
// (4, 13, 'lutff_2/in_1')
// (4, 16, 'sp4_v_t_45')
// (4, 17, 'sp4_v_b_45')
// (4, 18, 'glb2local_0')
// (4, 18, 'glb2local_1')
// (4, 18, 'local_g0_3')
// (4, 18, 'local_g0_4')
// (4, 18, 'local_g0_5')
// (4, 18, 'lutff_1/in_1')
// (4, 18, 'lutff_2/in_1')
// (4, 18, 'lutff_3/in_2')
// (4, 18, 'lutff_4/in_1')
// (4, 18, 'lutff_5/in_2')
// (4, 18, 'lutff_6/in_1')
// (4, 18, 'lutff_7/in_2')
// (4, 18, 'sp4_h_r_19')
// (4, 18, 'sp4_v_b_32')
// (4, 19, 'glb2local_2')
// (4, 19, 'glb2local_3')
// (4, 19, 'local_g0_5')
// (4, 19, 'local_g0_6')
// (4, 19, 'local_g0_7')
// (4, 19, 'lutff_0/in_2')
// (4, 19, 'lutff_1/in_2')
// (4, 19, 'lutff_2/in_1')
// (4, 19, 'lutff_3/in_1')
// (4, 19, 'sp4_v_b_21')
// (4, 20, 'sp4_h_r_8')
// (4, 20, 'sp4_v_b_8')
// (4, 21, 'local_g0_3')
// (4, 21, 'lutff_3/in_2')
// (4, 21, 'sp4_h_r_19')
// (5, 6, 'glb2local_0')
// (5, 6, 'local_g0_4')
// (5, 6, 'lutff_1/in_1')
// (5, 8, 'sp12_h_r_15')
// (5, 12, 'sp4_h_r_45')
// (5, 18, 'sp4_h_r_30')
// (5, 20, 'sp4_h_r_21')
// (5, 21, 'sp4_h_r_30')
// (6, 8, 'sp12_h_r_16')
// (6, 12, 'sp4_h_l_45')
// (6, 12, 'sp4_h_r_8')
// (6, 18, 'sp4_h_r_43')
// (6, 20, 'sp4_h_r_32')
// (6, 21, 'sp4_h_r_43')
// (7, 8, 'sp12_h_r_19')
// (7, 9, 'glb2local_0')
// (7, 9, 'glb2local_3')
// (7, 9, 'local_g0_4')
// (7, 9, 'local_g0_7')
// (7, 9, 'lutff_1/in_1')
// (7, 9, 'lutff_2/in_1')
// (7, 9, 'lutff_3/in_2')
// (7, 9, 'lutff_4/in_2')
// (7, 12, 'sp4_h_r_21')
// (7, 18, 'sp4_h_l_43')
// (7, 18, 'sp4_h_r_3')
// (7, 20, 'sp4_h_r_45')
// (7, 21, 'local_g1_2')
// (7, 21, 'lutff_1/in_2')
// (7, 21, 'sp4_h_l_43')
// (7, 21, 'sp4_h_r_10')
// (8, 8, 'sp12_h_r_20')
// (8, 12, 'sp4_h_r_32')
// (8, 17, 'glb2local_0')
// (8, 17, 'glb2local_1')
// (8, 17, 'local_g0_4')
// (8, 17, 'local_g0_5')
// (8, 17, 'lutff_5/in_1')
// (8, 17, 'lutff_6/in_1')
// (8, 18, 'sp4_h_r_14')
// (8, 19, 'glb2local_0')
// (8, 19, 'local_g0_4')
// (8, 19, 'lutff_7/in_1')
// (8, 20, 'glb2local_2')
// (8, 20, 'local_g0_6')
// (8, 20, 'lutff_6/in_2')
// (8, 20, 'sp4_h_l_45')
// (8, 20, 'sp4_h_r_5')
// (8, 21, 'sp4_h_r_23')
// (9, 8, 'sp12_h_r_23')
// (9, 12, 'glb2local_0')
// (9, 12, 'glb2local_1')
// (9, 12, 'local_g0_4')
// (9, 12, 'local_g0_5')
// (9, 12, 'lutff_1/in_1')
// (9, 12, 'lutff_2/in_1')
// (9, 12, 'sp4_h_r_45')
// (9, 16, 'glb2local_1')
// (9, 16, 'glb2local_2')
// (9, 16, 'local_g0_5')
// (9, 16, 'local_g0_6')
// (9, 16, 'lutff_5/in_2')
// (9, 16, 'lutff_6/in_2')
// (9, 18, 'glb2local_0')
// (9, 18, 'local_g0_4')
// (9, 18, 'lutff_7/in_1')
// (9, 18, 'sp4_h_r_27')
// (9, 20, 'glb2local_2')
// (9, 20, 'glb2local_3')
// (9, 20, 'local_g0_6')
// (9, 20, 'local_g0_7')
// (9, 20, 'lutff_1/in_2')
// (9, 20, 'lutff_2/in_1')
// (9, 20, 'lutff_3/in_1')
// (9, 20, 'lutff_4/in_2')
// (9, 20, 'lutff_5/in_2')
// (9, 20, 'lutff_6/in_1')
// (9, 20, 'lutff_7/in_2')
// (9, 20, 'sp4_h_r_16')
// (9, 21, 'glb2local_0')
// (9, 21, 'local_g0_4')
// (9, 21, 'lutff_0/in_0')
// (9, 21, 'sp4_h_r_34')
// (10, 8, 'sp12_h_l_23')
// (10, 8, 'sp12_h_r_0')
// (10, 11, 'sp4_r_v_b_46')
// (10, 12, 'sp4_h_l_45')
// (10, 12, 'sp4_h_r_5')
// (10, 12, 'sp4_r_v_b_35')
// (10, 13, 'sp4_r_v_b_22')
// (10, 14, 'sp4_r_v_b_11')
// (10, 15, 'sp4_r_v_b_45')
// (10, 16, 'sp4_r_v_b_32')
// (10, 17, 'sp4_r_v_b_21')
// (10, 18, 'sp4_h_r_38')
// (10, 18, 'sp4_r_v_b_8')
// (10, 20, 'sp4_h_r_29')
// (10, 21, 'sp4_h_r_47')
// (11, 1, 'glb2local_1')
// (11, 1, 'local_g0_5')
// (11, 1, 'lutff_2/in_1')
// (11, 1, 'lutff_3/in_2')
// (11, 1, 'lutff_4/in_1')
// (11, 8, 'sp12_h_r_3')
// (11, 10, 'sp4_v_t_46')
// (11, 11, 'glb2local_1')
// (11, 11, 'local_g0_5')
// (11, 11, 'local_g2_6')
// (11, 11, 'lutff_1/in_2')
// (11, 11, 'lutff_2/in_2')
// (11, 11, 'lutff_3/in_2')
// (11, 11, 'sp4_v_b_46')
// (11, 12, 'sp4_h_r_16')
// (11, 12, 'sp4_v_b_35')
// (11, 13, 'sp4_v_b_22')
// (11, 14, 'sp4_v_b_11')
// (11, 14, 'sp4_v_t_45')
// (11, 15, 'sp4_v_b_45')
// (11, 16, 'sp4_v_b_32')
// (11, 17, 'sp4_v_b_21')
// (11, 18, 'sp4_h_l_38')
// (11, 18, 'sp4_h_r_3')
// (11, 18, 'sp4_v_b_8')
// (11, 20, 'sp4_h_r_40')
// (11, 21, 'sp4_h_l_47')
// (11, 21, 'sp4_h_r_7')
// (12, 1, 'glb2local_2')
// (12, 1, 'local_g0_6')
// (12, 1, 'lutff_4/in_2')
// (12, 3, 'glb2local_0')
// (12, 3, 'local_g0_4')
// (12, 3, 'lutff_1/in_1')
// (12, 3, 'lutff_2/in_2')
// (12, 3, 'lutff_3/in_1')
// (12, 8, 'sp12_h_r_4')
// (12, 12, 'sp4_h_r_29')
// (12, 18, 'sp4_h_r_14')
// (12, 20, 'sp4_h_l_40')
// (12, 20, 'sp4_h_r_2')
// (12, 21, 'sp4_h_r_18')
// (13, 1, 'glb2local_3')
// (13, 1, 'local_g0_7')
// (13, 1, 'lutff_2/in_1')
// (13, 1, 'lutff_4/in_1')
// (13, 8, 'sp12_h_r_7')
// (13, 12, 'sp4_h_r_40')
// (13, 14, 'sp4_r_v_b_40')
// (13, 15, 'sp4_r_v_b_29')
// (13, 16, 'sp4_r_v_b_16')
// (13, 17, 'local_g1_5')
// (13, 17, 'lutff_2/in_2')
// (13, 17, 'lutff_4/in_2')
// (13, 17, 'lutff_6/in_2')
// (13, 17, 'sp4_r_v_b_5')
// (13, 18, 'sp4_h_r_27')
// (13, 20, 'glb2local_1')
// (13, 20, 'glb2local_2')
// (13, 20, 'local_g0_5')
// (13, 20, 'local_g0_6')
// (13, 20, 'lutff_1/in_2')
// (13, 20, 'lutff_2/in_2')
// (13, 20, 'lutff_3/in_1')
// (13, 20, 'lutff_4/in_1')
// (13, 20, 'lutff_5/in_2')
// (13, 20, 'lutff_6/in_0')
// (13, 20, 'sp4_h_r_15')
// (13, 21, 'sp4_h_r_31')
// (14, 8, 'sp12_h_r_8')
// (14, 12, 'sp4_h_l_40')
// (14, 12, 'sp4_h_r_5')
// (14, 13, 'sp4_v_t_40')
// (14, 14, 'sp4_v_b_40')
// (14, 15, 'sp4_v_b_29')
// (14, 16, 'sp4_v_b_16')
// (14, 17, 'sp4_h_r_5')
// (14, 17, 'sp4_v_b_5')
// (14, 18, 'sp4_h_r_38')
// (14, 20, 'sp4_h_r_26')
// (14, 21, 'sp4_h_r_42')
// (14, 22, 'glb2local_3')
// (14, 22, 'local_g0_7')
// (14, 22, 'lutff_6/in_1')
// (14, 23, 'glb2local_2')
// (14, 23, 'local_g0_6')
// (14, 23, 'lutff_4/in_2')
// (14, 23, 'lutff_5/in_1')
// (14, 23, 'lutff_6/in_2')
// (15, 8, 'sp12_h_r_11')
// (15, 12, 'sp4_h_r_16')
// (15, 17, 'sp4_h_r_16')
// (15, 17, 'sp4_r_v_b_41')
// (15, 18, 'glb2local_0')
// (15, 18, 'glb2local_1')
// (15, 18, 'local_g0_4')
// (15, 18, 'local_g0_5')
// (15, 18, 'local_g1_4')
// (15, 18, 'lutff_1/in_1')
// (15, 18, 'lutff_2/in_1')
// (15, 18, 'lutff_3/in_2')
// (15, 18, 'lutff_4/in_1')
// (15, 18, 'lutff_5/in_2')
// (15, 18, 'lutff_6/in_1')
// (15, 18, 'lutff_7/in_2')
// (15, 18, 'sp4_h_l_38')
// (15, 18, 'sp4_h_r_3')
// (15, 18, 'sp4_r_v_b_28')
// (15, 19, 'glb2local_0')
// (15, 19, 'local_g0_4')
// (15, 19, 'local_g3_1')
// (15, 19, 'lutff_0/in_2')
// (15, 19, 'lutff_1/in_1')
// (15, 19, 'lutff_2/in_2')
// (15, 19, 'lutff_3/in_1')
// (15, 19, 'sp4_r_v_b_17')
// (15, 20, 'glb2local_0')
// (15, 20, 'local_g0_4')
// (15, 20, 'lutff_3/in_3')
// (15, 20, 'sp4_h_r_39')
// (15, 20, 'sp4_r_v_b_4')
// (15, 21, 'sp4_h_l_42')
// (15, 21, 'sp4_h_r_7')
// (16, 8, 'sp12_h_r_12')
// (16, 12, 'sp4_h_r_29')
// (16, 16, 'sp4_v_t_41')
// (16, 17, 'sp4_h_r_29')
// (16, 17, 'sp4_r_v_b_36')
// (16, 17, 'sp4_v_b_41')
// (16, 18, 'local_g2_4')
// (16, 18, 'lutff_2/in_2')
// (16, 18, 'lutff_4/in_2')
// (16, 18, 'lutff_6/in_2')
// (16, 18, 'sp4_h_r_14')
// (16, 18, 'sp4_r_v_b_25')
// (16, 18, 'sp4_v_b_28')
// (16, 19, 'local_g1_1')
// (16, 19, 'lutff_0/in_2')
// (16, 19, 'lutff_2/in_2')
// (16, 19, 'sp4_r_v_b_12')
// (16, 19, 'sp4_v_b_17')
// (16, 20, 'sp4_h_l_39')
// (16, 20, 'sp4_h_r_11')
// (16, 20, 'sp4_r_v_b_1')
// (16, 20, 'sp4_v_b_4')
// (16, 21, 'sp4_h_r_18')
// (17, 1, 'sp4_r_v_b_45')
// (17, 2, 'sp4_r_v_b_32')
// (17, 3, 'sp4_r_v_b_21')
// (17, 4, 'sp4_r_v_b_8')
// (17, 5, 'sp4_r_v_b_39')
// (17, 5, 'sp4_r_v_b_40')
// (17, 6, 'local_g1_5')
// (17, 6, 'lutff_1/in_1')
// (17, 6, 'lutff_3/in_1')
// (17, 6, 'lutff_5/in_1')
// (17, 6, 'lutff_7/in_1')
// (17, 6, 'sp4_r_v_b_26')
// (17, 6, 'sp4_r_v_b_29')
// (17, 7, 'local_g2_7')
// (17, 7, 'lutff_1/in_2')
// (17, 7, 'lutff_3/in_2')
// (17, 7, 'sp4_r_v_b_15')
// (17, 7, 'sp4_r_v_b_16')
// (17, 8, 'sp12_h_r_15')
// (17, 8, 'sp4_r_v_b_2')
// (17, 8, 'sp4_r_v_b_5')
// (17, 9, 'sp4_r_v_b_39')
// (17, 10, 'glb2local_0')
// (17, 10, 'local_g0_4')
// (17, 10, 'lutff_6/in_0')
// (17, 10, 'sp4_r_v_b_26')
// (17, 11, 'sp4_r_v_b_15')
// (17, 12, 'sp4_h_r_40')
// (17, 12, 'sp4_r_v_b_2')
// (17, 16, 'sp4_v_t_36')
// (17, 17, 'sp4_h_r_40')
// (17, 17, 'sp4_v_b_36')
// (17, 18, 'sp4_h_r_27')
// (17, 18, 'sp4_v_b_25')
// (17, 19, 'local_g0_4')
// (17, 19, 'lutff_2/in_2')
// (17, 19, 'lutff_4/in_2')
// (17, 19, 'lutff_6/in_2')
// (17, 19, 'sp4_v_b_12')
// (17, 20, 'sp4_h_r_1')
// (17, 20, 'sp4_h_r_22')
// (17, 20, 'sp4_v_b_1')
// (17, 21, 'sp4_h_r_31')
// (18, 0, 'span4_horz_r_3')
// (18, 0, 'span4_vert_45')
// (18, 1, 'glb2local_1')
// (18, 1, 'local_g0_5')
// (18, 1, 'local_g3_5')
// (18, 1, 'lutff_1/in_2')
// (18, 1, 'lutff_2/in_1')
// (18, 1, 'lutff_3/in_2')
// (18, 1, 'lutff_4/in_2')
// (18, 1, 'sp4_v_b_45')
// (18, 2, 'sp4_v_b_32')
// (18, 3, 'sp4_v_b_21')
// (18, 4, 'sp4_h_r_8')
// (18, 4, 'sp4_v_b_8')
// (18, 4, 'sp4_v_t_39')
// (18, 4, 'sp4_v_t_40')
// (18, 5, 'sp4_v_b_39')
// (18, 5, 'sp4_v_b_40')
// (18, 6, 'sp4_v_b_26')
// (18, 6, 'sp4_v_b_29')
// (18, 7, 'sp4_v_b_15')
// (18, 7, 'sp4_v_b_16')
// (18, 8, 'sp12_h_r_16')
// (18, 8, 'sp4_h_r_0')
// (18, 8, 'sp4_v_b_2')
// (18, 8, 'sp4_v_b_5')
// (18, 8, 'sp4_v_t_39')
// (18, 9, 'sp4_v_b_39')
// (18, 10, 'sp4_v_b_26')
// (18, 11, 'sp4_v_b_15')
// (18, 12, 'sp4_h_l_40')
// (18, 12, 'sp4_h_r_9')
// (18, 12, 'sp4_v_b_2')
// (18, 17, 'sp4_h_l_40')
// (18, 17, 'sp4_h_r_5')
// (18, 18, 'sp4_h_r_38')
// (18, 20, 'sp4_h_r_12')
// (18, 20, 'sp4_h_r_35')
// (18, 21, 'sp4_h_r_42')
// (19, 0, 'fabout')
// (19, 0, 'local_g0_7')
// (19, 0, 'span4_horz_r_7')
// (19, 4, 'sp4_h_r_21')
// (19, 5, 'glb2local_0')
// (19, 5, 'local_g0_4')
// (19, 5, 'ram/RE')
// (19, 5, 'sp4_r_v_b_41')
// (19, 6, 'glb2local_0')
// (19, 6, 'local_g0_4')
// (19, 6, 'ram/WE')
// (19, 6, 'sp4_r_v_b_28')
// (19, 7, 'glb2local_0')
// (19, 7, 'glb2local_1')
// (19, 7, 'glb2local_2')
// (19, 7, 'local_g0_4')
// (19, 7, 'local_g0_5')
// (19, 7, 'local_g0_6')
// (19, 7, 'ram/MASK_10')
// (19, 7, 'ram/MASK_11')
// (19, 7, 'ram/MASK_12')
// (19, 7, 'ram/MASK_13')
// (19, 7, 'ram/MASK_14')
// (19, 7, 'ram/MASK_15')
// (19, 7, 'ram/MASK_8')
// (19, 7, 'ram/MASK_9')
// (19, 7, 'ram/RE')
// (19, 7, 'sp4_r_v_b_17')
// (19, 8, 'glb2local_0')
// (19, 8, 'glb2local_3')
// (19, 8, 'local_g0_4')
// (19, 8, 'local_g0_7')
// (19, 8, 'ram/MASK_4')
// (19, 8, 'ram/MASK_5')
// (19, 8, 'ram/MASK_6')
// (19, 8, 'ram/MASK_7')
// (19, 8, 'ram/WE')
// (19, 8, 'sp12_h_r_19')
// (19, 8, 'sp4_h_r_13')
// (19, 8, 'sp4_r_v_b_4')
// (19, 9, 'glb2local_0')
// (19, 9, 'glb2local_2')
// (19, 9, 'glb2local_3')
// (19, 9, 'local_g0_4')
// (19, 9, 'local_g0_6')
// (19, 9, 'local_g0_7')
// (19, 9, 'ram/MASK_10')
// (19, 9, 'ram/MASK_11')
// (19, 9, 'ram/MASK_12')
// (19, 9, 'ram/MASK_13')
// (19, 9, 'ram/MASK_14')
// (19, 9, 'ram/MASK_15')
// (19, 9, 'ram/MASK_8')
// (19, 9, 'ram/MASK_9')
// (19, 9, 'ram/RE')
// (19, 9, 'sp4_r_v_b_41')
// (19, 10, 'glb2local_0')
// (19, 10, 'glb2local_3')
// (19, 10, 'local_g0_4')
// (19, 10, 'local_g0_7')
// (19, 10, 'ram/MASK_4')
// (19, 10, 'ram/MASK_5')
// (19, 10, 'ram/MASK_6')
// (19, 10, 'ram/MASK_7')
// (19, 10, 'ram/WE')
// (19, 10, 'sp4_r_v_b_28')
// (19, 11, 'glb2local_0')
// (19, 11, 'local_g0_4')
// (19, 11, 'ram/RE')
// (19, 11, 'sp4_r_v_b_17')
// (19, 12, 'glb2local_0')
// (19, 12, 'local_g0_4')
// (19, 12, 'ram/WE')
// (19, 12, 'sp4_h_r_20')
// (19, 12, 'sp4_r_v_b_4')
// (19, 13, 'glb2local_0')
// (19, 13, 'local_g0_4')
// (19, 13, 'ram/RE')
// (19, 13, 'sp4_r_v_b_41')
// (19, 14, 'glb2local_0')
// (19, 14, 'local_g0_4')
// (19, 14, 'ram/WE')
// (19, 14, 'sp4_r_v_b_28')
// (19, 15, 'glb2local_0')
// (19, 15, 'local_g0_4')
// (19, 15, 'ram/RCLKE')
// (19, 15, 'ram/RE')
// (19, 15, 'sp4_r_v_b_17')
// (19, 16, 'glb2local_0')
// (19, 16, 'local_g0_4')
// (19, 16, 'ram/WE')
// (19, 16, 'sp4_r_v_b_4')
// (19, 17, 'sp4_h_r_16')
// (19, 17, 'sp4_r_v_b_36')
// (19, 18, 'sp4_h_l_38')
// (19, 18, 'sp4_h_r_3')
// (19, 18, 'sp4_r_v_b_25')
// (19, 19, 'sp4_r_v_b_12')
// (19, 20, 'sp4_h_r_25')
// (19, 20, 'sp4_h_r_46')
// (19, 20, 'sp4_r_v_b_1')
// (19, 21, 'sp4_h_l_42')
// (19, 21, 'sp4_h_r_4')
// (20, 0, 'span4_horz_r_11')
// (20, 4, 'sp4_h_r_32')
// (20, 4, 'sp4_v_t_41')
// (20, 5, 'sp4_v_b_41')
// (20, 6, 'sp4_v_b_28')
// (20, 7, 'glb2local_1')
// (20, 7, 'glb2local_2')
// (20, 7, 'local_g0_5')
// (20, 7, 'local_g0_6')
// (20, 7, 'local_g1_1')
// (20, 7, 'lutff_1/in_1')
// (20, 7, 'lutff_2/in_2')
// (20, 7, 'lutff_3/in_2')
// (20, 7, 'lutff_4/in_2')
// (20, 7, 'lutff_5/in_1')
// (20, 7, 'lutff_6/in_2')
// (20, 7, 'lutff_7/in_1')
// (20, 7, 'sp4_v_b_17')
// (20, 8, 'glb2local_2')
// (20, 8, 'glb2local_3')
// (20, 8, 'local_g0_6')
// (20, 8, 'local_g0_7')
// (20, 8, 'local_g3_0')
// (20, 8, 'lutff_0/in_1')
// (20, 8, 'lutff_1/in_2')
// (20, 8, 'lutff_2/in_1')
// (20, 8, 'lutff_3/in_1')
// (20, 8, 'sp12_h_r_20')
// (20, 8, 'sp4_h_r_24')
// (20, 8, 'sp4_v_b_4')
// (20, 8, 'sp4_v_t_41')
// (20, 9, 'sp4_v_b_41')
// (20, 10, 'sp4_v_b_28')
// (20, 11, 'sp4_v_b_17')
// (20, 12, 'sp4_h_r_33')
// (20, 12, 'sp4_v_b_4')
// (20, 12, 'sp4_v_t_41')
// (20, 13, 'sp4_v_b_41')
// (20, 14, 'glb2local_1')
// (20, 14, 'glb2local_2')
// (20, 14, 'local_g0_5')
// (20, 14, 'local_g0_6')
// (20, 14, 'lutff_1/in_2')
// (20, 14, 'lutff_2/in_2')
// (20, 14, 'sp4_v_b_28')
// (20, 15, 'sp4_v_b_17')
// (20, 16, 'sp4_v_b_4')
// (20, 16, 'sp4_v_t_36')
// (20, 17, 'sp4_h_r_29')
// (20, 17, 'sp4_v_b_36')
// (20, 18, 'sp4_h_r_14')
// (20, 18, 'sp4_v_b_25')
// (20, 19, 'sp4_v_b_12')
// (20, 20, 'sp4_h_l_46')
// (20, 20, 'sp4_h_r_36')
// (20, 20, 'sp4_h_r_8')
// (20, 20, 'sp4_v_b_1')
// (20, 21, 'sp4_h_r_17')
// (21, 0, 'span4_horz_r_15')
// (21, 1, 'sp4_r_v_b_43')
// (21, 2, 'sp4_r_v_b_30')
// (21, 3, 'glb2local_2')
// (21, 3, 'glb2local_3')
// (21, 3, 'local_g0_6')
// (21, 3, 'local_g0_7')
// (21, 3, 'lutff_1/in_2')
// (21, 3, 'lutff_2/in_2')
// (21, 3, 'lutff_3/in_2')
// (21, 3, 'lutff_4/in_2')
// (21, 3, 'lutff_5/in_2')
// (21, 3, 'lutff_6/in_1')
// (21, 3, 'lutff_7/in_1')
// (21, 3, 'sp4_r_v_b_19')
// (21, 4, 'glb2local_0')
// (21, 4, 'glb2local_1')
// (21, 4, 'local_g0_4')
// (21, 4, 'local_g0_5')
// (21, 4, 'lutff_0/in_2')
// (21, 4, 'lutff_1/in_1')
// (21, 4, 'lutff_2/in_1')
// (21, 4, 'lutff_3/in_1')
// (21, 4, 'lutff_4/in_2')
// (21, 4, 'lutff_5/in_1')
// (21, 4, 'lutff_6/in_1')
// (21, 4, 'lutff_7/in_1')
// (21, 4, 'sp4_h_r_45')
// (21, 4, 'sp4_r_v_b_6')
// (21, 5, 'glb2local_2')
// (21, 5, 'glb2local_3')
// (21, 5, 'local_g0_6')
// (21, 5, 'local_g0_7')
// (21, 5, 'lutff_0/in_2')
// (21, 5, 'lutff_1/in_2')
// (21, 5, 'lutff_2/in_2')
// (21, 5, 'lutff_3/in_2')
// (21, 5, 'lutff_4/in_1')
// (21, 5, 'lutff_5/in_2')
// (21, 5, 'lutff_6/in_0')
// (21, 5, 'sp4_r_v_b_39')
// (21, 5, 'sp4_r_v_b_43')
// (21, 5, 'sp4_r_v_b_44')
// (21, 6, 'sp4_r_v_b_26')
// (21, 6, 'sp4_r_v_b_30')
// (21, 6, 'sp4_r_v_b_33')
// (21, 7, 'local_g2_7')
// (21, 7, 'lutff_2/in_1')
// (21, 7, 'lutff_4/in_1')
// (21, 7, 'lutff_6/in_1')
// (21, 7, 'sp4_r_v_b_15')
// (21, 7, 'sp4_r_v_b_19')
// (21, 7, 'sp4_r_v_b_20')
// (21, 8, 'local_g2_1')
// (21, 8, 'lutff_0/in_1')
// (21, 8, 'lutff_2/in_1')
// (21, 8, 'sp12_h_r_23')
// (21, 8, 'sp4_h_r_37')
// (21, 8, 'sp4_r_v_b_2')
// (21, 8, 'sp4_r_v_b_6')
// (21, 8, 'sp4_r_v_b_9')
// (21, 9, 'sp4_r_v_b_43')
// (21, 10, 'sp4_r_v_b_30')
// (21, 11, 'sp4_r_v_b_19')
// (21, 12, 'sp4_h_r_44')
// (21, 12, 'sp4_r_v_b_6')
// (21, 13, 'glb2local_2')
// (21, 13, 'local_g0_6')
// (21, 13, 'lutff_7/in_1')
// (21, 13, 'sp4_r_v_b_37')
// (21, 13, 'sp4_r_v_b_38')
// (21, 14, 'sp4_r_v_b_24')
// (21, 14, 'sp4_r_v_b_27')
// (21, 15, 'sp4_r_v_b_13')
// (21, 15, 'sp4_r_v_b_14')
// (21, 16, 'sp4_r_v_b_0')
// (21, 16, 'sp4_r_v_b_3')
// (21, 17, 'sp4_h_r_40')
// (21, 17, 'sp4_r_v_b_37')
// (21, 18, 'sp4_h_r_27')
// (21, 18, 'sp4_r_v_b_24')
// (21, 18, 'sp4_r_v_b_40')
// (21, 19, 'neigh_op_tnr_0')
// (21, 19, 'sp4_r_v_b_13')
// (21, 19, 'sp4_r_v_b_29')
// (21, 20, 'neigh_op_rgt_0')
// (21, 20, 'sp4_h_l_36')
// (21, 20, 'sp4_h_r_21')
// (21, 20, 'sp4_h_r_5')
// (21, 20, 'sp4_r_v_b_0')
// (21, 20, 'sp4_r_v_b_16')
// (21, 21, 'neigh_op_bnr_0')
// (21, 21, 'sp4_h_r_28')
// (21, 21, 'sp4_r_v_b_5')
// (22, 0, 'span4_horz_l_15')
// (22, 0, 'span4_vert_43')
// (22, 1, 'sp4_v_b_43')
// (22, 2, 'sp4_r_v_b_45')
// (22, 2, 'sp4_v_b_30')
// (22, 3, 'sp4_r_v_b_32')
// (22, 3, 'sp4_v_b_19')
// (22, 4, 'sp4_h_l_45')
// (22, 4, 'sp4_r_v_b_21')
// (22, 4, 'sp4_v_b_6')
// (22, 4, 'sp4_v_t_39')
// (22, 4, 'sp4_v_t_43')
// (22, 4, 'sp4_v_t_44')
// (22, 5, 'sp4_r_v_b_8')
// (22, 5, 'sp4_v_b_39')
// (22, 5, 'sp4_v_b_43')
// (22, 5, 'sp4_v_b_44')
// (22, 6, 'sp4_r_v_b_37')
// (22, 6, 'sp4_v_b_26')
// (22, 6, 'sp4_v_b_30')
// (22, 6, 'sp4_v_b_33')
// (22, 7, 'sp4_r_v_b_24')
// (22, 7, 'sp4_v_b_15')
// (22, 7, 'sp4_v_b_19')
// (22, 7, 'sp4_v_b_20')
// (22, 8, 'sp12_h_l_23')
// (22, 8, 'sp12_v_t_23')
// (22, 8, 'sp4_h_l_37')
// (22, 8, 'sp4_r_v_b_13')
// (22, 8, 'sp4_v_b_2')
// (22, 8, 'sp4_v_b_6')
// (22, 8, 'sp4_v_b_9')
// (22, 8, 'sp4_v_t_43')
// (22, 9, 'sp12_v_b_23')
// (22, 9, 'sp4_r_v_b_0')
// (22, 9, 'sp4_v_b_43')
// (22, 10, 'sp12_v_b_20')
// (22, 10, 'sp4_r_v_b_37')
// (22, 10, 'sp4_v_b_30')
// (22, 11, 'sp12_v_b_19')
// (22, 11, 'sp4_r_v_b_24')
// (22, 11, 'sp4_v_b_19')
// (22, 12, 'sp12_v_b_16')
// (22, 12, 'sp4_h_l_44')
// (22, 12, 'sp4_r_v_b_13')
// (22, 12, 'sp4_v_b_6')
// (22, 12, 'sp4_v_t_37')
// (22, 12, 'sp4_v_t_38')
// (22, 13, 'sp12_v_b_15')
// (22, 13, 'sp4_r_v_b_0')
// (22, 13, 'sp4_v_b_37')
// (22, 13, 'sp4_v_b_38')
// (22, 14, 'glb2local_0')
// (22, 14, 'glb2local_3')
// (22, 14, 'local_g0_4')
// (22, 14, 'local_g0_7')
// (22, 14, 'local_g3_3')
// (22, 14, 'lutff_1/in_1')
// (22, 14, 'lutff_2/in_1')
// (22, 14, 'lutff_3/in_2')
// (22, 14, 'lutff_4/in_2')
// (22, 14, 'lutff_5/in_1')
// (22, 14, 'lutff_6/in_2')
// (22, 14, 'lutff_7/in_1')
// (22, 14, 'sp12_v_b_12')
// (22, 14, 'sp4_r_v_b_37')
// (22, 14, 'sp4_v_b_24')
// (22, 14, 'sp4_v_b_27')
// (22, 15, 'glb2local_0')
// (22, 15, 'glb2local_3')
// (22, 15, 'local_g0_4')
// (22, 15, 'local_g0_5')
// (22, 15, 'local_g0_7')
// (22, 15, 'lutff_0/in_2')
// (22, 15, 'lutff_1/in_2')
// (22, 15, 'lutff_2/in_2')
// (22, 15, 'lutff_3/in_2')
// (22, 15, 'lutff_4/in_2')
// (22, 15, 'sp12_v_b_11')
// (22, 15, 'sp4_r_v_b_24')
// (22, 15, 'sp4_v_b_13')
// (22, 15, 'sp4_v_b_14')
// (22, 16, 'sp12_v_b_8')
// (22, 16, 'sp4_r_v_b_13')
// (22, 16, 'sp4_v_b_0')
// (22, 16, 'sp4_v_b_3')
// (22, 16, 'sp4_v_t_37')
// (22, 17, 'sp12_v_b_7')
// (22, 17, 'sp4_h_l_40')
// (22, 17, 'sp4_r_v_b_0')
// (22, 17, 'sp4_v_b_37')
// (22, 17, 'sp4_v_t_40')
// (22, 18, 'sp12_v_b_4')
// (22, 18, 'sp4_h_r_38')
// (22, 18, 'sp4_r_v_b_41')
// (22, 18, 'sp4_v_b_24')
// (22, 18, 'sp4_v_b_40')
// (22, 19, 'neigh_op_top_0')
// (22, 19, 'sp12_v_b_3')
// (22, 19, 'sp4_r_v_b_28')
// (22, 19, 'sp4_r_v_b_44')
// (22, 19, 'sp4_v_b_13')
// (22, 19, 'sp4_v_b_29')
// (22, 20, 'lutff_0/out')
// (22, 20, 'sp12_v_b_0')
// (22, 20, 'sp4_h_r_16')
// (22, 20, 'sp4_h_r_32')
// (22, 20, 'sp4_r_v_b_17')
// (22, 20, 'sp4_r_v_b_33')
// (22, 20, 'sp4_v_b_0')
// (22, 20, 'sp4_v_b_16')
// (22, 21, 'neigh_op_bot_0')
// (22, 21, 'sp4_h_r_41')
// (22, 21, 'sp4_r_v_b_20')
// (22, 21, 'sp4_r_v_b_4')
// (22, 21, 'sp4_v_b_5')
// (22, 22, 'sp4_r_v_b_9')
// (23, 1, 'sp4_v_t_45')
// (23, 2, 'glb2local_0')
// (23, 2, 'glb2local_1')
// (23, 2, 'local_g0_4')
// (23, 2, 'local_g0_5')
// (23, 2, 'local_g2_5')
// (23, 2, 'lutff_1/in_1')
// (23, 2, 'lutff_2/in_2')
// (23, 2, 'lutff_3/in_2')
// (23, 2, 'lutff_4/in_1')
// (23, 2, 'lutff_5/in_2')
// (23, 2, 'lutff_6/in_1')
// (23, 2, 'lutff_7/in_2')
// (23, 2, 'sp4_v_b_45')
// (23, 3, 'glb2local_0')
// (23, 3, 'glb2local_1')
// (23, 3, 'local_g0_4')
// (23, 3, 'local_g0_5')
// (23, 3, 'local_g2_0')
// (23, 3, 'lutff_0/in_2')
// (23, 3, 'lutff_1/in_1')
// (23, 3, 'lutff_2/in_2')
// (23, 3, 'lutff_3/in_1')
// (23, 3, 'lutff_4/in_1')
// (23, 3, 'lutff_5/in_0')
// (23, 3, 'sp4_v_b_32')
// (23, 4, 'sp4_v_b_21')
// (23, 5, 'sp4_v_b_8')
// (23, 5, 'sp4_v_t_37')
// (23, 6, 'sp4_v_b_37')
// (23, 7, 'sp4_v_b_24')
// (23, 8, 'sp4_v_b_13')
// (23, 9, 'sp4_v_b_0')
// (23, 9, 'sp4_v_t_37')
// (23, 10, 'sp4_v_b_37')
// (23, 11, 'sp4_v_b_24')
// (23, 12, 'sp4_v_b_13')
// (23, 13, 'sp4_v_b_0')
// (23, 13, 'sp4_v_t_37')
// (23, 14, 'sp4_v_b_37')
// (23, 15, 'sp4_v_b_24')
// (23, 16, 'sp4_v_b_13')
// (23, 17, 'sp4_v_b_0')
// (23, 17, 'sp4_v_t_41')
// (23, 18, 'sp4_h_l_38')
// (23, 18, 'sp4_v_b_41')
// (23, 18, 'sp4_v_t_44')
// (23, 19, 'neigh_op_tnl_0')
// (23, 19, 'sp4_v_b_28')
// (23, 19, 'sp4_v_b_44')
// (23, 20, 'neigh_op_lft_0')
// (23, 20, 'sp4_h_r_29')
// (23, 20, 'sp4_h_r_45')
// (23, 20, 'sp4_v_b_17')
// (23, 20, 'sp4_v_b_33')
// (23, 21, 'neigh_op_bnl_0')
// (23, 21, 'sp4_h_l_41')
// (23, 21, 'sp4_v_b_20')
// (23, 21, 'sp4_v_b_4')
// (23, 22, 'sp4_v_b_9')
// (24, 3, 'glb2local_1')
// (24, 3, 'local_g0_5')
// (24, 3, 'lutff_0/in_3')
// (24, 20, 'sp4_h_l_45')
// (24, 20, 'sp4_h_r_40')
// (25, 20, 'sp4_h_l_40')

reg n9 = 0;
// (0, 1, 'neigh_op_tnr_1')
// (0, 2, 'neigh_op_rgt_1')
// (0, 3, 'neigh_op_bnr_1')
// (1, 1, 'neigh_op_top_1')
// (1, 2, 'lutff_1/out')
// (1, 3, 'local_g1_1')
// (1, 3, 'lutff_6/in_2')
// (1, 3, 'neigh_op_bot_1')
// (2, 1, 'neigh_op_tnl_1')
// (2, 2, 'neigh_op_lft_1')
// (2, 3, 'neigh_op_bnl_1')

reg n10 = 0;
// (0, 1, 'neigh_op_tnr_2')
// (0, 2, 'neigh_op_rgt_2')
// (0, 3, 'neigh_op_bnr_2')
// (1, 1, 'neigh_op_top_2')
// (1, 2, 'local_g3_2')
// (1, 2, 'lutff_2/out')
// (1, 2, 'lutff_6/in_3')
// (1, 3, 'local_g1_2')
// (1, 3, 'lutff_2/in_3')
// (1, 3, 'neigh_op_bot_2')
// (2, 1, 'neigh_op_tnl_2')
// (2, 2, 'neigh_op_lft_2')
// (2, 3, 'neigh_op_bnl_2')

reg n11 = 0;
// (0, 1, 'neigh_op_tnr_3')
// (0, 2, 'neigh_op_rgt_3')
// (0, 3, 'neigh_op_bnr_3')
// (1, 1, 'neigh_op_top_3')
// (1, 2, 'local_g1_3')
// (1, 2, 'lutff_3/out')
// (1, 2, 'lutff_7/in_3')
// (1, 3, 'local_g1_3')
// (1, 3, 'lutff_3/in_1')
// (1, 3, 'neigh_op_bot_3')
// (2, 1, 'neigh_op_tnl_3')
// (2, 2, 'neigh_op_lft_3')
// (2, 3, 'neigh_op_bnl_3')

reg n12 = 0;
// (0, 1, 'neigh_op_tnr_4')
// (0, 2, 'neigh_op_rgt_4')
// (0, 3, 'neigh_op_bnr_4')
// (1, 1, 'neigh_op_top_4')
// (1, 2, 'local_g2_4')
// (1, 2, 'lutff_1/in_3')
// (1, 2, 'lutff_4/out')
// (1, 3, 'local_g1_4')
// (1, 3, 'lutff_6/in_3')
// (1, 3, 'neigh_op_bot_4')
// (2, 1, 'neigh_op_tnl_4')
// (2, 2, 'neigh_op_lft_4')
// (2, 3, 'neigh_op_bnl_4')

reg n13 = 0;
// (0, 1, 'neigh_op_tnr_6')
// (0, 2, 'neigh_op_rgt_6')
// (0, 3, 'neigh_op_bnr_6')
// (1, 1, 'neigh_op_top_6')
// (1, 2, 'local_g2_6')
// (1, 2, 'lutff_4/in_2')
// (1, 2, 'lutff_6/out')
// (1, 3, 'local_g1_6')
// (1, 3, 'lutff_3/in_2')
// (1, 3, 'neigh_op_bot_6')
// (2, 1, 'neigh_op_tnl_6')
// (2, 2, 'neigh_op_lft_6')
// (2, 3, 'neigh_op_bnl_6')

reg n14 = 0;
// (0, 1, 'neigh_op_tnr_7')
// (0, 2, 'neigh_op_rgt_7')
// (0, 3, 'neigh_op_bnr_7')
// (1, 1, 'neigh_op_top_7')
// (1, 2, 'lutff_7/out')
// (1, 3, 'local_g0_7')
// (1, 3, 'lutff_5/in_2')
// (1, 3, 'lutff_7/in_2')
// (1, 3, 'neigh_op_bot_7')
// (2, 1, 'neigh_op_tnl_7')
// (2, 2, 'neigh_op_lft_7')
// (2, 3, 'neigh_op_bnl_7')

reg n15 = 0;
// (0, 1, 'sp4_h_r_4')
// (0, 1, 'sp4_h_r_7')
// (1, 1, 'sp4_h_r_17')
// (1, 1, 'sp4_h_r_18')
// (2, 1, 'local_g3_7')
// (2, 1, 'lutff_7/in_1')
// (2, 1, 'sp4_h_r_28')
// (2, 1, 'sp4_h_r_31')
// (3, 1, 'local_g2_1')
// (3, 1, 'lutff_5/in_0')
// (3, 1, 'sp4_h_r_41')
// (3, 1, 'sp4_h_r_42')
// (3, 2, 'sp4_r_v_b_39')
// (3, 3, 'local_g1_2')
// (3, 3, 'lutff_1/in_2')
// (3, 3, 'sp4_r_v_b_26')
// (3, 4, 'sp4_r_v_b_15')
// (3, 5, 'sp4_r_v_b_2')
// (3, 6, 'sp4_r_v_b_44')
// (3, 7, 'local_g0_2')
// (3, 7, 'lutff_6/in_0')
// (3, 7, 'sp4_r_v_b_33')
// (3, 8, 'sp4_r_v_b_20')
// (3, 9, 'sp4_r_v_b_9')
// (4, 1, 'sp4_h_l_41')
// (4, 1, 'sp4_h_l_42')
// (4, 1, 'sp4_h_r_4')
// (4, 1, 'sp4_v_t_39')
// (4, 2, 'sp4_h_r_6')
// (4, 2, 'sp4_v_b_39')
// (4, 3, 'sp4_v_b_26')
// (4, 4, 'sp4_v_b_15')
// (4, 5, 'sp4_h_r_9')
// (4, 5, 'sp4_r_v_b_45')
// (4, 5, 'sp4_v_b_2')
// (4, 5, 'sp4_v_t_44')
// (4, 6, 'sp4_r_v_b_32')
// (4, 6, 'sp4_v_b_44')
// (4, 7, 'sp4_r_v_b_21')
// (4, 7, 'sp4_v_b_33')
// (4, 8, 'sp4_r_v_b_8')
// (4, 8, 'sp4_v_b_20')
// (4, 9, 'sp4_r_v_b_39')
// (4, 9, 'sp4_v_b_9')
// (4, 10, 'local_g1_7')
// (4, 10, 'lutff_7/in_1')
// (4, 10, 'sp4_h_r_7')
// (4, 10, 'sp4_r_v_b_26')
// (4, 11, 'sp4_r_v_b_15')
// (4, 12, 'sp4_r_v_b_2')
// (4, 13, 'sp4_r_v_b_47')
// (4, 14, 'sp4_r_v_b_34')
// (4, 15, 'sp4_r_v_b_23')
// (4, 16, 'sp4_r_v_b_10')
// (4, 17, 'sp4_r_v_b_43')
// (4, 18, 'sp4_r_v_b_30')
// (4, 19, 'sp4_r_v_b_19')
// (4, 20, 'sp4_r_v_b_6')
// (5, 1, 'sp4_h_r_17')
// (5, 2, 'local_g0_3')
// (5, 2, 'lutff_6/in_3')
// (5, 2, 'sp4_h_r_19')
// (5, 4, 'sp4_v_t_45')
// (5, 5, 'local_g2_5')
// (5, 5, 'lutff_7/in_2')
// (5, 5, 'sp4_h_r_20')
// (5, 5, 'sp4_v_b_45')
// (5, 6, 'sp4_v_b_32')
// (5, 7, 'local_g1_5')
// (5, 7, 'lutff_4/in_2')
// (5, 7, 'sp4_v_b_21')
// (5, 8, 'sp4_h_r_8')
// (5, 8, 'sp4_v_b_8')
// (5, 8, 'sp4_v_t_39')
// (5, 9, 'sp4_v_b_39')
// (5, 10, 'sp4_h_r_18')
// (5, 10, 'sp4_v_b_26')
// (5, 11, 'sp4_v_b_15')
// (5, 12, 'sp4_v_b_2')
// (5, 12, 'sp4_v_t_47')
// (5, 13, 'sp4_v_b_47')
// (5, 14, 'sp4_v_b_34')
// (5, 15, 'sp4_v_b_23')
// (5, 16, 'sp4_v_b_10')
// (5, 16, 'sp4_v_t_43')
// (5, 17, 'sp4_v_b_43')
// (5, 18, 'sp4_v_b_30')
// (5, 19, 'sp4_v_b_19')
// (5, 20, 'local_g1_6')
// (5, 20, 'lutff_4/in_1')
// (5, 20, 'sp4_v_b_6')
// (6, 1, 'sp4_h_r_28')
// (6, 2, 'sp4_h_r_30')
// (6, 5, 'sp4_h_r_33')
// (6, 8, 'sp4_h_r_21')
// (6, 10, 'sp4_h_r_31')
// (7, 1, 'sp4_h_r_41')
// (7, 2, 'sp4_h_r_43')
// (7, 2, 'sp4_r_v_b_36')
// (7, 3, 'local_g0_1')
// (7, 3, 'lutff_0/in_1')
// (7, 3, 'sp4_r_v_b_25')
// (7, 4, 'sp4_r_v_b_12')
// (7, 5, 'sp4_h_r_44')
// (7, 5, 'sp4_r_v_b_1')
// (7, 8, 'sp4_h_r_32')
// (7, 10, 'sp4_h_r_42')
// (7, 11, 'sp4_r_v_b_36')
// (7, 12, 'sp4_r_v_b_25')
// (7, 13, 'sp4_r_v_b_12')
// (7, 14, 'sp4_r_v_b_1')
// (7, 15, 'sp4_r_v_b_44')
// (7, 16, 'sp4_r_v_b_33')
// (7, 17, 'sp4_r_v_b_20')
// (7, 18, 'sp4_r_v_b_9')
// (7, 19, 'sp4_r_v_b_40')
// (7, 20, 'sp4_r_v_b_29')
// (7, 21, 'local_g3_0')
// (7, 21, 'lutff_7/in_0')
// (7, 21, 'sp4_r_v_b_16')
// (7, 22, 'sp4_r_v_b_5')
// (8, 1, 'local_g0_2')
// (8, 1, 'lutff_0/in_2')
// (8, 1, 'sp4_h_l_41')
// (8, 1, 'sp4_h_r_10')
// (8, 1, 'sp4_h_r_4')
// (8, 1, 'sp4_v_t_36')
// (8, 2, 'local_g2_4')
// (8, 2, 'lutff_4/in_0')
// (8, 2, 'sp4_h_l_43')
// (8, 2, 'sp4_h_r_3')
// (8, 2, 'sp4_v_b_36')
// (8, 3, 'sp4_v_b_25')
// (8, 4, 'sp4_v_b_12')
// (8, 5, 'sp4_h_l_44')
// (8, 5, 'sp4_h_r_1')
// (8, 5, 'sp4_h_r_6')
// (8, 5, 'sp4_v_b_1')
// (8, 8, 'local_g3_5')
// (8, 8, 'lutff_1/in_3')
// (8, 8, 'sp4_h_r_45')
// (8, 9, 'sp4_r_v_b_37')
// (8, 10, 'sp4_h_l_42')
// (8, 10, 'sp4_h_r_7')
// (8, 10, 'sp4_r_v_b_24')
// (8, 10, 'sp4_v_t_36')
// (8, 11, 'sp4_r_v_b_13')
// (8, 11, 'sp4_v_b_36')
// (8, 12, 'local_g1_0')
// (8, 12, 'lutff_4/in_3')
// (8, 12, 'sp4_r_v_b_0')
// (8, 12, 'sp4_v_b_25')
// (8, 13, 'sp4_v_b_12')
// (8, 14, 'sp4_v_b_1')
// (8, 14, 'sp4_v_t_44')
// (8, 15, 'sp4_v_b_44')
// (8, 16, 'sp4_v_b_33')
// (8, 17, 'sp4_v_b_20')
// (8, 18, 'sp4_h_r_8')
// (8, 18, 'sp4_v_b_9')
// (8, 18, 'sp4_v_t_40')
// (8, 19, 'sp4_v_b_40')
// (8, 20, 'sp4_v_b_29')
// (8, 21, 'sp4_v_b_16')
// (8, 22, 'sp4_v_b_5')
// (9, 1, 'sp4_h_r_17')
// (9, 1, 'sp4_h_r_23')
// (9, 2, 'sp4_h_r_14')
// (9, 4, 'sp4_h_r_3')
// (9, 5, 'sp4_h_r_12')
// (9, 5, 'sp4_h_r_19')
// (9, 8, 'sp4_h_l_45')
// (9, 8, 'sp4_h_r_0')
// (9, 8, 'sp4_v_t_37')
// (9, 9, 'sp4_v_b_37')
// (9, 10, 'sp4_h_r_18')
// (9, 10, 'sp4_v_b_24')
// (9, 11, 'sp4_v_b_13')
// (9, 12, 'sp4_v_b_0')
// (9, 17, 'sp4_h_r_10')
// (9, 18, 'sp4_h_r_21')
// (9, 20, 'sp4_h_r_11')
// (10, 1, 'local_g2_2')
// (10, 1, 'lutff_2/in_2')
// (10, 1, 'sp4_h_r_28')
// (10, 1, 'sp4_h_r_34')
// (10, 1, 'sp4_r_v_b_47')
// (10, 2, 'sp4_h_r_27')
// (10, 2, 'sp4_r_v_b_34')
// (10, 3, 'local_g3_7')
// (10, 3, 'lutff_0/in_0')
// (10, 3, 'sp4_r_v_b_23')
// (10, 4, 'sp4_h_r_14')
// (10, 4, 'sp4_r_v_b_10')
// (10, 5, 'sp4_h_r_25')
// (10, 5, 'sp4_h_r_30')
// (10, 5, 'sp4_r_v_b_47')
// (10, 6, 'sp4_r_v_b_34')
// (10, 7, 'sp4_r_v_b_23')
// (10, 8, 'sp4_h_r_13')
// (10, 8, 'sp4_r_v_b_10')
// (10, 10, 'sp4_h_r_31')
// (10, 17, 'local_g0_7')
// (10, 17, 'lutff_4/in_1')
// (10, 17, 'sp4_h_r_23')
// (10, 18, 'local_g2_0')
// (10, 18, 'lutff_3/in_1')
// (10, 18, 'sp4_h_r_32')
// (10, 20, 'local_g0_6')
// (10, 20, 'lutff_1/in_1')
// (10, 20, 'sp4_h_r_22')
// (11, 0, 'span4_vert_47')
// (11, 1, 'sp4_h_r_41')
// (11, 1, 'sp4_h_r_47')
// (11, 1, 'sp4_v_b_47')
// (11, 2, 'sp4_h_r_38')
// (11, 2, 'sp4_r_v_b_47')
// (11, 2, 'sp4_v_b_34')
// (11, 3, 'sp4_r_v_b_34')
// (11, 3, 'sp4_v_b_23')
// (11, 4, 'local_g2_3')
// (11, 4, 'lutff_6/in_3')
// (11, 4, 'sp4_h_r_27')
// (11, 4, 'sp4_r_v_b_23')
// (11, 4, 'sp4_v_b_10')
// (11, 4, 'sp4_v_t_47')
// (11, 5, 'sp4_h_r_36')
// (11, 5, 'sp4_h_r_43')
// (11, 5, 'sp4_r_v_b_10')
// (11, 5, 'sp4_v_b_47')
// (11, 6, 'sp4_v_b_34')
// (11, 7, 'sp4_v_b_23')
// (11, 8, 'sp4_h_r_24')
// (11, 8, 'sp4_h_r_5')
// (11, 8, 'sp4_v_b_10')
// (11, 10, 'sp4_h_r_42')
// (11, 11, 'sp4_r_v_b_37')
// (11, 12, 'sp4_r_v_b_24')
// (11, 13, 'local_g2_5')
// (11, 13, 'lutff_7/in_2')
// (11, 13, 'sp4_r_v_b_13')
// (11, 14, 'sp4_r_v_b_0')
// (11, 15, 'sp4_r_v_b_45')
// (11, 16, 'sp4_r_v_b_32')
// (11, 17, 'local_g3_5')
// (11, 17, 'lutff_3/in_1')
// (11, 17, 'sp4_h_r_34')
// (11, 17, 'sp4_r_v_b_21')
// (11, 18, 'sp4_h_r_45')
// (11, 18, 'sp4_r_v_b_8')
// (11, 20, 'sp4_h_r_35')
// (12, 1, 'sp4_h_l_41')
// (12, 1, 'sp4_h_l_47')
// (12, 1, 'sp4_h_r_1')
// (12, 1, 'sp4_v_t_47')
// (12, 2, 'sp4_h_l_38')
// (12, 2, 'sp4_h_r_0')
// (12, 2, 'sp4_v_b_47')
// (12, 3, 'sp4_v_b_34')
// (12, 4, 'sp4_h_r_38')
// (12, 4, 'sp4_v_b_23')
// (12, 5, 'local_g0_3')
// (12, 5, 'lutff_4/in_1')
// (12, 5, 'sp4_h_l_36')
// (12, 5, 'sp4_h_l_43')
// (12, 5, 'sp4_h_r_10')
// (12, 5, 'sp4_h_r_3')
// (12, 5, 'sp4_v_b_10')
// (12, 8, 'local_g0_0')
// (12, 8, 'lutff_0/in_0')
// (12, 8, 'sp4_h_r_16')
// (12, 8, 'sp4_h_r_37')
// (12, 10, 'sp4_h_l_42')
// (12, 10, 'sp4_h_r_0')
// (12, 10, 'sp4_h_r_7')
// (12, 10, 'sp4_v_t_37')
// (12, 11, 'sp4_v_b_37')
// (12, 12, 'sp4_v_b_24')
// (12, 13, 'sp4_v_b_13')
// (12, 14, 'sp4_r_v_b_40')
// (12, 14, 'sp4_v_b_0')
// (12, 14, 'sp4_v_t_45')
// (12, 15, 'sp4_r_v_b_29')
// (12, 15, 'sp4_v_b_45')
// (12, 16, 'sp4_r_v_b_16')
// (12, 16, 'sp4_v_b_32')
// (12, 17, 'sp4_h_r_47')
// (12, 17, 'sp4_r_v_b_46')
// (12, 17, 'sp4_r_v_b_5')
// (12, 17, 'sp4_v_b_21')
// (12, 18, 'sp4_h_l_45')
// (12, 18, 'sp4_r_v_b_35')
// (12, 18, 'sp4_v_b_8')
// (12, 19, 'sp4_r_v_b_22')
// (12, 20, 'local_g2_3')
// (12, 20, 'lutff_4/in_1')
// (12, 20, 'sp4_h_r_46')
// (12, 20, 'sp4_r_v_b_11')
// (13, 1, 'sp4_h_r_12')
// (13, 2, 'sp4_h_r_13')
// (13, 4, 'local_g1_3')
// (13, 4, 'lutff_1/in_3')
// (13, 4, 'sp4_h_l_38')
// (13, 4, 'sp4_h_r_3')
// (13, 5, 'local_g1_7')
// (13, 5, 'lutff_7/in_3')
// (13, 5, 'sp4_h_r_14')
// (13, 5, 'sp4_h_r_23')
// (13, 8, 'sp4_h_l_37')
// (13, 8, 'sp4_h_r_29')
// (13, 8, 'sp4_h_r_9')
// (13, 10, 'sp4_h_r_13')
// (13, 10, 'sp4_h_r_18')
// (13, 13, 'sp4_h_r_11')
// (13, 13, 'sp4_v_t_40')
// (13, 14, 'sp4_v_b_40')
// (13, 15, 'sp4_v_b_29')
// (13, 16, 'sp4_h_r_11')
// (13, 16, 'sp4_v_b_16')
// (13, 16, 'sp4_v_t_46')
// (13, 17, 'sp4_h_l_47')
// (13, 17, 'sp4_v_b_46')
// (13, 17, 'sp4_v_b_5')
// (13, 18, 'sp4_v_b_35')
// (13, 19, 'sp4_v_b_22')
// (13, 20, 'sp4_h_l_46')
// (13, 20, 'sp4_v_b_11')
// (14, 1, 'local_g2_1')
// (14, 1, 'lutff_2/in_3')
// (14, 1, 'sp4_h_r_25')
// (14, 2, 'sp4_h_r_24')
// (14, 4, 'sp4_h_r_14')
// (14, 5, 'sp4_h_r_27')
// (14, 5, 'sp4_h_r_34')
// (14, 8, 'sp4_h_r_20')
// (14, 8, 'sp4_h_r_40')
// (14, 10, 'sp4_h_r_24')
// (14, 10, 'sp4_h_r_31')
// (14, 13, 'sp4_h_r_22')
// (14, 16, 'sp4_h_r_22')
// (15, 1, 'sp4_h_r_36')
// (15, 2, 'sp4_h_r_37')
// (15, 2, 'sp4_r_v_b_42')
// (15, 3, 'local_g0_7')
// (15, 3, 'lutff_4/in_1')
// (15, 3, 'sp4_r_v_b_31')
// (15, 4, 'sp4_h_r_27')
// (15, 4, 'sp4_r_v_b_18')
// (15, 5, 'sp4_h_r_38')
// (15, 5, 'sp4_h_r_47')
// (15, 5, 'sp4_r_v_b_7')
// (15, 8, 'sp4_h_l_40')
// (15, 8, 'sp4_h_r_33')
// (15, 8, 'sp4_h_r_9')
// (15, 10, 'sp4_h_r_37')
// (15, 10, 'sp4_h_r_42')
// (15, 13, 'sp4_h_r_35')
// (15, 16, 'sp4_h_r_35')
// (16, 1, 'sp4_h_l_36')
// (16, 1, 'sp4_h_r_1')
// (16, 1, 'sp4_v_t_42')
// (16, 2, 'local_g3_2')
// (16, 2, 'lutff_6/in_1')
// (16, 2, 'sp4_h_l_37')
// (16, 2, 'sp4_h_r_0')
// (16, 2, 'sp4_v_b_42')
// (16, 3, 'local_g3_7')
// (16, 3, 'lutff_0/in_0')
// (16, 3, 'sp4_v_b_31')
// (16, 4, 'sp4_h_r_38')
// (16, 4, 'sp4_v_b_18')
// (16, 5, 'local_g0_7')
// (16, 5, 'lutff_3/in_2')
// (16, 5, 'sp4_h_l_38')
// (16, 5, 'sp4_h_l_47')
// (16, 5, 'sp4_h_r_7')
// (16, 5, 'sp4_r_v_b_44')
// (16, 5, 'sp4_v_b_7')
// (16, 6, 'sp4_r_v_b_33')
// (16, 7, 'sp4_r_v_b_20')
// (16, 8, 'sp4_h_r_20')
// (16, 8, 'sp4_h_r_44')
// (16, 8, 'sp4_r_v_b_9')
// (16, 9, 'sp4_r_v_b_38')
// (16, 10, 'sp4_h_l_37')
// (16, 10, 'sp4_h_l_42')
// (16, 10, 'sp4_h_r_4')
// (16, 10, 'sp4_r_v_b_27')
// (16, 11, 'sp4_r_v_b_14')
// (16, 12, 'sp4_r_v_b_3')
// (16, 13, 'sp4_h_r_46')
// (16, 13, 'sp4_r_v_b_43')
// (16, 14, 'sp4_r_v_b_30')
// (16, 15, 'sp4_r_v_b_19')
// (16, 16, 'sp4_h_r_46')
// (16, 16, 'sp4_r_v_b_6')
// (17, 1, 'sp4_h_r_12')
// (17, 2, 'sp4_h_r_13')
// (17, 4, 'sp4_h_l_38')
// (17, 4, 'sp4_v_t_44')
// (17, 5, 'sp4_h_r_18')
// (17, 5, 'sp4_v_b_44')
// (17, 6, 'sp4_v_b_33')
// (17, 7, 'sp4_v_b_20')
// (17, 8, 'sp4_h_l_44')
// (17, 8, 'sp4_h_r_33')
// (17, 8, 'sp4_h_r_9')
// (17, 8, 'sp4_v_b_9')
// (17, 8, 'sp4_v_t_38')
// (17, 9, 'sp4_v_b_38')
// (17, 10, 'sp4_h_r_17')
// (17, 10, 'sp4_v_b_27')
// (17, 11, 'sp4_v_b_14')
// (17, 12, 'sp4_v_b_3')
// (17, 12, 'sp4_v_t_43')
// (17, 13, 'sp4_h_l_46')
// (17, 13, 'sp4_h_r_8')
// (17, 13, 'sp4_v_b_43')
// (17, 14, 'sp4_v_b_30')
// (17, 15, 'sp4_v_b_19')
// (17, 16, 'sp4_h_l_46')
// (17, 16, 'sp4_v_b_6')
// (18, 1, 'sp4_h_r_25')
// (18, 2, 'sp4_h_r_24')
// (18, 5, 'sp4_h_r_31')
// (18, 8, 'sp4_h_r_20')
// (18, 8, 'sp4_h_r_44')
// (18, 10, 'sp4_h_r_28')
// (18, 13, 'sp4_h_r_21')
// (19, 1, 'sp4_h_r_36')
// (19, 2, 'sp4_h_r_37')
// (19, 2, 'sp4_r_v_b_36')
// (19, 3, 'sp4_r_v_b_25')
// (19, 3, 'sp4_r_v_b_37')
// (19, 4, 'sp4_r_v_b_12')
// (19, 4, 'sp4_r_v_b_24')
// (19, 5, 'sp4_h_r_42')
// (19, 5, 'sp4_r_v_b_1')
// (19, 5, 'sp4_r_v_b_13')
// (19, 6, 'sp4_r_v_b_0')
// (19, 6, 'sp4_r_v_b_36')
// (19, 7, 'neigh_op_tnr_6')
// (19, 7, 'sp4_r_v_b_25')
// (19, 7, 'sp4_r_v_b_41')
// (19, 8, 'neigh_op_rgt_6')
// (19, 8, 'sp4_h_l_44')
// (19, 8, 'sp4_h_r_1')
// (19, 8, 'sp4_h_r_33')
// (19, 8, 'sp4_r_v_b_12')
// (19, 8, 'sp4_r_v_b_28')
// (19, 9, 'neigh_op_bnr_6')
// (19, 9, 'sp4_r_v_b_1')
// (19, 9, 'sp4_r_v_b_17')
// (19, 10, 'sp4_h_r_41')
// (19, 10, 'sp4_r_v_b_4')
// (19, 13, 'sp4_h_r_32')
// (20, 1, 'sp4_h_l_36')
// (20, 1, 'sp4_v_t_36')
// (20, 2, 'sp4_h_l_37')
// (20, 2, 'sp4_v_b_36')
// (20, 2, 'sp4_v_t_37')
// (20, 3, 'sp4_v_b_25')
// (20, 3, 'sp4_v_b_37')
// (20, 4, 'sp4_v_b_12')
// (20, 4, 'sp4_v_b_24')
// (20, 5, 'sp4_h_l_42')
// (20, 5, 'sp4_v_b_1')
// (20, 5, 'sp4_v_b_13')
// (20, 5, 'sp4_v_t_36')
// (20, 6, 'sp4_r_v_b_37')
// (20, 6, 'sp4_v_b_0')
// (20, 6, 'sp4_v_b_36')
// (20, 6, 'sp4_v_t_41')
// (20, 7, 'neigh_op_top_6')
// (20, 7, 'sp4_r_v_b_24')
// (20, 7, 'sp4_v_b_25')
// (20, 7, 'sp4_v_b_41')
// (20, 8, 'lutff_6/out')
// (20, 8, 'sp4_h_r_12')
// (20, 8, 'sp4_h_r_44')
// (20, 8, 'sp4_r_v_b_13')
// (20, 8, 'sp4_v_b_12')
// (20, 8, 'sp4_v_b_28')
// (20, 9, 'neigh_op_bot_6')
// (20, 9, 'sp4_r_v_b_0')
// (20, 9, 'sp4_v_b_1')
// (20, 9, 'sp4_v_b_17')
// (20, 10, 'sp4_h_l_41')
// (20, 10, 'sp4_r_v_b_45')
// (20, 10, 'sp4_v_b_4')
// (20, 11, 'sp4_r_v_b_32')
// (20, 12, 'sp4_r_v_b_21')
// (20, 13, 'sp4_h_r_45')
// (20, 13, 'sp4_r_v_b_8')
// (21, 5, 'sp4_v_t_37')
// (21, 6, 'sp4_v_b_37')
// (21, 7, 'neigh_op_tnl_6')
// (21, 7, 'sp4_v_b_24')
// (21, 8, 'neigh_op_lft_6')
// (21, 8, 'sp4_h_l_44')
// (21, 8, 'sp4_h_r_25')
// (21, 8, 'sp4_v_b_13')
// (21, 9, 'neigh_op_bnl_6')
// (21, 9, 'sp4_v_b_0')
// (21, 9, 'sp4_v_t_45')
// (21, 10, 'sp4_v_b_45')
// (21, 11, 'sp4_v_b_32')
// (21, 12, 'sp4_v_b_21')
// (21, 13, 'sp4_h_l_45')
// (21, 13, 'sp4_v_b_8')
// (22, 8, 'sp4_h_r_36')
// (23, 8, 'sp4_h_l_36')

reg n16 = 0;
// (0, 1, 'sp4_r_v_b_27')
// (0, 2, 'sp4_r_v_b_14')
// (0, 3, 'sp4_r_v_b_3')
// (0, 4, 'sp4_r_v_b_38')
// (0, 5, 'neigh_op_tnr_7')
// (0, 5, 'sp4_r_v_b_27')
// (0, 6, 'neigh_op_rgt_7')
// (0, 6, 'sp4_r_v_b_14')
// (0, 7, 'neigh_op_bnr_7')
// (0, 7, 'sp4_r_v_b_3')
// (1, 0, 'span4_vert_27')
// (1, 1, 'sp4_v_b_27')
// (1, 2, 'local_g0_6')
// (1, 2, 'lutff_3/in_3')
// (1, 2, 'sp4_v_b_14')
// (1, 3, 'sp4_v_b_3')
// (1, 3, 'sp4_v_t_38')
// (1, 4, 'local_g2_6')
// (1, 4, 'lutff_1/in_1')
// (1, 4, 'sp4_v_b_38')
// (1, 5, 'neigh_op_top_7')
// (1, 5, 'sp4_v_b_27')
// (1, 6, 'lutff_7/out')
// (1, 6, 'sp4_v_b_14')
// (1, 7, 'neigh_op_bot_7')
// (1, 7, 'sp4_v_b_3')
// (2, 5, 'neigh_op_tnl_7')
// (2, 6, 'neigh_op_lft_7')
// (2, 7, 'neigh_op_bnl_7')

wire n17;
// (0, 1, 'sp4_r_v_b_31')
// (0, 2, 'sp4_r_v_b_18')
// (0, 3, 'sp4_h_r_14')
// (0, 3, 'sp4_r_v_b_7')
// (0, 4, 'sp4_r_v_b_46')
// (0, 5, 'sp4_r_v_b_35')
// (0, 6, 'sp4_r_v_b_22')
// (0, 7, 'sp4_r_v_b_11')
// (0, 8, 'sp4_r_v_b_45')
// (0, 9, 'sp4_r_v_b_32')
// (0, 10, 'sp4_r_v_b_21')
// (0, 11, 'sp4_r_v_b_8')
// (1, 0, 'span4_vert_31')
// (1, 1, 'sp4_v_b_31')
// (1, 2, 'local_g0_2')
// (1, 2, 'lutff_global/cen')
// (1, 2, 'sp4_v_b_18')
// (1, 3, 'local_g3_3')
// (1, 3, 'lutff_global/cen')
// (1, 3, 'sp4_h_r_27')
// (1, 3, 'sp4_v_b_7')
// (1, 3, 'sp4_v_t_46')
// (1, 4, 'sp4_r_v_b_43')
// (1, 4, 'sp4_v_b_46')
// (1, 5, 'sp4_r_v_b_30')
// (1, 5, 'sp4_v_b_35')
// (1, 6, 'local_g3_3')
// (1, 6, 'lutff_global/cen')
// (1, 6, 'sp4_r_v_b_19')
// (1, 6, 'sp4_v_b_22')
// (1, 7, 'sp4_r_v_b_6')
// (1, 7, 'sp4_v_b_11')
// (1, 7, 'sp4_v_t_45')
// (1, 8, 'sp4_r_v_b_47')
// (1, 8, 'sp4_v_b_45')
// (1, 9, 'sp4_r_v_b_34')
// (1, 9, 'sp4_v_b_32')
// (1, 10, 'sp4_r_v_b_23')
// (1, 10, 'sp4_v_b_21')
// (1, 11, 'sp4_h_r_8')
// (1, 11, 'sp4_r_v_b_10')
// (1, 11, 'sp4_v_b_8')
// (2, 1, 'sp4_r_v_b_27')
// (2, 2, 'sp4_r_v_b_14')
// (2, 3, 'local_g1_3')
// (2, 3, 'lutff_global/cen')
// (2, 3, 'sp4_h_r_38')
// (2, 3, 'sp4_r_v_b_3')
// (2, 3, 'sp4_v_t_43')
// (2, 4, 'sp4_r_v_b_38')
// (2, 4, 'sp4_v_b_43')
// (2, 5, 'sp4_r_v_b_27')
// (2, 5, 'sp4_v_b_30')
// (2, 6, 'sp4_r_v_b_14')
// (2, 6, 'sp4_v_b_19')
// (2, 7, 'sp4_r_v_b_3')
// (2, 7, 'sp4_v_b_6')
// (2, 7, 'sp4_v_t_47')
// (2, 8, 'sp4_r_v_b_37')
// (2, 8, 'sp4_v_b_47')
// (2, 9, 'sp4_r_v_b_24')
// (2, 9, 'sp4_v_b_34')
// (2, 10, 'neigh_op_tnr_0')
// (2, 10, 'sp4_r_v_b_13')
// (2, 10, 'sp4_v_b_23')
// (2, 11, 'neigh_op_rgt_0')
// (2, 11, 'sp4_h_r_21')
// (2, 11, 'sp4_h_r_5')
// (2, 11, 'sp4_r_v_b_0')
// (2, 11, 'sp4_v_b_10')
// (2, 12, 'neigh_op_bnr_0')
// (3, 0, 'span4_vert_27')
// (3, 1, 'sp4_v_b_27')
// (3, 2, 'sp4_v_b_14')
// (3, 3, 'sp4_h_l_38')
// (3, 3, 'sp4_v_b_3')
// (3, 3, 'sp4_v_t_38')
// (3, 4, 'sp4_v_b_38')
// (3, 5, 'sp4_v_b_27')
// (3, 6, 'sp4_v_b_14')
// (3, 7, 'sp4_v_b_3')
// (3, 7, 'sp4_v_t_37')
// (3, 8, 'sp4_v_b_37')
// (3, 9, 'sp4_v_b_24')
// (3, 10, 'neigh_op_top_0')
// (3, 10, 'sp4_v_b_13')
// (3, 11, 'local_g1_0')
// (3, 11, 'lutff_0/out')
// (3, 11, 'lutff_6/in_1')
// (3, 11, 'sp4_h_r_16')
// (3, 11, 'sp4_h_r_32')
// (3, 11, 'sp4_v_b_0')
// (3, 12, 'neigh_op_bot_0')
// (4, 10, 'neigh_op_tnl_0')
// (4, 11, 'neigh_op_lft_0')
// (4, 11, 'sp4_h_r_29')
// (4, 11, 'sp4_h_r_45')
// (4, 12, 'neigh_op_bnl_0')
// (5, 11, 'sp4_h_l_45')
// (5, 11, 'sp4_h_r_40')
// (6, 11, 'sp4_h_l_40')

reg n18 = 0;
// (0, 2, 'neigh_op_tnr_0')
// (0, 3, 'neigh_op_rgt_0')
// (0, 4, 'neigh_op_bnr_0')
// (1, 2, 'neigh_op_top_0')
// (1, 3, 'local_g0_0')
// (1, 3, 'lutff_0/out')
// (1, 3, 'lutff_4/in_2')
// (1, 3, 'lutff_5/in_1')
// (1, 4, 'neigh_op_bot_0')
// (2, 2, 'neigh_op_tnl_0')
// (2, 3, 'neigh_op_lft_0')
// (2, 4, 'neigh_op_bnl_0')

wire n19;
// (0, 2, 'neigh_op_tnr_1')
// (0, 3, 'neigh_op_rgt_1')
// (0, 4, 'neigh_op_bnr_1')
// (1, 2, 'neigh_op_top_1')
// (1, 3, 'lutff_1/out')
// (1, 4, 'neigh_op_bot_1')
// (2, 2, 'neigh_op_tnl_1')
// (2, 3, 'local_g0_1')
// (2, 3, 'lutff_3/in_0')
// (2, 3, 'neigh_op_lft_1')
// (2, 4, 'neigh_op_bnl_1')

wire n20;
// (0, 2, 'neigh_op_tnr_2')
// (0, 3, 'neigh_op_rgt_2')
// (0, 4, 'neigh_op_bnr_2')
// (1, 2, 'neigh_op_top_2')
// (1, 3, 'lutff_2/out')
// (1, 4, 'neigh_op_bot_2')
// (2, 2, 'neigh_op_tnl_2')
// (2, 3, 'local_g1_2')
// (2, 3, 'lutff_3/in_2')
// (2, 3, 'neigh_op_lft_2')
// (2, 4, 'neigh_op_bnl_2')

wire n21;
// (0, 2, 'neigh_op_tnr_3')
// (0, 3, 'neigh_op_rgt_3')
// (0, 4, 'neigh_op_bnr_3')
// (1, 2, 'neigh_op_top_3')
// (1, 3, 'local_g2_3')
// (1, 3, 'lutff_1/in_0')
// (1, 3, 'lutff_3/out')
// (1, 4, 'neigh_op_bot_3')
// (2, 2, 'neigh_op_tnl_3')
// (2, 3, 'neigh_op_lft_3')
// (2, 4, 'neigh_op_bnl_3')

reg n22 = 0;
// (0, 2, 'neigh_op_tnr_4')
// (0, 3, 'neigh_op_rgt_4')
// (0, 4, 'neigh_op_bnr_4')
// (1, 2, 'local_g1_4')
// (1, 2, 'lutff_2/in_1')
// (1, 2, 'neigh_op_top_4')
// (1, 3, 'lutff_4/out')
// (1, 4, 'neigh_op_bot_4')
// (2, 2, 'neigh_op_tnl_4')
// (2, 3, 'neigh_op_lft_4')
// (2, 4, 'local_g3_4')
// (2, 4, 'lutff_2/in_3')
// (2, 4, 'neigh_op_bnl_4')

wire n23;
// (0, 2, 'neigh_op_tnr_5')
// (0, 3, 'neigh_op_rgt_5')
// (0, 4, 'neigh_op_bnr_5')
// (1, 2, 'neigh_op_top_5')
// (1, 3, 'local_g2_5')
// (1, 3, 'lutff_1/in_2')
// (1, 3, 'lutff_5/out')
// (1, 4, 'neigh_op_bot_5')
// (2, 2, 'neigh_op_tnl_5')
// (2, 3, 'neigh_op_lft_5')
// (2, 4, 'neigh_op_bnl_5')

wire n24;
// (0, 2, 'neigh_op_tnr_6')
// (0, 3, 'neigh_op_rgt_6')
// (0, 4, 'neigh_op_bnr_6')
// (1, 2, 'neigh_op_top_6')
// (1, 3, 'local_g0_6')
// (1, 3, 'lutff_1/in_3')
// (1, 3, 'lutff_6/out')
// (1, 4, 'neigh_op_bot_6')
// (2, 2, 'neigh_op_tnl_6')
// (2, 3, 'neigh_op_lft_6')
// (2, 4, 'neigh_op_bnl_6')

reg n25 = 0;
// (0, 2, 'neigh_op_tnr_7')
// (0, 3, 'neigh_op_rgt_7')
// (0, 4, 'neigh_op_bnr_7')
// (1, 2, 'neigh_op_top_7')
// (1, 3, 'lutff_7/out')
// (1, 4, 'local_g0_7')
// (1, 4, 'lutff_1/in_0')
// (1, 4, 'neigh_op_bot_7')
// (2, 2, 'neigh_op_tnl_7')
// (2, 3, 'local_g0_7')
// (2, 3, 'lutff_4/in_3')
// (2, 3, 'neigh_op_lft_7')
// (2, 4, 'neigh_op_bnl_7')

reg n26 = 0;
// (0, 2, 'sp4_r_v_b_45')
// (0, 3, 'sp4_r_v_b_32')
// (0, 4, 'neigh_op_tnr_4')
// (0, 4, 'sp4_r_v_b_21')
// (0, 5, 'neigh_op_rgt_4')
// (0, 5, 'sp4_r_v_b_8')
// (0, 6, 'neigh_op_bnr_4')
// (1, 1, 'sp4_v_t_45')
// (1, 2, 'sp4_v_b_45')
// (1, 3, 'local_g2_0')
// (1, 3, 'lutff_3/in_3')
// (1, 3, 'sp4_v_b_32')
// (1, 4, 'neigh_op_top_4')
// (1, 4, 'sp4_v_b_21')
// (1, 5, 'local_g0_4')
// (1, 5, 'lutff_4/out')
// (1, 5, 'lutff_7/in_1')
// (1, 5, 'sp4_v_b_8')
// (1, 6, 'neigh_op_bot_4')
// (2, 4, 'neigh_op_tnl_4')
// (2, 5, 'neigh_op_lft_4')
// (2, 6, 'local_g3_4')
// (2, 6, 'lutff_6/in_1')
// (2, 6, 'neigh_op_bnl_4')

reg n27 = 0;
// (0, 3, 'neigh_op_tnr_0')
// (0, 4, 'neigh_op_rgt_0')
// (0, 5, 'neigh_op_bnr_0')
// (1, 3, 'local_g1_0')
// (1, 3, 'lutff_3/in_0')
// (1, 3, 'neigh_op_top_0')
// (1, 4, 'local_g2_0')
// (1, 4, 'lutff_0/out')
// (1, 4, 'lutff_2/in_0')
// (1, 4, 'lutff_5/in_3')
// (1, 5, 'neigh_op_bot_0')
// (2, 3, 'neigh_op_tnl_0')
// (2, 4, 'neigh_op_lft_0')
// (2, 5, 'neigh_op_bnl_0')

wire n28;
// (0, 3, 'neigh_op_tnr_1')
// (0, 4, 'neigh_op_rgt_1')
// (0, 5, 'neigh_op_bnr_1')
// (1, 3, 'neigh_op_top_1')
// (1, 4, 'lutff_1/out')
// (1, 5, 'neigh_op_bot_1')
// (2, 3, 'local_g3_1')
// (2, 3, 'lutff_3/in_3')
// (2, 3, 'neigh_op_tnl_1')
// (2, 4, 'neigh_op_lft_1')
// (2, 5, 'neigh_op_bnl_1')

reg n29 = 0;
// (0, 3, 'neigh_op_tnr_2')
// (0, 4, 'neigh_op_rgt_2')
// (0, 5, 'neigh_op_bnr_2')
// (1, 3, 'local_g0_2')
// (1, 3, 'lutff_6/in_0')
// (1, 3, 'neigh_op_top_2')
// (1, 4, 'local_g3_2')
// (1, 4, 'lutff_2/out')
// (1, 4, 'lutff_3/in_0')
// (1, 4, 'lutff_5/in_0')
// (1, 5, 'neigh_op_bot_2')
// (2, 3, 'neigh_op_tnl_2')
// (2, 4, 'neigh_op_lft_2')
// (2, 5, 'neigh_op_bnl_2')

reg n30 = 0;
// (0, 3, 'neigh_op_tnr_3')
// (0, 4, 'neigh_op_rgt_3')
// (0, 5, 'neigh_op_bnr_3')
// (1, 3, 'local_g0_3')
// (1, 3, 'lutff_6/in_1')
// (1, 3, 'neigh_op_top_3')
// (1, 4, 'local_g1_3')
// (1, 4, 'lutff_3/out')
// (1, 4, 'lutff_4/in_2')
// (1, 5, 'local_g0_3')
// (1, 5, 'lutff_3/in_2')
// (1, 5, 'neigh_op_bot_3')
// (2, 3, 'neigh_op_tnl_3')
// (2, 4, 'neigh_op_lft_3')
// (2, 5, 'neigh_op_bnl_3')

wire n31;
// (0, 3, 'neigh_op_tnr_4')
// (0, 4, 'neigh_op_rgt_4')
// (0, 5, 'neigh_op_bnr_4')
// (1, 3, 'neigh_op_top_4')
// (1, 4, 'lutff_4/out')
// (1, 5, 'neigh_op_bot_4')
// (2, 3, 'neigh_op_tnl_4')
// (2, 4, 'local_g1_4')
// (2, 4, 'lutff_5/in_0')
// (2, 4, 'neigh_op_lft_4')
// (2, 5, 'neigh_op_bnl_4')

wire n32;
// (0, 3, 'neigh_op_tnr_5')
// (0, 4, 'neigh_op_rgt_5')
// (0, 5, 'neigh_op_bnr_5')
// (1, 3, 'neigh_op_top_5')
// (1, 4, 'lutff_5/out')
// (1, 5, 'neigh_op_bot_5')
// (2, 3, 'neigh_op_tnl_5')
// (2, 4, 'local_g0_5')
// (2, 4, 'lutff_5/in_2')
// (2, 4, 'neigh_op_lft_5')
// (2, 5, 'neigh_op_bnl_5')

reg n33 = 0;
// (0, 3, 'neigh_op_tnr_6')
// (0, 4, 'neigh_op_rgt_6')
// (0, 5, 'neigh_op_bnr_6')
// (1, 3, 'neigh_op_top_6')
// (1, 4, 'local_g3_6')
// (1, 4, 'lutff_1/in_2')
// (1, 4, 'lutff_6/out')
// (1, 5, 'neigh_op_bot_6')
// (2, 3, 'neigh_op_tnl_6')
// (2, 4, 'local_g1_6')
// (2, 4, 'lutff_4/in_3')
// (2, 4, 'lutff_7/in_0')
// (2, 4, 'neigh_op_lft_6')
// (2, 5, 'neigh_op_bnl_6')

reg n34 = 0;
// (0, 3, 'neigh_op_tnr_7')
// (0, 4, 'neigh_op_rgt_7')
// (0, 5, 'neigh_op_bnr_7')
// (1, 3, 'local_g1_7')
// (1, 3, 'lutff_2/in_2')
// (1, 3, 'neigh_op_top_7')
// (1, 4, 'local_g3_7')
// (1, 4, 'lutff_0/in_0')
// (1, 4, 'lutff_4/in_0')
// (1, 4, 'lutff_7/out')
// (1, 5, 'neigh_op_bot_7')
// (2, 3, 'neigh_op_tnl_7')
// (2, 4, 'neigh_op_lft_7')
// (2, 5, 'neigh_op_bnl_7')

reg n35 = 0;
// (0, 3, 'sp4_h_r_28')
// (1, 3, 'local_g3_1')
// (1, 3, 'lutff_5/in_3')
// (1, 3, 'sp4_h_r_41')
// (1, 4, 'neigh_op_tnr_6')
// (1, 4, 'sp4_r_v_b_41')
// (1, 5, 'local_g2_6')
// (1, 5, 'lutff_0/in_2')
// (1, 5, 'neigh_op_rgt_6')
// (1, 5, 'sp4_r_v_b_28')
// (1, 6, 'neigh_op_bnr_6')
// (1, 6, 'sp4_r_v_b_17')
// (1, 7, 'sp4_r_v_b_4')
// (2, 3, 'sp4_h_l_41')
// (2, 3, 'sp4_v_t_41')
// (2, 4, 'neigh_op_top_6')
// (2, 4, 'sp4_v_b_41')
// (2, 5, 'local_g2_6')
// (2, 5, 'lutff_5/in_1')
// (2, 5, 'lutff_6/out')
// (2, 5, 'sp4_v_b_28')
// (2, 6, 'neigh_op_bot_6')
// (2, 6, 'sp4_v_b_17')
// (2, 7, 'sp4_v_b_4')
// (3, 4, 'neigh_op_tnl_6')
// (3, 5, 'neigh_op_lft_6')
// (3, 6, 'neigh_op_bnl_6')

reg n36 = 0;
// (0, 4, 'neigh_op_tnr_0')
// (0, 5, 'neigh_op_rgt_0')
// (0, 6, 'neigh_op_bnr_0')
// (1, 4, 'local_g0_0')
// (1, 4, 'lutff_7/in_1')
// (1, 4, 'neigh_op_top_0')
// (1, 5, 'lutff_0/out')
// (1, 6, 'neigh_op_bot_0')
// (2, 4, 'local_g3_0')
// (2, 4, 'lutff_2/in_1')
// (2, 4, 'neigh_op_tnl_0')
// (2, 5, 'local_g1_0')
// (2, 5, 'lutff_3/in_0')
// (2, 5, 'neigh_op_lft_0')
// (2, 6, 'neigh_op_bnl_0')

wire n37;
// (0, 4, 'neigh_op_tnr_3')
// (0, 5, 'neigh_op_rgt_3')
// (0, 6, 'neigh_op_bnr_3')
// (1, 4, 'local_g0_3')
// (1, 4, 'lutff_3/in_2')
// (1, 4, 'lutff_6/in_1')
// (1, 4, 'neigh_op_top_3')
// (1, 5, 'local_g2_3')
// (1, 5, 'lutff_0/in_3')
// (1, 5, 'lutff_3/out')
// (1, 5, 'lutff_5/in_0')
// (1, 6, 'neigh_op_bot_3')
// (2, 4, 'local_g2_3')
// (2, 4, 'lutff_3/in_2')
// (2, 4, 'lutff_4/in_1')
// (2, 4, 'lutff_6/in_3')
// (2, 4, 'neigh_op_tnl_3')
// (2, 5, 'neigh_op_lft_3')
// (2, 6, 'neigh_op_bnl_3')

reg n38 = 0;
// (0, 4, 'neigh_op_tnr_5')
// (0, 5, 'neigh_op_rgt_5')
// (0, 6, 'neigh_op_bnr_5')
// (1, 4, 'local_g1_5')
// (1, 4, 'lutff_1/in_3')
// (1, 4, 'neigh_op_top_5')
// (1, 5, 'local_g0_5')
// (1, 5, 'lutff_4/in_1')
// (1, 5, 'lutff_5/out')
// (1, 5, 'lutff_6/in_3')
// (1, 6, 'neigh_op_bot_5')
// (2, 4, 'neigh_op_tnl_5')
// (2, 5, 'neigh_op_lft_5')
// (2, 6, 'neigh_op_bnl_5')

wire n39;
// (0, 4, 'neigh_op_tnr_6')
// (0, 5, 'neigh_op_rgt_6')
// (0, 6, 'neigh_op_bnr_6')
// (1, 4, 'neigh_op_top_6')
// (1, 5, 'lutff_6/out')
// (1, 6, 'neigh_op_bot_6')
// (2, 4, 'neigh_op_tnl_6')
// (2, 5, 'neigh_op_lft_6')
// (2, 6, 'local_g3_6')
// (2, 6, 'lutff_6/in_3')
// (2, 6, 'neigh_op_bnl_6')

reg n40 = 0;
// (0, 4, 'neigh_op_tnr_7')
// (0, 5, 'neigh_op_rgt_7')
// (0, 6, 'neigh_op_bnr_7')
// (1, 3, 'local_g2_7')
// (1, 3, 'lutff_5/in_0')
// (1, 3, 'sp4_r_v_b_39')
// (1, 4, 'local_g1_7')
// (1, 4, 'lutff_6/in_0')
// (1, 4, 'neigh_op_top_7')
// (1, 4, 'sp4_r_v_b_26')
// (1, 5, 'local_g1_7')
// (1, 5, 'lutff_6/in_0')
// (1, 5, 'lutff_7/out')
// (1, 5, 'sp4_r_v_b_15')
// (1, 6, 'neigh_op_bot_7')
// (1, 6, 'sp4_r_v_b_2')
// (2, 2, 'sp4_v_t_39')
// (2, 3, 'sp4_v_b_39')
// (2, 4, 'neigh_op_tnl_7')
// (2, 4, 'sp4_v_b_26')
// (2, 5, 'neigh_op_lft_7')
// (2, 5, 'sp4_v_b_15')
// (2, 6, 'neigh_op_bnl_7')
// (2, 6, 'sp4_v_b_2')

reg n41 = 0;
// (0, 4, 'sp4_h_r_30')
// (0, 5, 'sp4_h_r_30')
// (1, 1, 'sp4_r_v_b_38')
// (1, 2, 'sp4_r_v_b_27')
// (1, 3, 'sp4_r_v_b_14')
// (1, 4, 'local_g2_3')
// (1, 4, 'lutff_4/in_3')
// (1, 4, 'lutff_5/in_2')
// (1, 4, 'sp4_h_r_43')
// (1, 4, 'sp4_r_v_b_3')
// (1, 5, 'local_g3_3')
// (1, 5, 'lutff_6/in_2')
// (1, 5, 'sp4_h_r_43')
// (1, 5, 'sp4_r_v_b_44')
// (1, 6, 'sp4_r_v_b_33')
// (1, 7, 'sp4_h_r_8')
// (1, 7, 'sp4_r_v_b_20')
// (1, 8, 'sp4_r_v_b_9')
// (2, 0, 'span4_vert_38')
// (2, 1, 'local_g2_6')
// (2, 1, 'lutff_4/in_0')
// (2, 1, 'lutff_6/in_0')
// (2, 1, 'sp4_h_r_10')
// (2, 1, 'sp4_v_b_38')
// (2, 2, 'local_g3_3')
// (2, 2, 'lutff_5/in_3')
// (2, 2, 'sp4_v_b_27')
// (2, 3, 'sp4_v_b_14')
// (2, 4, 'local_g1_3')
// (2, 4, 'lutff_7/in_1')
// (2, 4, 'sp4_h_l_43')
// (2, 4, 'sp4_h_r_3')
// (2, 4, 'sp4_v_b_3')
// (2, 4, 'sp4_v_t_44')
// (2, 5, 'local_g0_3')
// (2, 5, 'lutff_3/in_2')
// (2, 5, 'lutff_5/in_2')
// (2, 5, 'lutff_7/in_0')
// (2, 5, 'sp4_h_l_43')
// (2, 5, 'sp4_h_r_3')
// (2, 5, 'sp4_v_b_44')
// (2, 6, 'local_g2_1')
// (2, 6, 'lutff_1/in_2')
// (2, 6, 'sp4_v_b_33')
// (2, 7, 'local_g1_5')
// (2, 7, 'lutff_1/in_3')
// (2, 7, 'sp4_h_r_21')
// (2, 7, 'sp4_v_b_20')
// (2, 8, 'sp4_v_b_9')
// (3, 1, 'local_g0_7')
// (3, 1, 'lutff_0/in_1')
// (3, 1, 'lutff_2/in_1')
// (3, 1, 'sp4_h_r_23')
// (3, 1, 'sp4_r_v_b_41')
// (3, 2, 'local_g0_4')
// (3, 2, 'lutff_2/in_0')
// (3, 2, 'lutff_4/in_2')
// (3, 2, 'sp4_r_v_b_28')
// (3, 3, 'sp4_r_v_b_17')
// (3, 4, 'local_g0_6')
// (3, 4, 'lutff_5/in_1')
// (3, 4, 'lutff_7/in_3')
// (3, 4, 'sp4_h_r_14')
// (3, 4, 'sp4_r_v_b_4')
// (3, 5, 'local_g1_6')
// (3, 5, 'lutff_1/in_0')
// (3, 5, 'lutff_6/in_1')
// (3, 5, 'sp4_h_r_14')
// (3, 5, 'sp4_r_v_b_46')
// (3, 6, 'local_g0_0')
// (3, 6, 'local_g2_3')
// (3, 6, 'lutff_1/in_2')
// (3, 6, 'lutff_2/in_1')
// (3, 6, 'lutff_7/in_1')
// (3, 6, 'sp4_r_v_b_35')
// (3, 7, 'local_g3_6')
// (3, 7, 'lutff_4/in_1')
// (3, 7, 'sp4_h_r_32')
// (3, 7, 'sp4_r_v_b_22')
// (3, 8, 'sp4_r_v_b_11')
// (4, 0, 'span4_vert_41')
// (4, 1, 'local_g3_3')
// (4, 1, 'lutff_2/in_2')
// (4, 1, 'lutff_3/in_3')
// (4, 1, 'lutff_6/in_0')
// (4, 1, 'sp4_h_r_34')
// (4, 1, 'sp4_r_v_b_43')
// (4, 1, 'sp4_v_b_41')
// (4, 2, 'local_g0_6')
// (4, 2, 'lutff_3/in_3')
// (4, 2, 'lutff_4/in_2')
// (4, 2, 'sp4_r_v_b_30')
// (4, 2, 'sp4_v_b_28')
// (4, 3, 'local_g2_3')
// (4, 3, 'local_g3_3')
// (4, 3, 'lutff_1/in_1')
// (4, 3, 'lutff_7/in_2')
// (4, 3, 'neigh_op_tnr_3')
// (4, 3, 'sp4_r_v_b_19')
// (4, 3, 'sp4_v_b_17')
// (4, 4, 'local_g3_3')
// (4, 4, 'lutff_1/in_1')
// (4, 4, 'lutff_3/in_3')
// (4, 4, 'neigh_op_rgt_3')
// (4, 4, 'sp4_h_r_11')
// (4, 4, 'sp4_h_r_27')
// (4, 4, 'sp4_r_v_b_38')
// (4, 4, 'sp4_r_v_b_6')
// (4, 4, 'sp4_v_b_4')
// (4, 4, 'sp4_v_t_46')
// (4, 5, 'local_g0_3')
// (4, 5, 'lutff_6/in_1')
// (4, 5, 'neigh_op_bnr_3')
// (4, 5, 'sp4_h_r_27')
// (4, 5, 'sp4_r_v_b_27')
// (4, 5, 'sp4_v_b_46')
// (4, 6, 'local_g2_6')
// (4, 6, 'lutff_0/in_2')
// (4, 6, 'sp4_r_v_b_14')
// (4, 6, 'sp4_v_b_35')
// (4, 7, 'local_g1_3')
// (4, 7, 'lutff_3/in_3')
// (4, 7, 'lutff_7/in_3')
// (4, 7, 'sp4_h_r_45')
// (4, 7, 'sp4_r_v_b_3')
// (4, 7, 'sp4_v_b_22')
// (4, 8, 'sp4_v_b_11')
// (5, 0, 'span4_vert_43')
// (5, 1, 'local_g2_3')
// (5, 1, 'lutff_0/in_3')
// (5, 1, 'lutff_7/in_2')
// (5, 1, 'sp4_h_r_47')
// (5, 1, 'sp4_v_b_43')
// (5, 2, 'local_g2_6')
// (5, 2, 'lutff_0/in_2')
// (5, 2, 'sp4_r_v_b_47')
// (5, 2, 'sp4_v_b_30')
// (5, 3, 'local_g0_3')
// (5, 3, 'lutff_4/in_1')
// (5, 3, 'lutff_5/in_0')
// (5, 3, 'lutff_7/in_2')
// (5, 3, 'neigh_op_top_3')
// (5, 3, 'sp4_r_v_b_34')
// (5, 3, 'sp4_v_b_19')
// (5, 3, 'sp4_v_t_38')
// (5, 4, 'local_g1_3')
// (5, 4, 'local_g2_3')
// (5, 4, 'lutff_1/in_0')
// (5, 4, 'lutff_3/in_2')
// (5, 4, 'lutff_3/out')
// (5, 4, 'lutff_4/in_2')
// (5, 4, 'lutff_6/in_0')
// (5, 4, 'lutff_7/in_2')
// (5, 4, 'sp4_h_r_22')
// (5, 4, 'sp4_h_r_38')
// (5, 4, 'sp4_h_r_6')
// (5, 4, 'sp4_r_v_b_23')
// (5, 4, 'sp4_r_v_b_39')
// (5, 4, 'sp4_v_b_38')
// (5, 4, 'sp4_v_b_6')
// (5, 5, 'local_g1_3')
// (5, 5, 'lutff_0/in_2')
// (5, 5, 'lutff_1/in_1')
// (5, 5, 'lutff_5/in_3')
// (5, 5, 'neigh_op_bot_3')
// (5, 5, 'sp4_h_r_38')
// (5, 5, 'sp4_r_v_b_10')
// (5, 5, 'sp4_r_v_b_26')
// (5, 5, 'sp4_v_b_27')
// (5, 6, 'local_g2_7')
// (5, 6, 'lutff_4/in_1')
// (5, 6, 'lutff_7/in_0')
// (5, 6, 'sp4_r_v_b_15')
// (5, 6, 'sp4_v_b_14')
// (5, 7, 'local_g0_3')
// (5, 7, 'lutff_5/in_2')
// (5, 7, 'sp4_h_l_45')
// (5, 7, 'sp4_r_v_b_2')
// (5, 7, 'sp4_v_b_3')
// (6, 1, 'sp4_h_l_47')
// (6, 1, 'sp4_h_r_10')
// (6, 1, 'sp4_v_t_47')
// (6, 2, 'sp4_v_b_47')
// (6, 3, 'neigh_op_tnl_3')
// (6, 3, 'sp4_h_r_7')
// (6, 3, 'sp4_v_b_34')
// (6, 3, 'sp4_v_t_39')
// (6, 4, 'neigh_op_lft_3')
// (6, 4, 'sp4_h_l_38')
// (6, 4, 'sp4_h_r_19')
// (6, 4, 'sp4_h_r_35')
// (6, 4, 'sp4_v_b_23')
// (6, 4, 'sp4_v_b_39')
// (6, 5, 'neigh_op_bnl_3')
// (6, 5, 'sp4_h_l_38')
// (6, 5, 'sp4_v_b_10')
// (6, 5, 'sp4_v_b_26')
// (6, 6, 'sp4_v_b_15')
// (6, 7, 'sp4_v_b_2')
// (7, 1, 'local_g0_7')
// (7, 1, 'local_g1_7')
// (7, 1, 'lutff_1/in_3')
// (7, 1, 'lutff_2/in_1')
// (7, 1, 'sp4_h_r_23')
// (7, 1, 'sp4_r_v_b_40')
// (7, 2, 'sp4_r_v_b_29')
// (7, 3, 'sp4_h_r_18')
// (7, 3, 'sp4_r_v_b_16')
// (7, 4, 'sp4_h_r_30')
// (7, 4, 'sp4_h_r_46')
// (7, 4, 'sp4_r_v_b_5')
// (8, 0, 'span4_vert_40')
// (8, 1, 'local_g3_2')
// (8, 1, 'lutff_1/in_2')
// (8, 1, 'lutff_6/in_3')
// (8, 1, 'sp4_h_r_34')
// (8, 1, 'sp4_r_v_b_43')
// (8, 1, 'sp4_v_b_40')
// (8, 2, 'local_g3_5')
// (8, 2, 'lutff_5/in_3')
// (8, 2, 'sp4_r_v_b_30')
// (8, 2, 'sp4_v_b_29')
// (8, 3, 'sp4_h_r_31')
// (8, 3, 'sp4_r_v_b_19')
// (8, 3, 'sp4_v_b_16')
// (8, 4, 'sp4_h_l_46')
// (8, 4, 'sp4_h_r_11')
// (8, 4, 'sp4_h_r_43')
// (8, 4, 'sp4_h_r_7')
// (8, 4, 'sp4_r_v_b_6')
// (8, 4, 'sp4_v_b_5')
// (9, 0, 'span4_vert_43')
// (9, 1, 'local_g2_7')
// (9, 1, 'lutff_1/in_0')
// (9, 1, 'lutff_4/in_3')
// (9, 1, 'sp4_h_r_47')
// (9, 1, 'sp4_r_v_b_31')
// (9, 1, 'sp4_v_b_43')
// (9, 2, 'local_g2_6')
// (9, 2, 'lutff_3/in_1')
// (9, 2, 'lutff_5/in_3')
// (9, 2, 'lutff_6/in_0')
// (9, 2, 'sp4_r_v_b_18')
// (9, 2, 'sp4_v_b_30')
// (9, 3, 'local_g1_3')
// (9, 3, 'lutff_5/in_3')
// (9, 3, 'sp4_h_r_42')
// (9, 3, 'sp4_r_v_b_7')
// (9, 3, 'sp4_v_b_19')
// (9, 4, 'local_g1_2')
// (9, 4, 'lutff_5/in_2')
// (9, 4, 'lutff_7/in_0')
// (9, 4, 'sp4_h_l_43')
// (9, 4, 'sp4_h_r_18')
// (9, 4, 'sp4_h_r_2')
// (9, 4, 'sp4_h_r_22')
// (9, 4, 'sp4_v_b_6')
// (10, 0, 'span4_vert_31')
// (10, 1, 'local_g0_6')
// (10, 1, 'lutff_0/in_0')
// (10, 1, 'lutff_4/in_0')
// (10, 1, 'lutff_6/in_0')
// (10, 1, 'sp4_h_l_47')
// (10, 1, 'sp4_h_r_6')
// (10, 1, 'sp4_v_b_31')
// (10, 2, 'local_g0_2')
// (10, 2, 'local_g1_2')
// (10, 2, 'lutff_2/in_0')
// (10, 2, 'lutff_6/in_3')
// (10, 2, 'sp4_v_b_18')
// (10, 3, 'local_g1_3')
// (10, 3, 'lutff_1/in_3')
// (10, 3, 'lutff_4/in_0')
// (10, 3, 'sp4_h_l_42')
// (10, 3, 'sp4_h_r_3')
// (10, 3, 'sp4_v_b_7')
// (10, 4, 'local_g3_7')
// (10, 4, 'lutff_4/in_2')
// (10, 4, 'sp4_h_r_15')
// (10, 4, 'sp4_h_r_31')
// (10, 4, 'sp4_h_r_35')
// (11, 1, 'sp4_h_r_19')
// (11, 1, 'sp4_r_v_b_40')
// (11, 2, 'local_g1_5')
// (11, 2, 'lutff_3/in_3')
// (11, 2, 'sp4_r_v_b_29')
// (11, 3, 'sp4_h_r_14')
// (11, 3, 'sp4_r_v_b_16')
// (11, 4, 'sp4_h_r_26')
// (11, 4, 'sp4_h_r_42')
// (11, 4, 'sp4_h_r_46')
// (11, 4, 'sp4_r_v_b_5')
// (12, 0, 'span4_vert_40')
// (12, 1, 'sp4_h_r_30')
// (12, 1, 'sp4_v_b_40')
// (12, 2, 'sp4_v_b_29')
// (12, 3, 'sp4_h_r_27')
// (12, 3, 'sp4_v_b_16')
// (12, 4, 'sp4_h_l_42')
// (12, 4, 'sp4_h_l_46')
// (12, 4, 'sp4_h_r_39')
// (12, 4, 'sp4_v_b_5')
// (13, 1, 'sp4_h_r_43')
// (13, 3, 'sp4_h_r_38')
// (13, 4, 'sp4_h_l_39')
// (14, 1, 'sp4_h_l_43')
// (14, 3, 'sp4_h_l_38')

wire n42;
// (0, 4, 'sp4_r_v_b_44')
// (0, 5, 'sp4_r_v_b_33')
// (0, 5, 'sp4_r_v_b_42')
// (0, 6, 'sp4_r_v_b_20')
// (0, 6, 'sp4_r_v_b_31')
// (0, 7, 'sp4_r_v_b_18')
// (0, 7, 'sp4_r_v_b_9')
// (0, 8, 'sp4_r_v_b_43')
// (0, 8, 'sp4_r_v_b_7')
// (0, 9, 'sp4_r_v_b_30')
// (0, 9, 'sp4_r_v_b_46')
// (0, 10, 'neigh_op_tnr_3')
// (0, 10, 'sp4_r_v_b_19')
// (0, 10, 'sp4_r_v_b_35')
// (0, 11, 'neigh_op_rgt_3')
// (0, 11, 'sp4_r_v_b_22')
// (0, 11, 'sp4_r_v_b_6')
// (0, 12, 'neigh_op_bnr_3')
// (0, 12, 'sp4_r_v_b_11')
// (1, 3, 'sp4_v_t_44')
// (1, 4, 'local_g2_4')
// (1, 4, 'lutff_global/s_r')
// (1, 4, 'sp4_h_r_0')
// (1, 4, 'sp4_v_b_44')
// (1, 4, 'sp4_v_t_42')
// (1, 5, 'local_g2_4')
// (1, 5, 'lutff_global/s_r')
// (1, 5, 'sp4_r_v_b_36')
// (1, 5, 'sp4_v_b_33')
// (1, 5, 'sp4_v_b_42')
// (1, 6, 'sp4_r_v_b_25')
// (1, 6, 'sp4_v_b_20')
// (1, 6, 'sp4_v_b_31')
// (1, 7, 'sp4_r_v_b_12')
// (1, 7, 'sp4_v_b_18')
// (1, 7, 'sp4_v_b_9')
// (1, 7, 'sp4_v_t_43')
// (1, 8, 'sp4_r_v_b_1')
// (1, 8, 'sp4_v_b_43')
// (1, 8, 'sp4_v_b_7')
// (1, 8, 'sp4_v_t_46')
// (1, 9, 'sp4_r_v_b_47')
// (1, 9, 'sp4_v_b_30')
// (1, 9, 'sp4_v_b_46')
// (1, 10, 'neigh_op_top_3')
// (1, 10, 'sp4_r_v_b_34')
// (1, 10, 'sp4_v_b_19')
// (1, 10, 'sp4_v_b_35')
// (1, 11, 'lutff_3/out')
// (1, 11, 'sp4_r_v_b_23')
// (1, 11, 'sp4_v_b_22')
// (1, 11, 'sp4_v_b_6')
// (1, 12, 'neigh_op_bot_3')
// (1, 12, 'sp4_r_v_b_10')
// (1, 12, 'sp4_v_b_11')
// (2, 4, 'local_g1_5')
// (2, 4, 'lutff_global/s_r')
// (2, 4, 'sp4_h_r_13')
// (2, 4, 'sp4_v_t_36')
// (2, 5, 'local_g2_4')
// (2, 5, 'lutff_global/s_r')
// (2, 5, 'sp4_v_b_36')
// (2, 6, 'sp4_v_b_25')
// (2, 7, 'sp4_v_b_12')
// (2, 8, 'sp4_v_b_1')
// (2, 8, 'sp4_v_t_47')
// (2, 9, 'sp4_v_b_47')
// (2, 10, 'local_g3_3')
// (2, 10, 'lutff_1/in_3')
// (2, 10, 'neigh_op_tnl_3')
// (2, 10, 'sp4_v_b_34')
// (2, 11, 'local_g1_3')
// (2, 11, 'lutff_0/in_0')
// (2, 11, 'neigh_op_lft_3')
// (2, 11, 'sp4_v_b_23')
// (2, 12, 'neigh_op_bnl_3')
// (2, 12, 'sp4_v_b_10')
// (3, 4, 'sp4_h_r_24')
// (4, 4, 'sp4_h_r_37')
// (5, 4, 'sp4_h_l_37')

wire n43;
// (0, 5, 'neigh_op_tnr_5')
// (0, 6, 'neigh_op_rgt_5')
// (0, 7, 'neigh_op_bnr_5')
// (1, 5, 'neigh_op_top_5')
// (1, 5, 'sp4_r_v_b_38')
// (1, 6, 'lutff_5/out')
// (1, 6, 'sp4_r_v_b_27')
// (1, 7, 'neigh_op_bot_5')
// (1, 7, 'sp4_r_v_b_14')
// (1, 8, 'sp4_r_v_b_3')
// (2, 4, 'sp4_v_t_38')
// (2, 5, 'neigh_op_tnl_5')
// (2, 5, 'sp4_v_b_38')
// (2, 6, 'neigh_op_lft_5')
// (2, 6, 'sp4_v_b_27')
// (2, 7, 'neigh_op_bnl_5')
// (2, 7, 'sp4_v_b_14')
// (2, 8, 'sp4_h_r_3')
// (2, 8, 'sp4_v_b_3')
// (3, 8, 'local_g0_6')
// (3, 8, 'local_g1_6')
// (3, 8, 'lutff_3/in_0')
// (3, 8, 'lutff_4/in_1')
// (3, 8, 'lutff_5/in_3')
// (3, 8, 'lutff_7/in_1')
// (3, 8, 'sp4_h_r_14')
// (4, 8, 'sp4_h_r_27')
// (5, 8, 'sp4_h_r_38')
// (6, 8, 'sp4_h_l_38')

reg n44 = 0;
// (0, 5, 'sp4_h_r_5')
// (1, 5, 'sp4_h_r_16')
// (2, 5, 'local_g3_5')
// (2, 5, 'lutff_7/in_1')
// (2, 5, 'sp4_h_r_29')
// (2, 6, 'neigh_op_tnr_6')
// (2, 7, 'neigh_op_rgt_6')
// (2, 8, 'neigh_op_bnr_6')
// (3, 5, 'sp4_h_r_40')
// (3, 6, 'neigh_op_top_6')
// (3, 6, 'sp4_r_v_b_40')
// (3, 7, 'lutff_6/out')
// (3, 7, 'sp4_r_v_b_29')
// (3, 8, 'neigh_op_bot_6')
// (3, 8, 'sp4_r_v_b_16')
// (3, 9, 'sp4_r_v_b_5')
// (4, 5, 'sp4_h_l_40')
// (4, 5, 'sp4_v_t_40')
// (4, 6, 'neigh_op_tnl_6')
// (4, 6, 'sp4_v_b_40')
// (4, 7, 'local_g0_6')
// (4, 7, 'lutff_3/in_1')
// (4, 7, 'neigh_op_lft_6')
// (4, 7, 'sp4_v_b_29')
// (4, 8, 'local_g2_6')
// (4, 8, 'local_g3_6')
// (4, 8, 'lutff_3/in_0')
// (4, 8, 'lutff_5/in_0')
// (4, 8, 'lutff_6/in_3')
// (4, 8, 'lutff_7/in_1')
// (4, 8, 'neigh_op_bnl_6')
// (4, 8, 'sp4_v_b_16')
// (4, 9, 'sp4_v_b_5')

reg n45 = 0;
// (0, 5, 'sp4_h_r_7')
// (1, 5, 'local_g1_2')
// (1, 5, 'lutff_3/in_0')
// (1, 5, 'sp4_h_r_18')
// (1, 5, 'sp4_r_v_b_46')
// (1, 6, 'local_g0_0')
// (1, 6, 'lutff_7/in_1')
// (1, 6, 'sp4_r_v_b_35')
// (1, 7, 'sp4_r_v_b_22')
// (1, 8, 'sp4_r_v_b_11')
// (1, 9, 'sp4_r_v_b_46')
// (1, 10, 'sp4_r_v_b_35')
// (1, 11, 'local_g3_6')
// (1, 11, 'lutff_6/in_3')
// (1, 11, 'lutff_7/in_0')
// (1, 11, 'sp4_r_v_b_22')
// (1, 12, 'sp4_r_v_b_11')
// (1, 13, 'sp4_r_v_b_40')
// (1, 13, 'sp4_r_v_b_46')
// (1, 14, 'local_g0_0')
// (1, 14, 'lutff_7/in_1')
// (1, 14, 'sp4_r_v_b_29')
// (1, 14, 'sp4_r_v_b_35')
// (1, 15, 'sp4_r_v_b_16')
// (1, 15, 'sp4_r_v_b_22')
// (1, 16, 'sp4_r_v_b_11')
// (1, 16, 'sp4_r_v_b_5')
// (1, 17, 'sp4_r_v_b_36')
// (1, 18, 'sp4_r_v_b_25')
// (1, 19, 'sp4_r_v_b_12')
// (1, 20, 'sp4_r_v_b_1')
// (2, 4, 'sp4_v_t_46')
// (2, 5, 'sp4_h_r_31')
// (2, 5, 'sp4_v_b_46')
// (2, 6, 'sp4_v_b_35')
// (2, 7, 'sp4_v_b_22')
// (2, 8, 'sp4_v_b_11')
// (2, 8, 'sp4_v_t_46')
// (2, 9, 'sp4_v_b_46')
// (2, 10, 'sp4_v_b_35')
// (2, 11, 'neigh_op_tnr_3')
// (2, 11, 'sp4_v_b_22')
// (2, 12, 'neigh_op_rgt_3')
// (2, 12, 'sp4_h_r_11')
// (2, 12, 'sp4_r_v_b_38')
// (2, 12, 'sp4_v_b_11')
// (2, 12, 'sp4_v_t_40')
// (2, 12, 'sp4_v_t_46')
// (2, 13, 'local_g1_3')
// (2, 13, 'lutff_7/in_1')
// (2, 13, 'neigh_op_bnr_3')
// (2, 13, 'sp4_r_v_b_27')
// (2, 13, 'sp4_r_v_b_37')
// (2, 13, 'sp4_v_b_40')
// (2, 13, 'sp4_v_b_46')
// (2, 14, 'local_g2_6')
// (2, 14, 'lutff_0/in_2')
// (2, 14, 'sp4_r_v_b_14')
// (2, 14, 'sp4_r_v_b_24')
// (2, 14, 'sp4_v_b_29')
// (2, 14, 'sp4_v_b_35')
// (2, 15, 'sp4_r_v_b_13')
// (2, 15, 'sp4_r_v_b_3')
// (2, 15, 'sp4_v_b_16')
// (2, 15, 'sp4_v_b_22')
// (2, 16, 'sp4_r_v_b_0')
// (2, 16, 'sp4_r_v_b_46')
// (2, 16, 'sp4_v_b_11')
// (2, 16, 'sp4_v_b_5')
// (2, 16, 'sp4_v_t_36')
// (2, 17, 'sp4_r_v_b_35')
// (2, 17, 'sp4_v_b_36')
// (2, 18, 'sp4_r_v_b_22')
// (2, 18, 'sp4_v_b_25')
// (2, 19, 'local_g2_3')
// (2, 19, 'lutff_4/in_3')
// (2, 19, 'sp4_r_v_b_11')
// (2, 19, 'sp4_v_b_12')
// (2, 20, 'local_g0_1')
// (2, 20, 'lutff_2/in_1')
// (2, 20, 'sp4_v_b_1')
// (3, 5, 'sp4_h_r_42')
// (3, 6, 'sp4_r_v_b_36')
// (3, 7, 'sp4_r_v_b_25')
// (3, 8, 'sp4_r_v_b_12')
// (3, 9, 'sp4_r_v_b_1')
// (3, 9, 'sp4_r_v_b_42')
// (3, 10, 'local_g0_7')
// (3, 10, 'lutff_4/in_3')
// (3, 10, 'sp4_r_v_b_31')
// (3, 10, 'sp4_r_v_b_47')
// (3, 11, 'neigh_op_top_3')
// (3, 11, 'sp12_v_t_22')
// (3, 11, 'sp4_r_v_b_18')
// (3, 11, 'sp4_r_v_b_34')
// (3, 11, 'sp4_v_t_38')
// (3, 12, 'lutff_3/out')
// (3, 12, 'sp12_v_b_22')
// (3, 12, 'sp4_h_r_22')
// (3, 12, 'sp4_h_r_6')
// (3, 12, 'sp4_r_v_b_23')
// (3, 12, 'sp4_r_v_b_39')
// (3, 12, 'sp4_r_v_b_7')
// (3, 12, 'sp4_v_b_38')
// (3, 12, 'sp4_v_t_37')
// (3, 13, 'neigh_op_bot_3')
// (3, 13, 'sp12_v_b_21')
// (3, 13, 'sp4_r_v_b_10')
// (3, 13, 'sp4_r_v_b_26')
// (3, 13, 'sp4_v_b_27')
// (3, 13, 'sp4_v_b_37')
// (3, 14, 'sp12_v_b_18')
// (3, 14, 'sp4_r_v_b_15')
// (3, 14, 'sp4_v_b_14')
// (3, 14, 'sp4_v_b_24')
// (3, 15, 'sp12_v_b_17')
// (3, 15, 'sp4_r_v_b_2')
// (3, 15, 'sp4_v_b_13')
// (3, 15, 'sp4_v_b_3')
// (3, 15, 'sp4_v_t_46')
// (3, 16, 'local_g0_0')
// (3, 16, 'lutff_2/in_0')
// (3, 16, 'sp12_v_b_14')
// (3, 16, 'sp4_v_b_0')
// (3, 16, 'sp4_v_b_46')
// (3, 17, 'sp12_v_b_13')
// (3, 17, 'sp4_v_b_35')
// (3, 18, 'sp12_v_b_10')
// (3, 18, 'sp4_v_b_22')
// (3, 19, 'sp12_v_b_9')
// (3, 19, 'sp4_v_b_11')
// (3, 20, 'sp12_v_b_6')
// (3, 21, 'local_g3_5')
// (3, 21, 'lutff_1/in_3')
// (3, 21, 'sp12_v_b_5')
// (3, 22, 'sp12_v_b_2')
// (3, 23, 'sp12_v_b_1')
// (4, 5, 'sp4_h_l_42')
// (4, 5, 'sp4_v_t_36')
// (4, 6, 'sp4_v_b_36')
// (4, 7, 'sp4_v_b_25')
// (4, 8, 'sp4_v_b_12')
// (4, 8, 'sp4_v_t_42')
// (4, 9, 'sp4_v_b_1')
// (4, 9, 'sp4_v_b_42')
// (4, 9, 'sp4_v_t_47')
// (4, 10, 'sp4_v_b_31')
// (4, 10, 'sp4_v_b_47')
// (4, 11, 'neigh_op_tnl_3')
// (4, 11, 'sp4_v_b_18')
// (4, 11, 'sp4_v_b_34')
// (4, 11, 'sp4_v_t_39')
// (4, 12, 'neigh_op_lft_3')
// (4, 12, 'sp4_h_r_19')
// (4, 12, 'sp4_h_r_35')
// (4, 12, 'sp4_v_b_23')
// (4, 12, 'sp4_v_b_39')
// (4, 12, 'sp4_v_b_7')
// (4, 13, 'neigh_op_bnl_3')
// (4, 13, 'sp4_h_r_10')
// (4, 13, 'sp4_v_b_10')
// (4, 13, 'sp4_v_b_26')
// (4, 14, 'local_g0_7')
// (4, 14, 'lutff_6/in_3')
// (4, 14, 'sp4_v_b_15')
// (4, 15, 'sp4_h_r_8')
// (4, 15, 'sp4_v_b_2')
// (5, 12, 'sp4_h_r_30')
// (5, 12, 'sp4_h_r_46')
// (5, 13, 'local_g1_7')
// (5, 13, 'lutff_2/in_0')
// (5, 13, 'sp4_h_r_23')
// (5, 15, 'sp4_h_r_21')
// (6, 12, 'sp4_h_l_46')
// (6, 12, 'sp4_h_r_43')
// (6, 12, 'sp4_h_r_7')
// (6, 13, 'sp4_h_r_34')
// (6, 15, 'sp4_h_r_32')
// (7, 12, 'sp4_h_l_43')
// (7, 12, 'sp4_h_r_18')
// (7, 12, 'sp4_h_r_6')
// (7, 12, 'sp4_r_v_b_39')
// (7, 13, 'sp4_h_r_47')
// (7, 13, 'sp4_r_v_b_26')
// (7, 14, 'sp4_r_v_b_15')
// (7, 15, 'sp4_h_r_45')
// (7, 15, 'sp4_r_v_b_2')
// (8, 11, 'sp4_v_t_39')
// (8, 12, 'sp4_h_r_19')
// (8, 12, 'sp4_h_r_31')
// (8, 12, 'sp4_v_b_39')
// (8, 13, 'sp4_h_l_47')
// (8, 13, 'sp4_h_r_6')
// (8, 13, 'sp4_v_b_26')
// (8, 14, 'local_g0_7')
// (8, 14, 'lutff_2/in_3')
// (8, 14, 'sp4_v_b_15')
// (8, 15, 'sp4_h_l_45')
// (8, 15, 'sp4_v_b_2')
// (9, 12, 'sp4_h_r_30')
// (9, 12, 'sp4_h_r_42')
// (9, 13, 'sp4_h_r_19')
// (10, 12, 'sp4_h_l_42')
// (10, 12, 'sp4_h_r_3')
// (10, 12, 'sp4_h_r_43')
// (10, 12, 'sp4_h_r_7')
// (10, 13, 'sp4_h_r_30')
// (11, 12, 'local_g1_2')
// (11, 12, 'lutff_1/in_2')
// (11, 12, 'lutff_6/in_1')
// (11, 12, 'sp4_h_l_43')
// (11, 12, 'sp4_h_r_14')
// (11, 12, 'sp4_h_r_18')
// (11, 12, 'sp4_h_r_2')
// (11, 13, 'sp4_h_r_43')
// (12, 12, 'sp4_h_r_15')
// (12, 12, 'sp4_h_r_27')
// (12, 12, 'sp4_h_r_31')
// (12, 13, 'sp4_h_l_43')
// (12, 13, 'sp4_h_r_9')
// (13, 9, 'sp4_r_v_b_36')
// (13, 10, 'sp4_r_v_b_25')
// (13, 11, 'sp4_r_v_b_12')
// (13, 12, 'local_g2_2')
// (13, 12, 'lutff_7/in_3')
// (13, 12, 'sp4_h_r_26')
// (13, 12, 'sp4_h_r_38')
// (13, 12, 'sp4_h_r_42')
// (13, 12, 'sp4_r_v_b_1')
// (13, 13, 'sp4_h_r_20')
// (13, 13, 'sp4_r_v_b_38')
// (13, 14, 'local_g1_3')
// (13, 14, 'lutff_6/in_0')
// (13, 14, 'sp4_r_v_b_27')
// (13, 15, 'sp4_r_v_b_14')
// (13, 16, 'sp4_r_v_b_3')
// (14, 8, 'sp4_v_t_36')
// (14, 9, 'sp4_v_b_36')
// (14, 10, 'local_g2_1')
// (14, 10, 'lutff_1/in_2')
// (14, 10, 'sp4_v_b_25')
// (14, 11, 'sp4_v_b_12')
// (14, 12, 'sp4_h_l_38')
// (14, 12, 'sp4_h_l_42')
// (14, 12, 'sp4_h_r_39')
// (14, 12, 'sp4_v_b_1')
// (14, 12, 'sp4_v_t_38')
// (14, 13, 'local_g3_1')
// (14, 13, 'lutff_0/in_2')
// (14, 13, 'sp4_h_r_33')
// (14, 13, 'sp4_v_b_38')
// (14, 14, 'sp4_v_b_27')
// (14, 15, 'sp4_v_b_14')
// (14, 16, 'sp4_v_b_3')
// (15, 12, 'sp4_h_l_39')
// (15, 13, 'sp4_h_r_44')
// (16, 13, 'sp4_h_l_44')

wire n46;
// (0, 6, 'neigh_op_tnr_1')
// (0, 7, 'neigh_op_rgt_1')
// (0, 8, 'neigh_op_bnr_1')
// (1, 6, 'neigh_op_top_1')
// (1, 7, 'lutff_1/out')
// (1, 8, 'local_g0_1')
// (1, 8, 'lutff_1/in_2')
// (1, 8, 'neigh_op_bot_1')
// (2, 6, 'neigh_op_tnl_1')
// (2, 7, 'neigh_op_lft_1')
// (2, 8, 'neigh_op_bnl_1')

wire n47;
// (0, 6, 'neigh_op_tnr_2')
// (0, 7, 'neigh_op_rgt_2')
// (0, 8, 'neigh_op_bnr_2')
// (1, 6, 'neigh_op_top_2')
// (1, 7, 'lutff_2/out')
// (1, 8, 'local_g0_2')
// (1, 8, 'lutff_2/in_2')
// (1, 8, 'neigh_op_bot_2')
// (2, 6, 'neigh_op_tnl_2')
// (2, 7, 'neigh_op_lft_2')
// (2, 8, 'neigh_op_bnl_2')

wire n48;
// (0, 6, 'neigh_op_tnr_4')
// (0, 7, 'neigh_op_rgt_4')
// (0, 8, 'neigh_op_bnr_4')
// (1, 6, 'local_g0_4')
// (1, 6, 'lutff_2/in_2')
// (1, 6, 'neigh_op_top_4')
// (1, 7, 'local_g0_4')
// (1, 7, 'lutff_2/in_2')
// (1, 7, 'lutff_4/out')
// (1, 8, 'neigh_op_bot_4')
// (2, 6, 'neigh_op_tnl_4')
// (2, 7, 'neigh_op_lft_4')
// (2, 8, 'neigh_op_bnl_4')

wire n49;
// (0, 6, 'neigh_op_tnr_5')
// (0, 7, 'neigh_op_rgt_5')
// (0, 8, 'neigh_op_bnr_5')
// (1, 6, 'local_g1_5')
// (1, 6, 'lutff_1/in_1')
// (1, 6, 'neigh_op_top_5')
// (1, 7, 'local_g1_5')
// (1, 7, 'lutff_1/in_1')
// (1, 7, 'lutff_5/out')
// (1, 8, 'neigh_op_bot_5')
// (2, 6, 'neigh_op_tnl_5')
// (2, 7, 'neigh_op_lft_5')
// (2, 8, 'neigh_op_bnl_5')

wire n50;
// (0, 6, 'neigh_op_tnr_6')
// (0, 7, 'neigh_op_rgt_6')
// (0, 8, 'neigh_op_bnr_6')
// (1, 6, 'local_g1_6')
// (1, 6, 'lutff_3/in_2')
// (1, 6, 'neigh_op_top_6')
// (1, 7, 'lutff_6/out')
// (1, 8, 'neigh_op_bot_6')
// (2, 6, 'neigh_op_tnl_6')
// (2, 7, 'neigh_op_lft_6')
// (2, 8, 'neigh_op_bnl_6')

reg n51 = 0;
// (0, 6, 'sp4_h_r_0')
// (0, 6, 'sp4_h_r_16')
// (1, 5, 'neigh_op_tnr_4')
// (1, 6, 'neigh_op_rgt_4')
// (1, 6, 'sp4_h_r_13')
// (1, 6, 'sp4_h_r_29')
// (1, 7, 'neigh_op_bnr_4')
// (2, 3, 'sp4_r_v_b_44')
// (2, 4, 'sp4_r_v_b_33')
// (2, 5, 'neigh_op_top_4')
// (2, 5, 'sp4_r_v_b_20')
// (2, 6, 'local_g1_4')
// (2, 6, 'lutff_4/in_1')
// (2, 6, 'lutff_4/out')
// (2, 6, 'sp4_h_r_24')
// (2, 6, 'sp4_h_r_40')
// (2, 6, 'sp4_h_r_8')
// (2, 6, 'sp4_r_v_b_9')
// (2, 7, 'local_g0_4')
// (2, 7, 'lutff_3/in_3')
// (2, 7, 'neigh_op_bot_4')
// (3, 1, 'sp4_r_v_b_14')
// (3, 2, 'local_g1_1')
// (3, 2, 'lutff_0/in_2')
// (3, 2, 'sp4_h_r_9')
// (3, 2, 'sp4_r_v_b_3')
// (3, 2, 'sp4_v_t_44')
// (3, 3, 'sp4_r_v_b_37')
// (3, 3, 'sp4_v_b_44')
// (3, 4, 'local_g2_1')
// (3, 4, 'lutff_1/in_0')
// (3, 4, 'sp4_r_v_b_24')
// (3, 4, 'sp4_v_b_33')
// (3, 5, 'local_g3_4')
// (3, 5, 'lutff_5/in_0')
// (3, 5, 'neigh_op_tnl_4')
// (3, 5, 'sp4_r_v_b_13')
// (3, 5, 'sp4_v_b_20')
// (3, 6, 'local_g0_4')
// (3, 6, 'lutff_6/in_2')
// (3, 6, 'neigh_op_lft_4')
// (3, 6, 'sp4_h_l_40')
// (3, 6, 'sp4_h_r_1')
// (3, 6, 'sp4_h_r_21')
// (3, 6, 'sp4_h_r_37')
// (3, 6, 'sp4_r_v_b_0')
// (3, 6, 'sp4_v_b_9')
// (3, 7, 'neigh_op_bnl_4')
// (3, 7, 'sp4_r_v_b_40')
// (3, 8, 'sp4_r_v_b_29')
// (3, 9, 'sp4_r_v_b_16')
// (3, 10, 'sp4_r_v_b_5')
// (4, 0, 'span4_vert_14')
// (4, 1, 'local_g1_6')
// (4, 1, 'lutff_5/in_0')
// (4, 1, 'sp4_v_b_14')
// (4, 2, 'sp4_h_r_20')
// (4, 2, 'sp4_v_b_3')
// (4, 2, 'sp4_v_t_37')
// (4, 3, 'sp4_v_b_37')
// (4, 4, 'sp4_v_b_24')
// (4, 5, 'sp4_v_b_13')
// (4, 6, 'local_g2_0')
// (4, 6, 'local_g3_0')
// (4, 6, 'lutff_5/in_2')
// (4, 6, 'lutff_6/in_0')
// (4, 6, 'sp4_h_l_37')
// (4, 6, 'sp4_h_r_12')
// (4, 6, 'sp4_h_r_32')
// (4, 6, 'sp4_h_r_8')
// (4, 6, 'sp4_v_b_0')
// (4, 6, 'sp4_v_t_40')
// (4, 7, 'sp4_v_b_40')
// (4, 8, 'local_g2_5')
// (4, 8, 'lutff_6/in_1')
// (4, 8, 'sp4_v_b_29')
// (4, 9, 'sp4_v_b_16')
// (4, 10, 'sp4_v_b_5')
// (5, 2, 'local_g2_1')
// (5, 2, 'lutff_5/in_0')
// (5, 2, 'sp4_h_r_33')
// (5, 6, 'sp4_h_r_21')
// (5, 6, 'sp4_h_r_25')
// (5, 6, 'sp4_h_r_45')
// (6, 1, 'sp4_r_v_b_14')
// (6, 2, 'sp4_h_r_44')
// (6, 2, 'sp4_r_v_b_3')
// (6, 3, 'sp4_r_v_b_36')
// (6, 4, 'sp4_r_v_b_25')
// (6, 5, 'sp4_r_v_b_12')
// (6, 6, 'sp4_h_l_45')
// (6, 6, 'sp4_h_r_32')
// (6, 6, 'sp4_h_r_36')
// (6, 6, 'sp4_r_v_b_1')
// (7, 0, 'span4_vert_14')
// (7, 1, 'local_g1_6')
// (7, 1, 'lutff_7/in_2')
// (7, 1, 'sp4_v_b_14')
// (7, 2, 'sp4_h_l_44')
// (7, 2, 'sp4_v_b_3')
// (7, 2, 'sp4_v_t_36')
// (7, 3, 'local_g2_4')
// (7, 3, 'lutff_4/in_2')
// (7, 3, 'sp4_r_v_b_39')
// (7, 3, 'sp4_v_b_36')
// (7, 4, 'sp4_r_v_b_26')
// (7, 4, 'sp4_v_b_25')
// (7, 5, 'sp4_r_v_b_15')
// (7, 5, 'sp4_v_b_12')
// (7, 6, 'sp4_h_l_36')
// (7, 6, 'sp4_h_r_45')
// (7, 6, 'sp4_r_v_b_2')
// (7, 6, 'sp4_v_b_1')
// (8, 2, 'sp4_v_t_39')
// (8, 3, 'sp4_v_b_39')
// (8, 4, 'local_g2_2')
// (8, 4, 'lutff_7/in_3')
// (8, 4, 'sp4_v_b_26')
// (8, 5, 'sp4_v_b_15')
// (8, 6, 'sp4_h_l_45')
// (8, 6, 'sp4_v_b_2')

reg n52 = 0;
// (0, 6, 'sp4_h_r_2')
// (1, 5, 'neigh_op_tnr_5')
// (1, 6, 'neigh_op_rgt_5')
// (1, 6, 'sp4_h_r_15')
// (1, 6, 'sp4_r_v_b_42')
// (1, 7, 'neigh_op_bnr_5')
// (1, 7, 'sp4_r_v_b_31')
// (1, 8, 'sp4_r_v_b_18')
// (1, 9, 'sp4_r_v_b_7')
// (2, 3, 'sp4_r_v_b_46')
// (2, 4, 'sp4_r_v_b_35')
// (2, 5, 'local_g0_5')
// (2, 5, 'lutff_2/in_1')
// (2, 5, 'neigh_op_top_5')
// (2, 5, 'sp4_h_r_0')
// (2, 5, 'sp4_r_v_b_22')
// (2, 5, 'sp4_r_v_b_38')
// (2, 5, 'sp4_v_t_42')
// (2, 6, 'local_g0_5')
// (2, 6, 'lutff_5/in_2')
// (2, 6, 'lutff_5/out')
// (2, 6, 'sp4_h_r_10')
// (2, 6, 'sp4_h_r_26')
// (2, 6, 'sp4_r_v_b_11')
// (2, 6, 'sp4_r_v_b_27')
// (2, 6, 'sp4_v_b_42')
// (2, 7, 'local_g0_5')
// (2, 7, 'lutff_3/in_2')
// (2, 7, 'neigh_op_bot_5')
// (2, 7, 'sp4_r_v_b_14')
// (2, 7, 'sp4_v_b_31')
// (2, 8, 'sp4_r_v_b_3')
// (2, 8, 'sp4_v_b_18')
// (2, 9, 'sp4_v_b_7')
// (3, 2, 'local_g1_4')
// (3, 2, 'lutff_7/in_2')
// (3, 2, 'sp4_h_r_4')
// (3, 2, 'sp4_v_t_46')
// (3, 3, 'sp4_v_b_46')
// (3, 4, 'local_g3_3')
// (3, 4, 'lutff_1/in_3')
// (3, 4, 'sp4_h_r_3')
// (3, 4, 'sp4_v_b_35')
// (3, 4, 'sp4_v_t_38')
// (3, 5, 'local_g3_5')
// (3, 5, 'lutff_3/in_1')
// (3, 5, 'neigh_op_tnl_5')
// (3, 5, 'sp4_h_r_13')
// (3, 5, 'sp4_v_b_22')
// (3, 5, 'sp4_v_b_38')
// (3, 6, 'local_g1_5')
// (3, 6, 'lutff_6/in_0')
// (3, 6, 'neigh_op_lft_5')
// (3, 6, 'sp4_h_r_23')
// (3, 6, 'sp4_h_r_39')
// (3, 6, 'sp4_v_b_11')
// (3, 6, 'sp4_v_b_27')
// (3, 7, 'neigh_op_bnl_5')
// (3, 7, 'sp4_r_v_b_42')
// (3, 7, 'sp4_v_b_14')
// (3, 8, 'sp4_h_r_9')
// (3, 8, 'sp4_r_v_b_31')
// (3, 8, 'sp4_v_b_3')
// (3, 9, 'sp4_r_v_b_18')
// (3, 10, 'sp4_r_v_b_7')
// (4, 2, 'local_g0_1')
// (4, 2, 'lutff_7/in_0')
// (4, 2, 'sp4_h_r_17')
// (4, 4, 'sp4_h_r_14')
// (4, 5, 'local_g2_0')
// (4, 5, 'lutff_4/in_2')
// (4, 5, 'sp4_h_r_24')
// (4, 6, 'sp4_h_l_39')
// (4, 6, 'sp4_h_r_34')
// (4, 6, 'sp4_v_t_42')
// (4, 7, 'local_g3_2')
// (4, 7, 'lutff_1/in_0')
// (4, 7, 'sp4_v_b_42')
// (4, 8, 'local_g1_4')
// (4, 8, 'lutff_7/in_0')
// (4, 8, 'sp4_h_r_20')
// (4, 8, 'sp4_v_b_31')
// (4, 9, 'sp4_v_b_18')
// (4, 10, 'sp4_v_b_7')
// (5, 2, 'local_g3_4')
// (5, 2, 'lutff_5/in_2')
// (5, 2, 'lutff_7/in_2')
// (5, 2, 'sp4_h_r_28')
// (5, 4, 'sp4_h_r_27')
// (5, 5, 'sp4_h_r_37')
// (5, 6, 'local_g3_7')
// (5, 6, 'lutff_2/in_2')
// (5, 6, 'sp4_h_r_47')
// (5, 8, 'sp4_h_r_33')
// (6, 1, 'sp4_r_v_b_17')
// (6, 2, 'sp4_h_r_41')
// (6, 2, 'sp4_r_v_b_4')
// (6, 4, 'sp4_h_r_38')
// (6, 5, 'sp4_h_l_37')
// (6, 6, 'sp4_h_l_47')
// (6, 8, 'sp4_h_r_44')
// (7, 0, 'span4_vert_17')
// (7, 1, 'local_g0_1')
// (7, 1, 'lutff_7/in_0')
// (7, 1, 'sp4_v_b_17')
// (7, 2, 'local_g0_4')
// (7, 2, 'local_g1_4')
// (7, 2, 'lutff_1/in_3')
// (7, 2, 'lutff_5/in_2')
// (7, 2, 'lutff_6/in_3')
// (7, 2, 'sp4_h_l_41')
// (7, 2, 'sp4_h_r_4')
// (7, 2, 'sp4_v_b_4')
// (7, 4, 'sp4_h_l_38')
// (7, 4, 'sp4_h_r_6')
// (7, 8, 'sp4_h_l_44')
// (8, 2, 'sp4_h_r_17')
// (8, 4, 'local_g0_3')
// (8, 4, 'lutff_7/in_0')
// (8, 4, 'sp4_h_r_19')
// (9, 2, 'sp4_h_r_28')
// (9, 4, 'sp4_h_r_30')
// (10, 2, 'sp4_h_r_41')
// (10, 4, 'sp4_h_r_43')
// (11, 2, 'sp4_h_l_41')
// (11, 4, 'sp4_h_l_43')

reg n53 = 0;
// (0, 6, 'sp4_r_v_b_37')
// (0, 7, 'sp4_r_v_b_24')
// (0, 8, 'neigh_op_tnr_0')
// (0, 8, 'sp4_r_v_b_13')
// (0, 9, 'neigh_op_rgt_0')
// (0, 9, 'sp4_h_r_5')
// (0, 9, 'sp4_r_v_b_0')
// (0, 10, 'neigh_op_bnr_0')
// (1, 5, 'sp4_v_t_37')
// (1, 6, 'sp4_v_b_37')
// (1, 7, 'local_g2_0')
// (1, 7, 'lutff_5/in_3')
// (1, 7, 'sp4_v_b_24')
// (1, 8, 'neigh_op_top_0')
// (1, 8, 'sp4_v_b_13')
// (1, 9, 'local_g2_0')
// (1, 9, 'lutff_0/in_2')
// (1, 9, 'lutff_0/out')
// (1, 9, 'sp4_h_r_16')
// (1, 9, 'sp4_v_b_0')
// (1, 10, 'neigh_op_bot_0')
// (2, 8, 'local_g3_0')
// (2, 8, 'lutff_1/in_2')
// (2, 8, 'neigh_op_tnl_0')
// (2, 9, 'local_g1_0')
// (2, 9, 'lutff_5/in_2')
// (2, 9, 'neigh_op_lft_0')
// (2, 9, 'sp4_h_r_29')
// (2, 10, 'neigh_op_bnl_0')
// (3, 6, 'sp4_r_v_b_46')
// (3, 7, 'sp4_r_v_b_35')
// (3, 8, 'local_g3_6')
// (3, 8, 'lutff_1/in_2')
// (3, 8, 'sp4_r_v_b_22')
// (3, 9, 'local_g3_0')
// (3, 9, 'lutff_6/in_1')
// (3, 9, 'sp4_h_r_40')
// (3, 9, 'sp4_r_v_b_11')
// (4, 5, 'sp4_v_t_46')
// (4, 6, 'sp4_v_b_46')
// (4, 7, 'sp4_v_b_35')
// (4, 8, 'sp4_v_b_22')
// (4, 9, 'sp4_h_l_40')
// (4, 9, 'sp4_v_b_11')

wire n54;
// (0, 7, 'neigh_op_tnr_3')
// (0, 8, 'neigh_op_rgt_3')
// (0, 9, 'neigh_op_bnr_3')
// (1, 7, 'neigh_op_top_3')
// (1, 8, 'local_g1_3')
// (1, 8, 'lutff_3/out')
// (1, 8, 'lutff_7/in_3')
// (1, 9, 'neigh_op_bot_3')
// (2, 7, 'neigh_op_tnl_3')
// (2, 8, 'neigh_op_lft_3')
// (2, 9, 'neigh_op_bnl_3')

wire n55;
// (0, 7, 'neigh_op_tnr_4')
// (0, 8, 'neigh_op_rgt_4')
// (0, 9, 'neigh_op_bnr_4')
// (1, 7, 'neigh_op_top_4')
// (1, 8, 'lutff_4/out')
// (1, 9, 'local_g0_4')
// (1, 9, 'lutff_2/in_0')
// (1, 9, 'neigh_op_bot_4')
// (2, 7, 'neigh_op_tnl_4')
// (2, 8, 'neigh_op_lft_4')
// (2, 9, 'neigh_op_bnl_4')

reg n56 = 0;
// (0, 7, 'neigh_op_tnr_5')
// (0, 8, 'neigh_op_rgt_5')
// (0, 9, 'neigh_op_bnr_5')
// (1, 7, 'neigh_op_top_5')
// (1, 8, 'local_g3_5')
// (1, 8, 'lutff_4/in_0')
// (1, 8, 'lutff_5/in_3')
// (1, 8, 'lutff_5/out')
// (1, 9, 'neigh_op_bot_5')
// (2, 7, 'neigh_op_tnl_5')
// (2, 8, 'neigh_op_lft_5')
// (2, 9, 'neigh_op_bnl_5')

wire n57;
// (0, 7, 'neigh_op_tnr_6')
// (0, 8, 'neigh_op_rgt_6')
// (0, 9, 'neigh_op_bnr_6')
// (1, 7, 'neigh_op_top_6')
// (1, 8, 'local_g2_6')
// (1, 8, 'lutff_0/in_2')
// (1, 8, 'lutff_6/out')
// (1, 9, 'neigh_op_bot_6')
// (2, 7, 'neigh_op_tnl_6')
// (2, 8, 'neigh_op_lft_6')
// (2, 9, 'neigh_op_bnl_6')

wire n58;
// (0, 7, 'neigh_op_tnr_7')
// (0, 8, 'neigh_op_rgt_7')
// (0, 9, 'neigh_op_bnr_7')
// (1, 7, 'neigh_op_top_7')
// (1, 8, 'local_g1_7')
// (1, 8, 'lutff_5/in_1')
// (1, 8, 'lutff_7/out')
// (1, 9, 'neigh_op_bot_7')
// (2, 7, 'neigh_op_tnl_7')
// (2, 8, 'neigh_op_lft_7')
// (2, 9, 'neigh_op_bnl_7')

wire n59;
// (0, 7, 'sp12_h_r_2')
// (1, 7, 'sp12_h_r_5')
// (2, 7, 'local_g1_6')
// (2, 7, 'lutff_6/in_1')
// (2, 7, 'sp12_h_r_6')
// (3, 6, 'neigh_op_tnr_1')
// (3, 7, 'neigh_op_rgt_1')
// (3, 7, 'sp12_h_r_9')
// (3, 8, 'neigh_op_bnr_1')
// (4, 6, 'neigh_op_top_1')
// (4, 7, 'lutff_1/out')
// (4, 7, 'sp12_h_r_10')
// (4, 8, 'neigh_op_bot_1')
// (5, 6, 'neigh_op_tnl_1')
// (5, 7, 'neigh_op_lft_1')
// (5, 7, 'sp12_h_r_13')
// (5, 8, 'neigh_op_bnl_1')
// (6, 7, 'sp12_h_r_14')
// (7, 7, 'sp12_h_r_17')
// (8, 7, 'sp12_h_r_18')
// (9, 7, 'sp12_h_r_21')
// (10, 7, 'sp12_h_r_22')
// (11, 7, 'sp12_h_l_22')

reg n60 = 0;
// (0, 7, 'sp4_h_r_12')
// (0, 8, 'sp4_h_r_23')
// (1, 7, 'local_g3_1')
// (1, 7, 'lutff_0/in_2')
// (1, 7, 'sp4_h_r_25')
// (1, 8, 'local_g2_2')
// (1, 8, 'lutff_6/in_0')
// (1, 8, 'sp4_h_r_34')
// (2, 7, 'sp4_h_r_36')
// (2, 8, 'sp4_h_r_47')
// (2, 8, 'sp4_r_v_b_42')
// (2, 9, 'local_g3_1')
// (2, 9, 'lutff_5/in_3')
// (2, 9, 'neigh_op_tnr_1')
// (2, 9, 'sp4_r_v_b_31')
// (2, 9, 'sp4_r_v_b_47')
// (2, 10, 'neigh_op_rgt_1')
// (2, 10, 'sp4_r_v_b_18')
// (2, 10, 'sp4_r_v_b_34')
// (2, 11, 'neigh_op_bnr_1')
// (2, 11, 'sp4_r_v_b_23')
// (2, 11, 'sp4_r_v_b_7')
// (2, 12, 'sp4_r_v_b_10')
// (3, 7, 'sp4_h_l_36')
// (3, 7, 'sp4_v_t_42')
// (3, 8, 'sp4_h_l_47')
// (3, 8, 'sp4_h_r_3')
// (3, 8, 'sp4_r_v_b_43')
// (3, 8, 'sp4_v_b_42')
// (3, 8, 'sp4_v_t_47')
// (3, 9, 'neigh_op_top_1')
// (3, 9, 'sp4_r_v_b_30')
// (3, 9, 'sp4_v_b_31')
// (3, 9, 'sp4_v_b_47')
// (3, 10, 'lutff_1/out')
// (3, 10, 'sp4_r_v_b_19')
// (3, 10, 'sp4_v_b_18')
// (3, 10, 'sp4_v_b_34')
// (3, 11, 'neigh_op_bot_1')
// (3, 11, 'sp4_r_v_b_6')
// (3, 11, 'sp4_v_b_23')
// (3, 11, 'sp4_v_b_7')
// (3, 12, 'sp4_v_b_10')
// (4, 7, 'sp4_v_t_43')
// (4, 8, 'sp4_h_r_14')
// (4, 8, 'sp4_v_b_43')
// (4, 9, 'neigh_op_tnl_1')
// (4, 9, 'sp4_v_b_30')
// (4, 10, 'neigh_op_lft_1')
// (4, 10, 'sp4_v_b_19')
// (4, 11, 'neigh_op_bnl_1')
// (4, 11, 'sp4_h_r_6')
// (4, 11, 'sp4_v_b_6')
// (5, 8, 'local_g3_3')
// (5, 8, 'lutff_2/in_0')
// (5, 8, 'sp4_h_r_27')
// (5, 11, 'sp4_h_r_19')
// (6, 8, 'sp4_h_r_38')
// (6, 11, 'sp4_h_r_30')
// (7, 8, 'sp4_h_l_38')
// (7, 11, 'sp4_h_r_43')
// (8, 11, 'sp4_h_l_43')
// (8, 11, 'sp4_h_r_6')
// (9, 11, 'local_g0_3')
// (9, 11, 'lutff_1/in_2')
// (9, 11, 'sp4_h_r_19')
// (10, 11, 'sp4_h_r_30')
// (11, 11, 'sp4_h_r_43')
// (12, 11, 'sp4_h_l_43')

wire n61;
// (0, 7, 'sp4_h_r_14')
// (1, 7, 'sp4_h_r_27')
// (1, 10, 'neigh_op_tnr_4')
// (1, 11, 'neigh_op_rgt_4')
// (1, 12, 'neigh_op_bnr_4')
// (2, 7, 'local_g2_6')
// (2, 7, 'lutff_6/in_2')
// (2, 7, 'sp4_h_r_38')
// (2, 8, 'sp4_r_v_b_44')
// (2, 9, 'sp4_r_v_b_33')
// (2, 10, 'neigh_op_top_4')
// (2, 10, 'sp4_r_v_b_20')
// (2, 11, 'lutff_4/out')
// (2, 11, 'sp4_r_v_b_9')
// (2, 12, 'neigh_op_bot_4')
// (3, 7, 'sp4_h_l_38')
// (3, 7, 'sp4_v_t_44')
// (3, 8, 'sp4_v_b_44')
// (3, 9, 'sp4_v_b_33')
// (3, 10, 'neigh_op_tnl_4')
// (3, 10, 'sp4_v_b_20')
// (3, 11, 'neigh_op_lft_4')
// (3, 11, 'sp4_v_b_9')
// (3, 12, 'neigh_op_bnl_4')

reg n62 = 0;
// (0, 7, 'sp4_h_r_18')
// (1, 7, 'sp4_h_r_31')
// (1, 13, 'local_g1_2')
// (1, 13, 'lutff_4/in_1')
// (1, 13, 'sp4_h_r_10')
// (2, 4, 'sp4_r_v_b_44')
// (2, 5, 'local_g2_1')
// (2, 5, 'lutff_4/in_1')
// (2, 5, 'sp4_r_v_b_33')
// (2, 6, 'sp4_r_v_b_20')
// (2, 7, 'local_g2_2')
// (2, 7, 'lutff_1/in_1')
// (2, 7, 'sp4_h_r_42')
// (2, 7, 'sp4_r_v_b_9')
// (2, 8, 'sp4_r_v_b_36')
// (2, 9, 'sp4_r_v_b_25')
// (2, 10, 'sp4_r_v_b_12')
// (2, 11, 'sp4_r_v_b_1')
// (2, 13, 'sp4_h_r_23')
// (3, 1, 'sp4_r_v_b_37')
// (3, 2, 'sp4_r_v_b_24')
// (3, 3, 'sp4_r_v_b_13')
// (3, 3, 'sp4_v_t_44')
// (3, 4, 'sp4_r_v_b_0')
// (3, 4, 'sp4_v_b_44')
// (3, 5, 'sp4_r_v_b_44')
// (3, 5, 'sp4_v_b_33')
// (3, 6, 'sp4_r_v_b_33')
// (3, 6, 'sp4_v_b_20')
// (3, 7, 'sp4_h_l_42')
// (3, 7, 'sp4_r_v_b_20')
// (3, 7, 'sp4_v_b_9')
// (3, 7, 'sp4_v_t_36')
// (3, 8, 'sp4_r_v_b_9')
// (3, 8, 'sp4_v_b_36')
// (3, 9, 'sp4_r_v_b_36')
// (3, 9, 'sp4_v_b_25')
// (3, 10, 'neigh_op_tnr_6')
// (3, 10, 'sp4_r_v_b_25')
// (3, 10, 'sp4_v_b_12')
// (3, 11, 'neigh_op_rgt_6')
// (3, 11, 'sp4_h_r_1')
// (3, 11, 'sp4_r_v_b_12')
// (3, 11, 'sp4_v_b_1')
// (3, 12, 'neigh_op_bnr_6')
// (3, 12, 'sp4_r_v_b_1')
// (3, 13, 'sp4_h_r_34')
// (4, 0, 'span4_vert_37')
// (4, 1, 'sp4_v_b_37')
// (4, 2, 'local_g2_0')
// (4, 2, 'lutff_6/in_0')
// (4, 2, 'sp4_v_b_24')
// (4, 3, 'sp4_v_b_13')
// (4, 4, 'sp4_v_b_0')
// (4, 4, 'sp4_v_t_44')
// (4, 5, 'sp4_v_b_44')
// (4, 6, 'sp4_v_b_33')
// (4, 7, 'sp4_v_b_20')
// (4, 8, 'sp4_v_b_9')
// (4, 8, 'sp4_v_t_36')
// (4, 9, 'sp4_v_b_36')
// (4, 10, 'neigh_op_top_6')
// (4, 10, 'sp4_r_v_b_40')
// (4, 10, 'sp4_v_b_25')
// (4, 11, 'local_g1_6')
// (4, 11, 'local_g2_6')
// (4, 11, 'lutff_6/in_2')
// (4, 11, 'lutff_6/out')
// (4, 11, 'lutff_7/in_2')
// (4, 11, 'sp4_h_r_12')
// (4, 11, 'sp4_r_v_b_29')
// (4, 11, 'sp4_v_b_12')
// (4, 12, 'neigh_op_bot_6')
// (4, 12, 'sp4_r_v_b_16')
// (4, 12, 'sp4_v_b_1')
// (4, 13, 'sp4_h_r_47')
// (4, 13, 'sp4_r_v_b_5')
// (5, 9, 'sp4_v_t_40')
// (5, 10, 'neigh_op_tnl_6')
// (5, 10, 'sp4_v_b_40')
// (5, 11, 'neigh_op_lft_6')
// (5, 11, 'sp4_h_r_25')
// (5, 11, 'sp4_v_b_29')
// (5, 12, 'local_g2_6')
// (5, 12, 'lutff_1/in_1')
// (5, 12, 'neigh_op_bnl_6')
// (5, 12, 'sp4_v_b_16')
// (5, 13, 'sp4_h_l_47')
// (5, 13, 'sp4_v_b_5')
// (6, 11, 'sp4_h_r_36')
// (7, 11, 'sp4_h_l_36')

reg n63 = 0;
// (0, 7, 'sp4_h_r_20')
// (1, 7, 'local_g2_1')
// (1, 7, 'lutff_1/in_2')
// (1, 7, 'sp4_h_r_33')
// (2, 7, 'sp4_h_r_44')
// (2, 8, 'sp4_r_v_b_38')
// (2, 9, 'local_g3_7')
// (2, 9, 'lutff_5/in_1')
// (2, 9, 'neigh_op_tnr_7')
// (2, 9, 'sp4_r_v_b_27')
// (2, 10, 'neigh_op_rgt_7')
// (2, 10, 'sp4_h_r_3')
// (2, 10, 'sp4_r_v_b_14')
// (2, 11, 'neigh_op_bnr_7')
// (2, 11, 'sp4_r_v_b_3')
// (3, 7, 'sp4_h_l_44')
// (3, 7, 'sp4_v_t_38')
// (3, 8, 'sp4_v_b_38')
// (3, 9, 'neigh_op_top_7')
// (3, 9, 'sp4_v_b_27')
// (3, 10, 'lutff_7/out')
// (3, 10, 'sp4_h_r_14')
// (3, 10, 'sp4_v_b_14')
// (3, 11, 'neigh_op_bot_7')
// (3, 11, 'sp4_v_b_3')
// (4, 9, 'neigh_op_tnl_7')
// (4, 10, 'neigh_op_lft_7')
// (4, 10, 'sp4_h_r_27')
// (4, 11, 'neigh_op_bnl_7')
// (5, 10, 'local_g2_6')
// (5, 10, 'lutff_3/in_3')
// (5, 10, 'sp4_h_r_38')
// (6, 10, 'sp4_h_l_38')

reg n64 = 0;
// (0, 7, 'sp4_r_v_b_42')
// (0, 8, 'sp4_r_v_b_31')
// (0, 9, 'sp4_r_v_b_18')
// (0, 10, 'sp4_r_v_b_7')
// (1, 6, 'sp4_v_t_42')
// (1, 7, 'local_g3_2')
// (1, 7, 'lutff_2/in_1')
// (1, 7, 'sp4_r_v_b_42')
// (1, 7, 'sp4_v_b_42')
// (1, 8, 'sp4_r_v_b_31')
// (1, 8, 'sp4_v_b_31')
// (1, 9, 'sp4_r_v_b_18')
// (1, 9, 'sp4_v_b_18')
// (1, 10, 'sp4_h_r_7')
// (1, 10, 'sp4_r_v_b_7')
// (1, 10, 'sp4_v_b_7')
// (2, 6, 'sp4_v_t_42')
// (2, 7, 'sp4_v_b_42')
// (2, 8, 'sp4_v_b_31')
// (2, 9, 'local_g1_2')
// (2, 9, 'lutff_6/in_1')
// (2, 9, 'sp4_v_b_18')
// (2, 10, 'sp4_h_r_18')
// (2, 10, 'sp4_h_r_2')
// (2, 10, 'sp4_v_b_7')
// (3, 9, 'neigh_op_tnr_5')
// (3, 10, 'neigh_op_rgt_5')
// (3, 10, 'sp4_h_r_15')
// (3, 10, 'sp4_h_r_31')
// (3, 11, 'neigh_op_bnr_5')
// (4, 9, 'neigh_op_top_5')
// (4, 10, 'lutff_5/out')
// (4, 10, 'sp4_h_r_26')
// (4, 10, 'sp4_h_r_42')
// (4, 11, 'neigh_op_bot_5')
// (5, 9, 'neigh_op_tnl_5')
// (5, 10, 'local_g1_5')
// (5, 10, 'lutff_7/in_1')
// (5, 10, 'neigh_op_lft_5')
// (5, 10, 'sp4_h_l_42')
// (5, 10, 'sp4_h_r_39')
// (5, 11, 'neigh_op_bnl_5')
// (6, 10, 'sp4_h_l_39')

wire n65;
// (0, 8, 'neigh_op_tnr_2')
// (0, 9, 'neigh_op_rgt_2')
// (0, 10, 'neigh_op_bnr_2')
// (1, 8, 'local_g1_2')
// (1, 8, 'lutff_5/in_0')
// (1, 8, 'neigh_op_top_2')
// (1, 9, 'local_g3_2')
// (1, 9, 'lutff_2/out')
// (1, 9, 'lutff_6/in_1')
// (1, 10, 'neigh_op_bot_2')
// (2, 8, 'neigh_op_tnl_2')
// (2, 9, 'neigh_op_lft_2')
// (2, 10, 'local_g2_2')
// (2, 10, 'lutff_0/in_2')
// (2, 10, 'neigh_op_bnl_2')

reg n66 = 0;
// (0, 8, 'neigh_op_tnr_3')
// (0, 9, 'neigh_op_rgt_3')
// (0, 9, 'sp4_r_v_b_38')
// (0, 10, 'neigh_op_bnr_3')
// (0, 10, 'sp4_r_v_b_27')
// (0, 11, 'sp4_r_v_b_14')
// (0, 12, 'sp4_r_v_b_3')
// (1, 8, 'neigh_op_top_3')
// (1, 8, 'sp4_h_r_3')
// (1, 8, 'sp4_v_t_38')
// (1, 9, 'local_g0_3')
// (1, 9, 'lutff_0/in_1')
// (1, 9, 'lutff_3/in_2')
// (1, 9, 'lutff_3/out')
// (1, 9, 'sp4_h_r_6')
// (1, 9, 'sp4_v_b_38')
// (1, 10, 'neigh_op_bot_3')
// (1, 10, 'sp4_v_b_27')
// (1, 11, 'sp4_v_b_14')
// (1, 12, 'sp4_v_b_3')
// (2, 8, 'local_g2_3')
// (2, 8, 'lutff_0/in_1')
// (2, 8, 'lutff_5/in_0')
// (2, 8, 'neigh_op_tnl_3')
// (2, 8, 'sp4_h_r_14')
// (2, 9, 'local_g0_3')
// (2, 9, 'lutff_5/in_0')
// (2, 9, 'neigh_op_lft_3')
// (2, 9, 'sp4_h_r_19')
// (2, 10, 'neigh_op_bnl_3')
// (3, 8, 'local_g3_3')
// (3, 8, 'lutff_0/in_2')
// (3, 8, 'lutff_1/in_3')
// (3, 8, 'lutff_4/in_2')
// (3, 8, 'sp4_h_r_27')
// (3, 9, 'local_g3_6')
// (3, 9, 'lutff_5/in_0')
// (3, 9, 'sp4_h_r_30')
// (4, 8, 'sp4_h_r_38')
// (4, 9, 'sp4_h_r_43')
// (5, 8, 'sp4_h_l_38')
// (5, 9, 'sp4_h_l_43')

reg n67 = 0;
// (0, 8, 'neigh_op_tnr_5')
// (0, 9, 'neigh_op_rgt_5')
// (0, 10, 'neigh_op_bnr_5')
// (1, 8, 'neigh_op_top_5')
// (1, 9, 'local_g1_5')
// (1, 9, 'lutff_2/in_2')
// (1, 9, 'lutff_5/out')
// (1, 10, 'neigh_op_bot_5')
// (2, 8, 'neigh_op_tnl_5')
// (2, 9, 'neigh_op_lft_5')
// (2, 10, 'neigh_op_bnl_5')

wire n68;
// (0, 8, 'neigh_op_tnr_6')
// (0, 9, 'neigh_op_rgt_6')
// (0, 10, 'neigh_op_bnr_6')
// (1, 8, 'neigh_op_top_6')
// (1, 9, 'lutff_6/out')
// (1, 10, 'neigh_op_bot_6')
// (2, 8, 'local_g2_6')
// (2, 8, 'lutff_6/in_0')
// (2, 8, 'neigh_op_tnl_6')
// (2, 9, 'local_g1_6')
// (2, 9, 'lutff_4/in_3')
// (2, 9, 'lutff_7/in_2')
// (2, 9, 'neigh_op_lft_6')
// (2, 10, 'neigh_op_bnl_6')

wire n69;
// (0, 8, 'sp4_h_r_13')
// (0, 8, 'sp4_h_r_19')
// (0, 12, 'sp4_h_r_16')
// (1, 8, 'local_g2_0')
// (1, 8, 'local_g3_6')
// (1, 8, 'lutff_4/in_2')
// (1, 8, 'lutff_7/in_2')
// (1, 8, 'sp4_h_r_24')
// (1, 8, 'sp4_h_r_30')
// (1, 10, 'local_g1_0')
// (1, 10, 'lutff_0/in_3')
// (1, 10, 'lutff_1/in_2')
// (1, 10, 'sp4_h_r_0')
// (1, 12, 'local_g3_5')
// (1, 12, 'lutff_1/in_3')
// (1, 12, 'sp4_h_r_29')
// (2, 8, 'sp4_h_r_37')
// (2, 8, 'sp4_h_r_43')
// (2, 9, 'neigh_op_tnr_4')
// (2, 9, 'sp4_r_v_b_37')
// (2, 10, 'neigh_op_rgt_4')
// (2, 10, 'sp4_h_r_13')
// (2, 10, 'sp4_r_v_b_24')
// (2, 11, 'neigh_op_bnr_4')
// (2, 11, 'sp4_r_v_b_13')
// (2, 12, 'sp4_h_r_40')
// (2, 12, 'sp4_r_v_b_0')
// (3, 8, 'sp4_h_l_37')
// (3, 8, 'sp4_h_l_43')
// (3, 8, 'sp4_v_t_37')
// (3, 9, 'local_g0_4')
// (3, 9, 'lutff_7/in_3')
// (3, 9, 'neigh_op_top_4')
// (3, 9, 'sp4_v_b_37')
// (3, 10, 'lutff_4/out')
// (3, 10, 'sp4_h_r_24')
// (3, 10, 'sp4_v_b_24')
// (3, 11, 'neigh_op_bot_4')
// (3, 11, 'sp4_v_b_13')
// (3, 12, 'sp4_h_l_40')
// (3, 12, 'sp4_v_b_0')
// (4, 9, 'neigh_op_tnl_4')
// (4, 10, 'neigh_op_lft_4')
// (4, 10, 'sp4_h_r_37')
// (4, 11, 'neigh_op_bnl_4')
// (5, 10, 'sp4_h_l_37')

reg n70 = 0;
// (0, 8, 'sp4_h_r_18')
// (0, 9, 'sp4_h_r_23')
// (0, 9, 'sp4_r_v_b_40')
// (0, 9, 'sp4_r_v_b_47')
// (0, 10, 'sp4_r_v_b_29')
// (0, 10, 'sp4_r_v_b_34')
// (0, 11, 'sp4_r_v_b_16')
// (0, 11, 'sp4_r_v_b_23')
// (0, 12, 'sp4_r_v_b_10')
// (0, 12, 'sp4_r_v_b_5')
// (1, 8, 'sp4_h_r_31')
// (1, 8, 'sp4_v_t_40')
// (1, 8, 'sp4_v_t_47')
// (1, 9, 'local_g2_2')
// (1, 9, 'local_g3_0')
// (1, 9, 'lutff_2/in_1')
// (1, 9, 'lutff_global/cen')
// (1, 9, 'sp4_h_r_34')
// (1, 9, 'sp4_v_b_40')
// (1, 9, 'sp4_v_b_47')
// (1, 10, 'local_g2_2')
// (1, 10, 'lutff_global/cen')
// (1, 10, 'sp4_v_b_29')
// (1, 10, 'sp4_v_b_34')
// (1, 11, 'local_g2_0')
// (1, 11, 'lutff_0/in_2')
// (1, 11, 'lutff_2/in_2')
// (1, 11, 'neigh_op_tnr_0')
// (1, 11, 'sp4_v_b_16')
// (1, 11, 'sp4_v_b_23')
// (1, 12, 'neigh_op_rgt_0')
// (1, 12, 'sp4_h_r_5')
// (1, 12, 'sp4_v_b_10')
// (1, 12, 'sp4_v_b_5')
// (1, 13, 'neigh_op_bnr_0')
// (2, 8, 'local_g2_2')
// (2, 8, 'lutff_global/cen')
// (2, 8, 'sp4_h_r_42')
// (2, 9, 'sp4_h_r_47')
// (2, 9, 'sp4_r_v_b_36')
// (2, 9, 'sp4_r_v_b_43')
// (2, 10, 'sp4_r_v_b_25')
// (2, 10, 'sp4_r_v_b_30')
// (2, 10, 'sp4_r_v_b_41')
// (2, 11, 'local_g1_0')
// (2, 11, 'lutff_3/in_0')
// (2, 11, 'neigh_op_top_0')
// (2, 11, 'sp4_r_v_b_12')
// (2, 11, 'sp4_r_v_b_19')
// (2, 11, 'sp4_r_v_b_28')
// (2, 12, 'lutff_0/out')
// (2, 12, 'sp4_h_r_16')
// (2, 12, 'sp4_r_v_b_1')
// (2, 12, 'sp4_r_v_b_17')
// (2, 12, 'sp4_r_v_b_6')
// (2, 13, 'neigh_op_bot_0')
// (2, 13, 'sp4_r_v_b_4')
// (3, 8, 'sp4_h_l_42')
// (3, 8, 'sp4_h_r_6')
// (3, 8, 'sp4_v_t_36')
// (3, 8, 'sp4_v_t_43')
// (3, 9, 'local_g3_3')
// (3, 9, 'lutff_global/cen')
// (3, 9, 'sp4_h_l_47')
// (3, 9, 'sp4_v_b_36')
// (3, 9, 'sp4_v_b_43')
// (3, 9, 'sp4_v_t_41')
// (3, 10, 'sp4_v_b_25')
// (3, 10, 'sp4_v_b_30')
// (3, 10, 'sp4_v_b_41')
// (3, 11, 'local_g1_3')
// (3, 11, 'lutff_global/cen')
// (3, 11, 'neigh_op_tnl_0')
// (3, 11, 'sp4_v_b_12')
// (3, 11, 'sp4_v_b_19')
// (3, 11, 'sp4_v_b_28')
// (3, 12, 'neigh_op_lft_0')
// (3, 12, 'sp4_h_r_29')
// (3, 12, 'sp4_v_b_1')
// (3, 12, 'sp4_v_b_17')
// (3, 12, 'sp4_v_b_6')
// (3, 13, 'neigh_op_bnl_0')
// (3, 13, 'sp4_v_b_4')
// (4, 8, 'sp4_h_r_19')
// (4, 12, 'sp4_h_r_40')
// (5, 8, 'sp4_h_r_30')
// (5, 12, 'sp4_h_l_40')
// (6, 8, 'sp4_h_r_43')
// (7, 8, 'sp4_h_l_43')

wire n71;
// (0, 8, 'sp4_h_r_4')
// (1, 7, 'neigh_op_tnr_6')
// (1, 8, 'neigh_op_rgt_6')
// (1, 8, 'sp4_h_r_17')
// (1, 9, 'neigh_op_bnr_6')
// (2, 7, 'neigh_op_top_6')
// (2, 8, 'lutff_6/out')
// (2, 8, 'sp4_h_r_28')
// (2, 9, 'neigh_op_bot_6')
// (3, 5, 'sp4_r_v_b_47')
// (3, 6, 'sp4_r_v_b_34')
// (3, 7, 'neigh_op_tnl_6')
// (3, 7, 'sp4_r_v_b_23')
// (3, 8, 'local_g2_2')
// (3, 8, 'lutff_global/cen')
// (3, 8, 'neigh_op_lft_6')
// (3, 8, 'sp4_h_r_41')
// (3, 8, 'sp4_r_v_b_10')
// (3, 9, 'neigh_op_bnl_6')
// (4, 4, 'sp4_v_t_47')
// (4, 5, 'sp4_v_b_47')
// (4, 6, 'sp4_v_b_34')
// (4, 7, 'sp4_v_b_23')
// (4, 8, 'sp4_h_l_41')
// (4, 8, 'sp4_v_b_10')

wire n72;
// (0, 9, 'neigh_op_tnr_0')
// (0, 10, 'neigh_op_rgt_0')
// (0, 11, 'neigh_op_bnr_0')
// (1, 9, 'local_g1_0')
// (1, 9, 'lutff_5/in_2')
// (1, 9, 'lutff_6/in_3')
// (1, 9, 'neigh_op_top_0')
// (1, 10, 'lutff_0/out')
// (1, 11, 'neigh_op_bot_0')
// (2, 9, 'neigh_op_tnl_0')
// (2, 10, 'neigh_op_lft_0')
// (2, 11, 'neigh_op_bnl_0')

wire n73;
// (0, 9, 'neigh_op_tnr_1')
// (0, 10, 'neigh_op_rgt_1')
// (0, 11, 'neigh_op_bnr_1')
// (1, 9, 'neigh_op_top_1')
// (1, 10, 'lutff_1/out')
// (1, 11, 'neigh_op_bot_1')
// (2, 9, 'neigh_op_tnl_1')
// (2, 10, 'neigh_op_lft_1')
// (2, 11, 'local_g3_1')
// (2, 11, 'lutff_3/in_1')
// (2, 11, 'neigh_op_bnl_1')

reg n74 = 0;
// (0, 9, 'neigh_op_tnr_7')
// (0, 9, 'sp4_r_v_b_43')
// (0, 10, 'neigh_op_rgt_7')
// (0, 10, 'sp4_r_v_b_30')
// (0, 11, 'neigh_op_bnr_7')
// (0, 11, 'sp4_r_v_b_19')
// (0, 12, 'sp4_r_v_b_6')
// (1, 8, 'sp4_r_v_b_39')
// (1, 8, 'sp4_v_t_43')
// (1, 9, 'neigh_op_top_7')
// (1, 9, 'sp4_r_v_b_26')
// (1, 9, 'sp4_v_b_43')
// (1, 10, 'lutff_7/out')
// (1, 10, 'sp4_r_v_b_15')
// (1, 10, 'sp4_v_b_30')
// (1, 11, 'neigh_op_bot_7')
// (1, 11, 'sp4_r_v_b_2')
// (1, 11, 'sp4_v_b_19')
// (1, 12, 'sp4_h_r_0')
// (1, 12, 'sp4_v_b_6')
// (2, 7, 'sp4_v_t_39')
// (2, 8, 'sp4_v_b_39')
// (2, 9, 'neigh_op_tnl_7')
// (2, 9, 'sp4_v_b_26')
// (2, 10, 'neigh_op_lft_7')
// (2, 10, 'sp4_v_b_15')
// (2, 11, 'neigh_op_bnl_7')
// (2, 11, 'sp4_h_r_2')
// (2, 11, 'sp4_v_b_2')
// (2, 12, 'sp4_h_r_13')
// (3, 11, 'local_g0_7')
// (3, 11, 'lutff_2/in_3')
// (3, 11, 'sp4_h_r_15')
// (3, 12, 'local_g3_0')
// (3, 12, 'lutff_3/in_2')
// (3, 12, 'sp4_h_r_24')
// (4, 11, 'sp4_h_r_26')
// (4, 12, 'sp4_h_r_37')
// (5, 11, 'sp4_h_r_39')
// (5, 12, 'sp4_h_l_37')
// (6, 11, 'sp4_h_l_39')

wire n75;
// (0, 9, 'sp4_r_v_b_36')
// (0, 10, 'neigh_op_tnr_6')
// (0, 10, 'sp4_r_v_b_25')
// (0, 11, 'neigh_op_rgt_6')
// (0, 11, 'sp4_r_v_b_12')
// (0, 12, 'neigh_op_bnr_6')
// (0, 12, 'sp4_r_v_b_1')
// (1, 8, 'sp4_v_t_36')
// (1, 9, 'local_g3_4')
// (1, 9, 'lutff_2/in_3')
// (1, 9, 'sp4_v_b_36')
// (1, 10, 'local_g0_6')
// (1, 10, 'lutff_1/in_1')
// (1, 10, 'neigh_op_top_6')
// (1, 10, 'sp4_v_b_25')
// (1, 11, 'local_g0_6')
// (1, 11, 'lutff_0/in_0')
// (1, 11, 'lutff_2/in_0')
// (1, 11, 'lutff_3/in_3')
// (1, 11, 'lutff_6/out')
// (1, 11, 'sp4_v_b_12')
// (1, 12, 'neigh_op_bot_6')
// (1, 12, 'sp4_v_b_1')
// (2, 10, 'neigh_op_tnl_6')
// (2, 11, 'neigh_op_lft_6')
// (2, 12, 'neigh_op_bnl_6')

wire n76;
// (0, 10, 'neigh_op_tnr_0')
// (0, 11, 'neigh_op_rgt_0')
// (0, 11, 'sp4_h_r_21')
// (0, 12, 'neigh_op_bnr_0')
// (0, 12, 'sp4_r_v_b_37')
// (0, 13, 'sp4_r_v_b_24')
// (0, 14, 'sp4_r_v_b_13')
// (0, 15, 'sp4_r_v_b_0')
// (1, 10, 'local_g0_0')
// (1, 10, 'lutff_0/in_2')
// (1, 10, 'neigh_op_top_0')
// (1, 11, 'lutff_0/out')
// (1, 11, 'sp4_h_r_0')
// (1, 11, 'sp4_h_r_32')
// (1, 11, 'sp4_v_t_37')
// (1, 12, 'neigh_op_bot_0')
// (1, 12, 'sp4_v_b_37')
// (1, 13, 'sp4_v_b_24')
// (1, 14, 'local_g0_5')
// (1, 14, 'lutff_1/in_0')
// (1, 14, 'sp4_v_b_13')
// (1, 15, 'sp4_v_b_0')
// (2, 10, 'neigh_op_tnl_0')
// (2, 11, 'neigh_op_lft_0')
// (2, 11, 'sp4_h_r_13')
// (2, 11, 'sp4_h_r_45')
// (2, 12, 'neigh_op_bnl_0')
// (2, 12, 'sp4_r_v_b_45')
// (2, 13, 'sp4_r_v_b_32')
// (2, 14, 'sp4_r_v_b_21')
// (2, 15, 'sp4_r_v_b_8')
// (3, 11, 'sp4_h_l_45')
// (3, 11, 'sp4_h_r_24')
// (3, 11, 'sp4_v_t_45')
// (3, 12, 'sp4_v_b_45')
// (3, 13, 'sp4_v_b_32')
// (3, 14, 'local_g1_5')
// (3, 14, 'lutff_5/in_3')
// (3, 14, 'sp4_v_b_21')
// (3, 15, 'sp4_v_b_8')
// (4, 11, 'sp4_h_r_37')
// (5, 11, 'sp4_h_l_37')

wire n77;
// (0, 10, 'neigh_op_tnr_2')
// (0, 11, 'neigh_op_rgt_2')
// (0, 12, 'neigh_op_bnr_2')
// (1, 10, 'neigh_op_top_2')
// (1, 11, 'lutff_2/out')
// (1, 12, 'neigh_op_bot_2')
// (2, 10, 'local_g3_2')
// (2, 10, 'lutff_4/in_1')
// (2, 10, 'neigh_op_tnl_2')
// (2, 11, 'neigh_op_lft_2')
// (2, 12, 'neigh_op_bnl_2')

reg n78 = 0;
// (0, 10, 'neigh_op_tnr_7')
// (0, 11, 'neigh_op_rgt_7')
// (0, 11, 'sp4_r_v_b_46')
// (0, 12, 'neigh_op_bnr_7')
// (0, 12, 'sp4_r_v_b_35')
// (0, 13, 'sp4_r_v_b_22')
// (0, 14, 'sp4_r_v_b_11')
// (1, 10, 'neigh_op_top_7')
// (1, 10, 'sp4_v_t_46')
// (1, 11, 'lutff_7/out')
// (1, 11, 'sp4_v_b_46')
// (1, 12, 'neigh_op_bot_7')
// (1, 12, 'sp4_v_b_35')
// (1, 13, 'sp4_v_b_22')
// (1, 14, 'local_g0_3')
// (1, 14, 'lutff_7/in_0')
// (1, 14, 'sp4_v_b_11')
// (2, 10, 'neigh_op_tnl_7')
// (2, 11, 'neigh_op_lft_7')
// (2, 12, 'neigh_op_bnl_7')

reg n79 = 0;
// (0, 10, 'sp12_h_r_17')
// (0, 11, 'sp4_h_r_5')
// (1, 10, 'local_g1_2')
// (1, 10, 'lutff_7/in_0')
// (1, 10, 'sp12_h_r_18')
// (1, 11, 'local_g1_0')
// (1, 11, 'lutff_6/in_1')
// (1, 11, 'sp4_h_r_16')
// (2, 10, 'sp12_h_r_21')
// (2, 11, 'sp4_h_r_29')
// (3, 2, 'sp4_r_v_b_38')
// (3, 3, 'sp4_r_v_b_27')
// (3, 4, 'sp4_r_v_b_14')
// (3, 5, 'sp4_r_v_b_3')
// (3, 6, 'sp4_r_v_b_38')
// (3, 7, 'sp4_r_v_b_27')
// (3, 8, 'sp4_r_v_b_14')
// (3, 8, 'sp4_r_v_b_40')
// (3, 9, 'sp4_r_v_b_29')
// (3, 9, 'sp4_r_v_b_3')
// (3, 10, 'local_g3_0')
// (3, 10, 'lutff_4/in_1')
// (3, 10, 'sp12_h_r_22')
// (3, 10, 'sp4_r_v_b_16')
// (3, 10, 'sp4_r_v_b_43')
// (3, 11, 'sp4_h_r_40')
// (3, 11, 'sp4_r_v_b_30')
// (3, 11, 'sp4_r_v_b_5')
// (3, 12, 'local_g3_3')
// (3, 12, 'lutff_3/in_1')
// (3, 12, 'sp4_r_v_b_19')
// (3, 13, 'sp4_r_v_b_6')
// (4, 1, 'sp4_h_r_3')
// (4, 1, 'sp4_v_t_38')
// (4, 2, 'sp4_v_b_38')
// (4, 3, 'sp4_v_b_27')
// (4, 4, 'sp4_v_b_14')
// (4, 5, 'sp4_v_b_3')
// (4, 5, 'sp4_v_t_38')
// (4, 6, 'sp4_v_b_38')
// (4, 7, 'sp4_h_r_5')
// (4, 7, 'sp4_v_b_27')
// (4, 7, 'sp4_v_t_40')
// (4, 8, 'sp4_v_b_14')
// (4, 8, 'sp4_v_b_40')
// (4, 9, 'sp4_v_b_29')
// (4, 9, 'sp4_v_b_3')
// (4, 9, 'sp4_v_t_43')
// (4, 10, 'sp12_h_l_22')
// (4, 10, 'sp12_h_r_1')
// (4, 10, 'sp4_v_b_16')
// (4, 10, 'sp4_v_b_43')
// (4, 11, 'sp4_h_l_40')
// (4, 11, 'sp4_v_b_30')
// (4, 11, 'sp4_v_b_5')
// (4, 12, 'sp4_v_b_19')
// (4, 13, 'sp4_v_b_6')
// (5, 1, 'sp4_h_r_14')
// (5, 7, 'sp4_h_r_16')
// (5, 10, 'sp12_h_r_2')
// (6, 1, 'sp4_h_r_27')
// (6, 7, 'sp4_h_r_29')
// (6, 10, 'sp12_h_r_5')
// (7, 1, 'sp4_h_r_38')
// (7, 4, 'sp4_r_v_b_40')
// (7, 5, 'sp4_r_v_b_29')
// (7, 6, 'sp4_r_v_b_16')
// (7, 7, 'sp4_h_r_40')
// (7, 7, 'sp4_r_v_b_5')
// (7, 10, 'sp12_h_r_6')
// (8, 1, 'sp4_h_l_38')
// (8, 1, 'sp4_h_r_3')
// (8, 3, 'sp4_h_r_11')
// (8, 3, 'sp4_v_t_40')
// (8, 4, 'sp4_v_b_40')
// (8, 5, 'sp4_v_b_29')
// (8, 6, 'sp4_v_b_16')
// (8, 7, 'sp4_h_l_40')
// (8, 7, 'sp4_v_b_5')
// (8, 10, 'sp12_h_r_9')
// (9, 1, 'sp4_h_r_14')
// (9, 3, 'sp4_h_r_22')
// (9, 10, 'sp12_h_r_10')
// (10, 1, 'sp4_h_r_27')
// (10, 3, 'sp4_h_r_35')
// (10, 10, 'sp12_h_r_13')
// (11, 1, 'sp4_h_r_38')
// (11, 3, 'sp4_h_r_46')
// (11, 10, 'sp12_h_r_14')
// (12, 1, 'sp4_h_l_38')
// (12, 1, 'sp4_h_r_7')
// (12, 3, 'sp4_h_l_46')
// (12, 3, 'sp4_h_r_3')
// (12, 10, 'sp12_h_r_17')
// (13, 1, 'sp4_h_r_18')
// (13, 3, 'sp4_h_r_14')
// (13, 10, 'sp12_h_r_18')
// (14, 1, 'sp4_h_r_31')
// (14, 3, 'sp4_h_r_27')
// (14, 10, 'sp12_h_r_21')
// (15, 0, 'logic_op_tnr_1')
// (15, 1, 'neigh_op_rgt_1')
// (15, 1, 'sp4_h_r_42')
// (15, 1, 'sp4_r_v_b_2')
// (15, 1, 'sp4_r_v_b_34')
// (15, 2, 'neigh_op_bnr_1')
// (15, 2, 'sp4_r_v_b_23')
// (15, 3, 'sp4_h_r_38')
// (15, 3, 'sp4_r_v_b_10')
// (15, 10, 'sp12_h_r_22')
// (16, 0, 'logic_op_top_1')
// (16, 0, 'span12_vert_18')
// (16, 0, 'span4_vert_2')
// (16, 0, 'span4_vert_34')
// (16, 1, 'lutff_1/out')
// (16, 1, 'sp12_v_b_18')
// (16, 1, 'sp4_h_l_42')
// (16, 1, 'sp4_v_b_2')
// (16, 1, 'sp4_v_b_34')
// (16, 2, 'neigh_op_bot_1')
// (16, 2, 'sp12_v_b_17')
// (16, 2, 'sp4_v_b_23')
// (16, 3, 'sp12_v_b_14')
// (16, 3, 'sp4_h_l_38')
// (16, 3, 'sp4_v_b_10')
// (16, 4, 'sp12_v_b_13')
// (16, 5, 'sp12_v_b_10')
// (16, 6, 'sp12_v_b_9')
// (16, 7, 'sp12_v_b_6')
// (16, 8, 'sp12_v_b_5')
// (16, 9, 'sp12_v_b_2')
// (16, 10, 'sp12_h_l_22')
// (16, 10, 'sp12_v_b_1')
// (17, 0, 'logic_op_tnl_1')
// (17, 1, 'neigh_op_lft_1')
// (17, 2, 'neigh_op_bnl_1')

reg n80 = 0;
// (0, 10, 'sp4_h_r_5')
// (0, 15, 'sp4_r_v_b_39')
// (0, 16, 'sp4_r_v_b_26')
// (0, 17, 'sp4_r_v_b_15')
// (0, 18, 'sp4_r_v_b_2')
// (0, 19, 'sp4_r_v_b_40')
// (0, 20, 'sp4_r_v_b_29')
// (0, 21, 'sp4_h_r_7')
// (0, 21, 'sp4_r_v_b_16')
// (0, 22, 'sp4_r_v_b_5')
// (1, 10, 'sp4_h_r_16')
// (1, 14, 'local_g1_2')
// (1, 14, 'lutff_0/in_1')
// (1, 14, 'lutff_3/in_2')
// (1, 14, 'sp4_h_r_2')
// (1, 14, 'sp4_v_t_39')
// (1, 15, 'sp4_v_b_39')
// (1, 16, 'sp4_v_b_26')
// (1, 17, 'sp4_v_b_15')
// (1, 18, 'sp4_v_b_2')
// (1, 18, 'sp4_v_t_40')
// (1, 19, 'sp4_v_b_40')
// (1, 20, 'local_g2_5')
// (1, 20, 'lutff_3/in_0')
// (1, 20, 'sp4_v_b_29')
// (1, 21, 'local_g0_2')
// (1, 21, 'lutff_global/cen')
// (1, 21, 'sp4_h_r_18')
// (1, 21, 'sp4_v_b_16')
// (1, 22, 'sp4_v_b_5')
// (2, 10, 'local_g3_5')
// (2, 10, 'lutff_3/in_1')
// (2, 10, 'sp4_h_r_29')
// (2, 13, 'local_g2_5')
// (2, 13, 'lutff_1/in_0')
// (2, 13, 'lutff_7/in_0')
// (2, 13, 'neigh_op_tnr_5')
// (2, 13, 'sp4_r_v_b_39')
// (2, 14, 'local_g3_5')
// (2, 14, 'lutff_0/in_0')
// (2, 14, 'neigh_op_rgt_5')
// (2, 14, 'sp4_h_r_15')
// (2, 14, 'sp4_r_v_b_26')
// (2, 15, 'neigh_op_bnr_5')
// (2, 15, 'sp4_r_v_b_15')
// (2, 16, 'local_g1_2')
// (2, 16, 'lutff_0/in_3')
// (2, 16, 'lutff_5/in_0')
// (2, 16, 'sp4_r_v_b_2')
// (2, 17, 'sp4_r_v_b_40')
// (2, 18, 'sp4_r_v_b_29')
// (2, 19, 'sp4_r_v_b_16')
// (2, 20, 'local_g1_5')
// (2, 20, 'lutff_6/in_0')
// (2, 20, 'sp4_r_v_b_5')
// (2, 21, 'sp4_h_r_31')
// (3, 10, 'sp4_h_r_40')
// (3, 11, 'sp4_r_v_b_46')
// (3, 12, 'sp4_r_v_b_35')
// (3, 12, 'sp4_v_t_39')
// (3, 13, 'neigh_op_top_5')
// (3, 13, 'sp4_r_v_b_22')
// (3, 13, 'sp4_v_b_39')
// (3, 14, 'local_g2_5')
// (3, 14, 'lutff_5/in_0')
// (3, 14, 'lutff_5/out')
// (3, 14, 'sp4_h_r_10')
// (3, 14, 'sp4_h_r_26')
// (3, 14, 'sp4_r_v_b_11')
// (3, 14, 'sp4_r_v_b_43')
// (3, 14, 'sp4_v_b_26')
// (3, 15, 'local_g1_5')
// (3, 15, 'lutff_4/in_0')
// (3, 15, 'neigh_op_bot_5')
// (3, 15, 'sp4_r_v_b_30')
// (3, 15, 'sp4_v_b_15')
// (3, 16, 'local_g3_3')
// (3, 16, 'lutff_1/in_3')
// (3, 16, 'lutff_3/in_1')
// (3, 16, 'lutff_5/in_1')
// (3, 16, 'lutff_7/in_3')
// (3, 16, 'sp4_r_v_b_19')
// (3, 16, 'sp4_v_b_2')
// (3, 16, 'sp4_v_t_40')
// (3, 17, 'sp4_r_v_b_6')
// (3, 17, 'sp4_v_b_40')
// (3, 18, 'sp4_r_v_b_39')
// (3, 18, 'sp4_r_v_b_44')
// (3, 18, 'sp4_v_b_29')
// (3, 19, 'sp4_r_v_b_26')
// (3, 19, 'sp4_r_v_b_33')
// (3, 19, 'sp4_v_b_16')
// (3, 20, 'local_g3_4')
// (3, 20, 'lutff_1/in_2')
// (3, 20, 'sp4_r_v_b_15')
// (3, 20, 'sp4_r_v_b_20')
// (3, 20, 'sp4_v_b_5')
// (3, 21, 'sp4_h_r_42')
// (3, 21, 'sp4_r_v_b_2')
// (3, 21, 'sp4_r_v_b_9')
// (4, 10, 'sp4_h_l_40')
// (4, 10, 'sp4_v_t_46')
// (4, 11, 'sp4_v_b_46')
// (4, 12, 'sp4_v_b_35')
// (4, 13, 'neigh_op_tnl_5')
// (4, 13, 'sp4_v_b_22')
// (4, 13, 'sp4_v_t_43')
// (4, 14, 'neigh_op_lft_5')
// (4, 14, 'sp4_h_r_23')
// (4, 14, 'sp4_h_r_39')
// (4, 14, 'sp4_v_b_11')
// (4, 14, 'sp4_v_b_43')
// (4, 15, 'local_g2_5')
// (4, 15, 'lutff_2/in_3')
// (4, 15, 'neigh_op_bnl_5')
// (4, 15, 'sp4_r_v_b_39')
// (4, 15, 'sp4_v_b_30')
// (4, 16, 'sp4_r_v_b_26')
// (4, 16, 'sp4_v_b_19')
// (4, 17, 'local_g1_6')
// (4, 17, 'lutff_6/in_3')
// (4, 17, 'sp4_r_v_b_15')
// (4, 17, 'sp4_v_b_6')
// (4, 17, 'sp4_v_t_39')
// (4, 17, 'sp4_v_t_44')
// (4, 18, 'sp4_r_v_b_2')
// (4, 18, 'sp4_v_b_39')
// (4, 18, 'sp4_v_b_44')
// (4, 19, 'sp4_r_v_b_40')
// (4, 19, 'sp4_v_b_26')
// (4, 19, 'sp4_v_b_33')
// (4, 20, 'sp4_r_v_b_29')
// (4, 20, 'sp4_v_b_15')
// (4, 20, 'sp4_v_b_20')
// (4, 21, 'sp4_h_l_42')
// (4, 21, 'sp4_r_v_b_16')
// (4, 21, 'sp4_v_b_2')
// (4, 21, 'sp4_v_b_9')
// (4, 22, 'sp4_r_v_b_5')
// (5, 14, 'sp4_h_l_39')
// (5, 14, 'sp4_h_r_34')
// (5, 14, 'sp4_v_t_39')
// (5, 15, 'sp4_v_b_39')
// (5, 16, 'local_g2_2')
// (5, 16, 'lutff_global/cen')
// (5, 16, 'sp4_v_b_26')
// (5, 17, 'sp4_v_b_15')
// (5, 18, 'sp4_v_b_2')
// (5, 18, 'sp4_v_t_40')
// (5, 19, 'local_g3_0')
// (5, 19, 'lutff_1/in_2')
// (5, 19, 'sp4_v_b_40')
// (5, 20, 'sp4_v_b_29')
// (5, 21, 'sp4_v_b_16')
// (5, 22, 'sp4_v_b_5')
// (6, 14, 'sp4_h_r_47')
// (7, 14, 'sp4_h_l_47')
// (7, 14, 'sp4_h_r_6')
// (8, 14, 'sp4_h_r_19')
// (9, 14, 'sp4_h_r_30')
// (10, 14, 'sp4_h_r_43')
// (10, 15, 'sp4_r_v_b_46')
// (10, 16, 'sp4_r_v_b_35')
// (10, 17, 'sp4_r_v_b_22')
// (10, 18, 'sp4_r_v_b_11')
// (10, 19, 'sp4_r_v_b_39')
// (10, 20, 'local_g0_2')
// (10, 20, 'lutff_5/in_1')
// (10, 20, 'sp4_r_v_b_26')
// (10, 21, 'sp4_r_v_b_15')
// (10, 22, 'sp4_r_v_b_2')
// (11, 14, 'sp4_h_l_43')
// (11, 14, 'sp4_v_t_46')
// (11, 15, 'sp4_v_b_46')
// (11, 16, 'sp4_v_b_35')
// (11, 17, 'sp4_v_b_22')
// (11, 18, 'sp4_v_b_11')
// (11, 18, 'sp4_v_t_39')
// (11, 19, 'sp4_v_b_39')
// (11, 20, 'local_g3_2')
// (11, 20, 'lutff_3/in_0')
// (11, 20, 'lutff_4/in_1')
// (11, 20, 'lutff_6/in_1')
// (11, 20, 'sp4_v_b_26')
// (11, 21, 'local_g1_7')
// (11, 21, 'lutff_2/in_2')
// (11, 21, 'lutff_4/in_2')
// (11, 21, 'sp4_v_b_15')
// (11, 22, 'sp4_v_b_2')

wire n81;
// (0, 10, 'sp4_r_v_b_45')
// (0, 11, 'sp4_r_v_b_32')
// (0, 12, 'sp4_r_v_b_21')
// (0, 13, 'sp4_r_v_b_8')
// (1, 9, 'sp4_v_t_45')
// (1, 10, 'sp4_v_b_45')
// (1, 11, 'sp4_v_b_32')
// (1, 12, 'local_g0_5')
// (1, 12, 'lutff_5/in_0')
// (1, 12, 'sp4_v_b_21')
// (1, 13, 'sp4_h_r_8')
// (1, 13, 'sp4_v_b_8')
// (2, 13, 'local_g1_5')
// (2, 13, 'lutff_2/in_0')
// (2, 13, 'sp4_h_r_21')
// (3, 10, 'neigh_op_tnr_5')
// (3, 11, 'neigh_op_rgt_5')
// (3, 12, 'neigh_op_bnr_5')
// (3, 13, 'sp4_h_r_32')
// (4, 10, 'neigh_op_top_5')
// (4, 10, 'sp4_r_v_b_38')
// (4, 11, 'lutff_5/out')
// (4, 11, 'sp4_r_v_b_27')
// (4, 12, 'neigh_op_bot_5')
// (4, 12, 'sp4_r_v_b_14')
// (4, 13, 'sp4_h_r_45')
// (4, 13, 'sp4_r_v_b_3')
// (5, 9, 'sp4_v_t_38')
// (5, 10, 'neigh_op_tnl_5')
// (5, 10, 'sp4_v_b_38')
// (5, 11, 'neigh_op_lft_5')
// (5, 11, 'sp4_v_b_27')
// (5, 12, 'neigh_op_bnl_5')
// (5, 12, 'sp4_v_b_14')
// (5, 13, 'sp4_h_l_45')
// (5, 13, 'sp4_v_b_3')

wire n82;
// (0, 11, 'neigh_op_tnr_0')
// (0, 12, 'neigh_op_rgt_0')
// (0, 13, 'neigh_op_bnr_0')
// (1, 11, 'neigh_op_top_0')
// (1, 12, 'lutff_0/out')
// (1, 13, 'neigh_op_bot_0')
// (2, 11, 'local_g2_0')
// (2, 11, 'lutff_1/in_1')
// (2, 11, 'neigh_op_tnl_0')
// (2, 12, 'neigh_op_lft_0')
// (2, 13, 'neigh_op_bnl_0')

wire n83;
// (0, 11, 'neigh_op_tnr_1')
// (0, 12, 'neigh_op_rgt_1')
// (0, 13, 'neigh_op_bnr_1')
// (1, 9, 'sp4_r_v_b_38')
// (1, 10, 'sp4_r_v_b_27')
// (1, 11, 'neigh_op_top_1')
// (1, 11, 'sp4_r_v_b_14')
// (1, 12, 'lutff_1/out')
// (1, 12, 'sp4_r_v_b_3')
// (1, 13, 'neigh_op_bot_1')
// (2, 8, 'local_g1_0')
// (2, 8, 'lutff_6/in_3')
// (2, 8, 'sp4_h_r_8')
// (2, 8, 'sp4_v_t_38')
// (2, 9, 'sp4_v_b_38')
// (2, 10, 'sp4_v_b_27')
// (2, 11, 'neigh_op_tnl_1')
// (2, 11, 'sp4_v_b_14')
// (2, 12, 'neigh_op_lft_1')
// (2, 12, 'sp4_v_b_3')
// (2, 13, 'neigh_op_bnl_1')
// (3, 8, 'local_g0_5')
// (3, 8, 'lutff_3/in_2')
// (3, 8, 'lutff_4/in_3')
// (3, 8, 'lutff_5/in_2')
// (3, 8, 'lutff_7/in_2')
// (3, 8, 'sp4_h_r_21')
// (4, 8, 'sp4_h_r_32')
// (5, 8, 'sp4_h_r_45')
// (6, 8, 'sp4_h_l_45')

wire n84;
// (0, 11, 'neigh_op_tnr_2')
// (0, 12, 'neigh_op_rgt_2')
// (0, 13, 'neigh_op_bnr_2')
// (1, 11, 'neigh_op_top_2')
// (1, 12, 'local_g1_2')
// (1, 12, 'lutff_1/in_0')
// (1, 12, 'lutff_2/out')
// (1, 13, 'neigh_op_bot_2')
// (2, 11, 'neigh_op_tnl_2')
// (2, 12, 'neigh_op_lft_2')
// (2, 13, 'neigh_op_bnl_2')

reg io_4_31_0 = 0;
// (0, 11, 'neigh_op_tnr_3')
// (0, 12, 'neigh_op_rgt_3')
// (0, 12, 'sp4_h_r_11')
// (0, 13, 'neigh_op_bnr_3')
// (1, 11, 'neigh_op_top_3')
// (1, 12, 'local_g0_3')
// (1, 12, 'local_g1_3')
// (1, 12, 'lutff_2/in_1')
// (1, 12, 'lutff_3/in_3')
// (1, 12, 'lutff_3/out')
// (1, 12, 'sp4_h_r_22')
// (1, 12, 'sp4_r_v_b_39')
// (1, 13, 'neigh_op_bot_3')
// (1, 13, 'sp4_r_v_b_26')
// (1, 14, 'sp4_r_v_b_15')
// (1, 15, 'local_g1_2')
// (1, 15, 'lutff_2/in_1')
// (1, 15, 'sp4_r_v_b_2')
// (1, 16, 'sp4_r_v_b_39')
// (1, 17, 'sp4_r_v_b_26')
// (1, 18, 'sp4_r_v_b_15')
// (1, 19, 'sp4_r_v_b_2')
// (2, 11, 'neigh_op_tnl_3')
// (2, 11, 'sp4_v_t_39')
// (2, 12, 'neigh_op_lft_3')
// (2, 12, 'sp4_h_r_35')
// (2, 12, 'sp4_v_b_39')
// (2, 13, 'neigh_op_bnl_3')
// (2, 13, 'sp4_v_b_26')
// (2, 14, 'sp4_v_b_15')
// (2, 15, 'sp4_v_b_2')
// (2, 15, 'sp4_v_t_39')
// (2, 16, 'sp4_v_b_39')
// (2, 17, 'local_g2_2')
// (2, 17, 'lutff_7/in_1')
// (2, 17, 'sp4_v_b_26')
// (2, 18, 'sp4_v_b_15')
// (2, 19, 'sp4_v_b_2')
// (3, 12, 'sp4_h_r_46')
// (3, 13, 'sp4_r_v_b_41')
// (3, 14, 'sp4_r_v_b_28')
// (3, 15, 'sp4_r_v_b_17')
// (3, 16, 'local_g1_4')
// (3, 16, 'lutff_2/in_1')
// (3, 16, 'sp4_r_v_b_4')
// (3, 17, 'sp4_r_v_b_42')
// (3, 18, 'sp4_r_v_b_31')
// (3, 19, 'sp4_r_v_b_18')
// (3, 20, 'sp4_r_v_b_7')
// (3, 21, 'sp4_r_v_b_47')
// (3, 22, 'sp4_r_v_b_34')
// (3, 23, 'sp4_r_v_b_23')
// (3, 24, 'sp4_r_v_b_10')
// (3, 25, 'sp4_r_v_b_43')
// (3, 26, 'sp4_r_v_b_30')
// (3, 27, 'sp4_r_v_b_19')
// (3, 28, 'sp4_r_v_b_6')
// (3, 29, 'sp4_r_v_b_39')
// (3, 30, 'sp4_r_v_b_26')
// (4, 12, 'sp4_h_l_46')
// (4, 12, 'sp4_v_t_41')
// (4, 13, 'sp4_v_b_41')
// (4, 14, 'sp4_v_b_28')
// (4, 15, 'sp4_v_b_17')
// (4, 16, 'sp4_h_r_4')
// (4, 16, 'sp4_v_b_4')
// (4, 16, 'sp4_v_t_42')
// (4, 17, 'sp4_v_b_42')
// (4, 18, 'sp4_v_b_31')
// (4, 19, 'sp4_v_b_18')
// (4, 20, 'sp4_v_b_7')
// (4, 20, 'sp4_v_t_47')
// (4, 21, 'sp4_v_b_47')
// (4, 22, 'sp4_v_b_34')
// (4, 23, 'sp4_v_b_23')
// (4, 24, 'sp4_v_b_10')
// (4, 24, 'sp4_v_t_43')
// (4, 25, 'sp4_v_b_43')
// (4, 26, 'sp4_v_b_30')
// (4, 27, 'sp4_v_b_19')
// (4, 28, 'sp4_v_b_6')
// (4, 28, 'sp4_v_t_39')
// (4, 29, 'sp4_v_b_39')
// (4, 30, 'sp4_v_b_26')
// (4, 31, 'io_0/D_OUT_0')
// (4, 31, 'io_0/PAD')
// (4, 31, 'local_g1_7')
// (4, 31, 'span4_vert_15')
// (5, 16, 'local_g1_1')
// (5, 16, 'lutff_6/in_2')
// (5, 16, 'sp4_h_r_17')
// (6, 16, 'sp4_h_r_28')
// (7, 16, 'sp4_h_r_41')
// (8, 16, 'sp4_h_l_41')

wire n86;
// (0, 11, 'neigh_op_tnr_4')
// (0, 12, 'neigh_op_rgt_4')
// (0, 13, 'neigh_op_bnr_4')
// (1, 9, 'sp4_r_v_b_44')
// (1, 10, 'sp4_r_v_b_33')
// (1, 11, 'neigh_op_top_4')
// (1, 11, 'sp4_r_v_b_20')
// (1, 12, 'lutff_4/out')
// (1, 12, 'sp4_r_v_b_9')
// (1, 13, 'neigh_op_bot_4')
// (2, 8, 'sp4_v_t_44')
// (2, 9, 'sp4_v_b_44')
// (2, 10, 'local_g3_1')
// (2, 10, 'lutff_4/in_0')
// (2, 10, 'sp4_v_b_33')
// (2, 11, 'neigh_op_tnl_4')
// (2, 11, 'sp4_v_b_20')
// (2, 12, 'neigh_op_lft_4')
// (2, 12, 'sp4_v_b_9')
// (2, 13, 'neigh_op_bnl_4')

reg n87 = 0;
// (0, 11, 'neigh_op_tnr_5')
// (0, 12, 'neigh_op_rgt_5')
// (0, 12, 'sp4_h_r_15')
// (0, 12, 'sp4_r_v_b_42')
// (0, 13, 'neigh_op_bnr_5')
// (0, 13, 'sp4_r_v_b_31')
// (0, 14, 'sp4_r_v_b_18')
// (0, 15, 'sp4_r_v_b_7')
// (1, 11, 'neigh_op_top_5')
// (1, 11, 'sp4_v_t_42')
// (1, 12, 'local_g1_5')
// (1, 12, 'lutff_5/in_3')
// (1, 12, 'lutff_5/out')
// (1, 12, 'sp4_h_r_10')
// (1, 12, 'sp4_h_r_26')
// (1, 12, 'sp4_v_b_42')
// (1, 13, 'local_g0_5')
// (1, 13, 'lutff_4/in_3')
// (1, 13, 'neigh_op_bot_5')
// (1, 13, 'sp4_v_b_31')
// (1, 14, 'sp4_v_b_18')
// (1, 15, 'sp4_h_r_1')
// (1, 15, 'sp4_v_b_7')
// (2, 9, 'sp4_r_v_b_45')
// (2, 10, 'sp4_r_v_b_32')
// (2, 11, 'neigh_op_tnl_5')
// (2, 11, 'sp4_r_v_b_21')
// (2, 12, 'neigh_op_lft_5')
// (2, 12, 'sp4_h_r_23')
// (2, 12, 'sp4_h_r_39')
// (2, 12, 'sp4_r_v_b_8')
// (2, 13, 'neigh_op_bnl_5')
// (2, 15, 'sp4_h_r_12')
// (3, 8, 'sp4_v_t_45')
// (3, 9, 'sp4_v_b_45')
// (3, 10, 'sp4_v_b_32')
// (3, 11, 'local_g0_5')
// (3, 11, 'lutff_3/in_2')
// (3, 11, 'sp4_v_b_21')
// (3, 12, 'sp4_h_l_39')
// (3, 12, 'sp4_h_r_34')
// (3, 12, 'sp4_v_b_8')
// (3, 15, 'sp4_h_r_25')
// (4, 9, 'sp4_r_v_b_47')
// (4, 10, 'sp4_r_v_b_34')
// (4, 11, 'local_g3_7')
// (4, 11, 'lutff_7/in_1')
// (4, 11, 'sp4_r_v_b_23')
// (4, 12, 'sp4_h_r_47')
// (4, 12, 'sp4_r_v_b_10')
// (4, 15, 'local_g3_4')
// (4, 15, 'lutff_0/in_1')
// (4, 15, 'sp4_h_r_36')
// (5, 8, 'sp4_v_t_47')
// (5, 9, 'sp4_v_b_47')
// (5, 10, 'sp4_v_b_34')
// (5, 11, 'sp4_v_b_23')
// (5, 12, 'sp4_h_l_47')
// (5, 12, 'sp4_v_b_10')
// (5, 15, 'sp4_h_l_36')

wire n88;
// (0, 11, 'neigh_op_tnr_6')
// (0, 12, 'neigh_op_rgt_6')
// (0, 13, 'neigh_op_bnr_6')
// (1, 11, 'neigh_op_top_6')
// (1, 12, 'lutff_6/out')
// (1, 12, 'sp4_r_v_b_45')
// (1, 13, 'neigh_op_bot_6')
// (1, 13, 'sp4_r_v_b_32')
// (1, 14, 'sp4_r_v_b_21')
// (1, 15, 'sp4_r_v_b_8')
// (2, 11, 'neigh_op_tnl_6')
// (2, 11, 'sp4_h_r_8')
// (2, 11, 'sp4_v_t_45')
// (2, 12, 'neigh_op_lft_6')
// (2, 12, 'sp4_v_b_45')
// (2, 13, 'neigh_op_bnl_6')
// (2, 13, 'sp4_v_b_32')
// (2, 14, 'sp4_v_b_21')
// (2, 15, 'sp4_v_b_8')
// (3, 11, 'sp4_h_r_21')
// (4, 11, 'local_g2_0')
// (4, 11, 'local_g3_0')
// (4, 11, 'lutff_4/in_3')
// (4, 11, 'lutff_5/in_1')
// (4, 11, 'lutff_6/in_1')
// (4, 11, 'sp4_h_r_32')
// (5, 11, 'sp4_h_r_45')
// (6, 11, 'sp4_h_l_45')

wire n89;
// (0, 11, 'neigh_op_tnr_7')
// (0, 12, 'neigh_op_rgt_7')
// (0, 13, 'neigh_op_bnr_7')
// (1, 11, 'local_g0_7')
// (1, 11, 'lutff_2/in_3')
// (1, 11, 'neigh_op_top_7')
// (1, 12, 'lutff_7/out')
// (1, 13, 'neigh_op_bot_7')
// (2, 11, 'neigh_op_tnl_7')
// (2, 12, 'neigh_op_lft_7')
// (2, 13, 'neigh_op_bnl_7')

reg n90 = 0;
// (0, 11, 'sp4_h_r_10')
// (1, 10, 'sp4_r_v_b_40')
// (1, 11, 'sp4_h_r_23')
// (1, 11, 'sp4_r_v_b_29')
// (1, 12, 'sp4_r_v_b_16')
// (1, 13, 'sp4_r_v_b_5')
// (2, 9, 'sp4_h_r_11')
// (2, 9, 'sp4_v_t_40')
// (2, 10, 'sp4_v_b_40')
// (2, 11, 'local_g3_2')
// (2, 11, 'lutff_3/in_2')
// (2, 11, 'sp4_h_r_34')
// (2, 11, 'sp4_v_b_29')
// (2, 12, 'local_g0_0')
// (2, 12, 'lutff_0/in_2')
// (2, 12, 'sp4_v_b_16')
// (2, 13, 'sp4_v_b_5')
// (3, 9, 'sp4_h_r_22')
// (3, 11, 'sp4_h_r_47')
// (4, 9, 'sp4_h_r_35')
// (4, 11, 'sp4_h_l_47')
// (4, 11, 'sp4_h_r_7')
// (5, 9, 'sp4_h_r_46')
// (5, 11, 'sp4_h_r_18')
// (6, 8, 'neigh_op_tnr_7')
// (6, 9, 'neigh_op_rgt_7')
// (6, 9, 'sp4_h_l_46')
// (6, 9, 'sp4_h_r_3')
// (6, 10, 'neigh_op_bnr_7')
// (6, 11, 'sp4_h_r_31')
// (7, 8, 'neigh_op_top_7')
// (7, 8, 'sp4_r_v_b_42')
// (7, 9, 'lutff_7/out')
// (7, 9, 'sp4_h_r_14')
// (7, 9, 'sp4_r_v_b_31')
// (7, 10, 'neigh_op_bot_7')
// (7, 10, 'sp4_r_v_b_18')
// (7, 11, 'sp4_h_r_42')
// (7, 11, 'sp4_r_v_b_7')
// (8, 7, 'sp4_v_t_42')
// (8, 8, 'neigh_op_tnl_7')
// (8, 8, 'sp4_v_b_42')
// (8, 9, 'neigh_op_lft_7')
// (8, 9, 'sp4_h_r_27')
// (8, 9, 'sp4_v_b_31')
// (8, 10, 'neigh_op_bnl_7')
// (8, 10, 'sp4_v_b_18')
// (8, 11, 'sp4_h_l_42')
// (8, 11, 'sp4_v_b_7')
// (9, 9, 'sp4_h_r_38')
// (10, 9, 'sp4_h_l_38')

reg n91 = 0;
// (0, 11, 'sp4_h_r_6')
// (1, 10, 'neigh_op_tnr_7')
// (1, 11, 'neigh_op_rgt_7')
// (1, 11, 'sp4_h_r_19')
// (1, 11, 'sp4_r_v_b_46')
// (1, 12, 'neigh_op_bnr_7')
// (1, 12, 'sp4_r_v_b_35')
// (1, 13, 'sp4_r_v_b_22')
// (1, 14, 'sp4_r_v_b_11')
// (2, 10, 'neigh_op_top_7')
// (2, 10, 'sp4_v_t_46')
// (2, 11, 'local_g2_7')
// (2, 11, 'local_g3_7')
// (2, 11, 'lutff_4/in_3')
// (2, 11, 'lutff_7/in_1')
// (2, 11, 'lutff_7/out')
// (2, 11, 'sp4_h_r_30')
// (2, 11, 'sp4_r_v_b_47')
// (2, 11, 'sp4_v_b_46')
// (2, 12, 'neigh_op_bot_7')
// (2, 12, 'sp4_r_v_b_34')
// (2, 12, 'sp4_v_b_35')
// (2, 13, 'sp4_r_v_b_23')
// (2, 13, 'sp4_v_b_22')
// (2, 14, 'local_g1_3')
// (2, 14, 'lutff_4/in_0')
// (2, 14, 'lutff_5/in_3')
// (2, 14, 'sp4_r_v_b_10')
// (2, 14, 'sp4_v_b_11')
// (2, 15, 'sp4_r_v_b_47')
// (2, 16, 'sp4_r_v_b_34')
// (2, 17, 'sp4_r_v_b_23')
// (2, 18, 'sp4_r_v_b_10')
// (3, 10, 'neigh_op_tnl_7')
// (3, 10, 'sp4_v_t_47')
// (3, 11, 'neigh_op_lft_7')
// (3, 11, 'sp4_h_r_43')
// (3, 11, 'sp4_v_b_47')
// (3, 12, 'neigh_op_bnl_7')
// (3, 12, 'sp4_r_v_b_46')
// (3, 12, 'sp4_v_b_34')
// (3, 13, 'sp4_r_v_b_35')
// (3, 13, 'sp4_v_b_23')
// (3, 14, 'sp4_r_v_b_22')
// (3, 14, 'sp4_v_b_10')
// (3, 14, 'sp4_v_t_47')
// (3, 15, 'local_g2_3')
// (3, 15, 'lutff_6/in_1')
// (3, 15, 'sp4_r_v_b_11')
// (3, 15, 'sp4_v_b_47')
// (3, 16, 'local_g3_2')
// (3, 16, 'lutff_4/in_3')
// (3, 16, 'sp4_r_v_b_46')
// (3, 16, 'sp4_v_b_34')
// (3, 17, 'sp4_r_v_b_35')
// (3, 17, 'sp4_v_b_23')
// (3, 18, 'sp4_r_v_b_22')
// (3, 18, 'sp4_v_b_10')
// (3, 19, 'sp4_r_v_b_11')
// (4, 11, 'sp4_h_l_43')
// (4, 11, 'sp4_v_t_46')
// (4, 12, 'sp4_v_b_46')
// (4, 13, 'sp4_v_b_35')
// (4, 14, 'sp4_v_b_22')
// (4, 15, 'sp4_v_b_11')
// (4, 15, 'sp4_v_t_46')
// (4, 16, 'local_g2_6')
// (4, 16, 'lutff_2/in_2')
// (4, 16, 'sp4_v_b_46')
// (4, 17, 'sp4_v_b_35')
// (4, 18, 'sp4_v_b_22')
// (4, 19, 'sp4_v_b_11')

wire n92;
// (0, 11, 'sp4_r_v_b_37')
// (0, 12, 'sp4_r_v_b_24')
// (0, 13, 'sp4_r_v_b_13')
// (0, 14, 'sp4_r_v_b_0')
// (1, 10, 'sp4_v_t_37')
// (1, 11, 'local_g3_5')
// (1, 11, 'lutff_6/in_0')
// (1, 11, 'sp4_v_b_37')
// (1, 12, 'local_g3_0')
// (1, 12, 'lutff_7/in_0')
// (1, 12, 'sp4_v_b_24')
// (1, 13, 'sp4_v_b_13')
// (1, 14, 'sp4_h_r_0')
// (1, 14, 'sp4_v_b_0')
// (2, 11, 'sp4_r_v_b_45')
// (2, 12, 'sp4_r_v_b_32')
// (2, 13, 'neigh_op_tnr_4')
// (2, 13, 'sp4_r_v_b_21')
// (2, 14, 'neigh_op_rgt_4')
// (2, 14, 'sp4_h_r_13')
// (2, 14, 'sp4_r_v_b_8')
// (2, 15, 'neigh_op_bnr_4')
// (3, 10, 'local_g1_1')
// (3, 10, 'lutff_4/in_2')
// (3, 10, 'sp4_h_r_1')
// (3, 10, 'sp4_v_t_45')
// (3, 11, 'sp4_v_b_45')
// (3, 12, 'sp4_v_b_32')
// (3, 13, 'neigh_op_top_4')
// (3, 13, 'sp4_v_b_21')
// (3, 14, 'lutff_4/out')
// (3, 14, 'sp4_h_r_24')
// (3, 14, 'sp4_v_b_8')
// (3, 15, 'neigh_op_bot_4')
// (4, 10, 'sp4_h_r_12')
// (4, 13, 'neigh_op_tnl_4')
// (4, 14, 'neigh_op_lft_4')
// (4, 14, 'sp4_h_r_37')
// (4, 15, 'local_g2_4')
// (4, 15, 'lutff_1/in_3')
// (4, 15, 'neigh_op_bnl_4')
// (5, 10, 'sp4_h_r_25')
// (5, 14, 'sp4_h_l_37')
// (6, 10, 'sp4_h_r_36')
// (7, 10, 'sp4_h_l_36')

reg n93 = 0;
// (0, 11, 'sp4_r_v_b_42')
// (0, 12, 'sp4_r_v_b_31')
// (0, 13, 'sp4_r_v_b_18')
// (0, 14, 'sp4_r_v_b_7')
// (0, 15, 'sp4_r_v_b_47')
// (0, 16, 'sp4_r_v_b_34')
// (0, 17, 'sp4_r_v_b_23')
// (0, 18, 'sp4_r_v_b_10')
// (1, 8, 'sp4_r_v_b_36')
// (1, 9, 'neigh_op_tnr_6')
// (1, 9, 'sp4_r_v_b_25')
// (1, 9, 'sp4_r_v_b_41')
// (1, 10, 'neigh_op_rgt_6')
// (1, 10, 'sp4_h_r_1')
// (1, 10, 'sp4_r_v_b_12')
// (1, 10, 'sp4_r_v_b_28')
// (1, 10, 'sp4_r_v_b_44')
// (1, 10, 'sp4_v_t_42')
// (1, 11, 'neigh_op_bnr_6')
// (1, 11, 'sp4_r_v_b_1')
// (1, 11, 'sp4_r_v_b_17')
// (1, 11, 'sp4_r_v_b_33')
// (1, 11, 'sp4_v_b_42')
// (1, 12, 'local_g1_4')
// (1, 12, 'lutff_3/in_0')
// (1, 12, 'sp4_r_v_b_20')
// (1, 12, 'sp4_r_v_b_4')
// (1, 12, 'sp4_v_b_31')
// (1, 13, 'sp4_r_v_b_41')
// (1, 13, 'sp4_r_v_b_9')
// (1, 13, 'sp4_v_b_18')
// (1, 14, 'sp4_r_v_b_28')
// (1, 14, 'sp4_r_v_b_40')
// (1, 14, 'sp4_v_b_7')
// (1, 14, 'sp4_v_t_47')
// (1, 15, 'local_g3_1')
// (1, 15, 'lutff_3/in_1')
// (1, 15, 'sp4_r_v_b_17')
// (1, 15, 'sp4_r_v_b_29')
// (1, 15, 'sp4_v_b_47')
// (1, 16, 'sp4_r_v_b_16')
// (1, 16, 'sp4_r_v_b_4')
// (1, 16, 'sp4_v_b_34')
// (1, 17, 'sp4_r_v_b_41')
// (1, 17, 'sp4_r_v_b_42')
// (1, 17, 'sp4_r_v_b_5')
// (1, 17, 'sp4_v_b_23')
// (1, 18, 'local_g1_2')
// (1, 18, 'lutff_5/in_0')
// (1, 18, 'sp4_r_v_b_28')
// (1, 18, 'sp4_r_v_b_31')
// (1, 18, 'sp4_r_v_b_40')
// (1, 18, 'sp4_v_b_10')
// (1, 19, 'local_g3_2')
// (1, 19, 'lutff_6/in_3')
// (1, 19, 'sp4_r_v_b_17')
// (1, 19, 'sp4_r_v_b_18')
// (1, 19, 'sp4_r_v_b_29')
// (1, 20, 'sp4_r_v_b_16')
// (1, 20, 'sp4_r_v_b_4')
// (1, 20, 'sp4_r_v_b_7')
// (1, 21, 'sp4_r_v_b_5')
// (2, 7, 'sp4_h_r_6')
// (2, 7, 'sp4_v_t_36')
// (2, 8, 'sp4_v_b_36')
// (2, 8, 'sp4_v_t_41')
// (2, 9, 'neigh_op_top_6')
// (2, 9, 'sp4_v_b_25')
// (2, 9, 'sp4_v_b_41')
// (2, 9, 'sp4_v_t_44')
// (2, 10, 'local_g0_6')
// (2, 10, 'lutff_4/in_2')
// (2, 10, 'lutff_6/in_2')
// (2, 10, 'lutff_6/out')
// (2, 10, 'sp4_h_r_12')
// (2, 10, 'sp4_v_b_12')
// (2, 10, 'sp4_v_b_28')
// (2, 10, 'sp4_v_b_44')
// (2, 11, 'local_g0_6')
// (2, 11, 'lutff_4/in_2')
// (2, 11, 'neigh_op_bot_6')
// (2, 11, 'sp4_v_b_1')
// (2, 11, 'sp4_v_b_17')
// (2, 11, 'sp4_v_b_33')
// (2, 12, 'sp4_v_b_20')
// (2, 12, 'sp4_v_b_4')
// (2, 12, 'sp4_v_t_41')
// (2, 13, 'sp4_v_b_41')
// (2, 13, 'sp4_v_b_9')
// (2, 13, 'sp4_v_t_40')
// (2, 14, 'sp4_v_b_28')
// (2, 14, 'sp4_v_b_40')
// (2, 15, 'sp4_v_b_17')
// (2, 15, 'sp4_v_b_29')
// (2, 16, 'sp4_v_b_16')
// (2, 16, 'sp4_v_b_4')
// (2, 16, 'sp4_v_t_41')
// (2, 16, 'sp4_v_t_42')
// (2, 17, 'sp4_v_b_41')
// (2, 17, 'sp4_v_b_42')
// (2, 17, 'sp4_v_b_5')
// (2, 17, 'sp4_v_t_40')
// (2, 18, 'sp4_v_b_28')
// (2, 18, 'sp4_v_b_31')
// (2, 18, 'sp4_v_b_40')
// (2, 19, 'local_g0_1')
// (2, 19, 'lutff_5/in_2')
// (2, 19, 'sp4_v_b_17')
// (2, 19, 'sp4_v_b_18')
// (2, 19, 'sp4_v_b_29')
// (2, 20, 'local_g0_0')
// (2, 20, 'lutff_1/in_1')
// (2, 20, 'lutff_4/in_0')
// (2, 20, 'lutff_5/in_1')
// (2, 20, 'sp4_v_b_16')
// (2, 20, 'sp4_v_b_4')
// (2, 20, 'sp4_v_b_7')
// (2, 21, 'sp4_v_b_5')
// (3, 7, 'local_g0_3')
// (3, 7, 'lutff_1/in_2')
// (3, 7, 'sp4_h_r_19')
// (3, 9, 'neigh_op_tnl_6')
// (3, 10, 'neigh_op_lft_6')
// (3, 10, 'sp4_h_r_25')
// (3, 11, 'neigh_op_bnl_6')
// (4, 7, 'sp4_h_r_30')
// (4, 10, 'sp4_h_r_36')
// (4, 11, 'sp4_r_v_b_43')
// (4, 12, 'sp4_r_v_b_30')
// (4, 13, 'sp4_r_v_b_19')
// (4, 14, 'sp4_r_v_b_6')
// (4, 15, 'sp4_r_v_b_43')
// (4, 16, 'sp4_r_v_b_30')
// (4, 17, 'sp4_r_v_b_19')
// (4, 18, 'sp4_r_v_b_6')
// (5, 7, 'sp4_h_r_43')
// (5, 10, 'sp4_h_l_36')
// (5, 10, 'sp4_v_t_43')
// (5, 11, 'sp4_v_b_43')
// (5, 12, 'sp4_v_b_30')
// (5, 13, 'sp4_v_b_19')
// (5, 14, 'sp4_v_b_6')
// (5, 14, 'sp4_v_t_43')
// (5, 15, 'sp4_v_b_43')
// (5, 16, 'sp4_v_b_30')
// (5, 17, 'local_g0_3')
// (5, 17, 'lutff_1/in_2')
// (5, 17, 'sp4_v_b_19')
// (5, 18, 'sp4_v_b_6')
// (6, 7, 'sp4_h_l_43')

reg n94 = 0;
// (0, 12, 'neigh_op_tnr_1')
// (0, 13, 'neigh_op_rgt_1')
// (0, 14, 'neigh_op_bnr_1')
// (1, 12, 'neigh_op_top_1')
// (1, 13, 'local_g2_1')
// (1, 13, 'lutff_1/in_2')
// (1, 13, 'lutff_1/out')
// (1, 14, 'neigh_op_bot_1')
// (2, 12, 'neigh_op_tnl_1')
// (2, 13, 'local_g0_1')
// (2, 13, 'lutff_1/in_2')
// (2, 13, 'neigh_op_lft_1')
// (2, 14, 'neigh_op_bnl_1')

reg n95 = 0;
// (0, 12, 'neigh_op_tnr_2')
// (0, 13, 'neigh_op_rgt_2')
// (0, 13, 'sp4_h_r_9')
// (0, 14, 'neigh_op_bnr_2')
// (1, 12, 'neigh_op_top_2')
// (1, 13, 'local_g2_2')
// (1, 13, 'lutff_2/in_0')
// (1, 13, 'lutff_2/out')
// (1, 13, 'sp4_h_r_20')
// (1, 14, 'neigh_op_bot_2')
// (2, 12, 'neigh_op_tnl_2')
// (2, 13, 'local_g3_1')
// (2, 13, 'lutff_1/in_1')
// (2, 13, 'neigh_op_lft_2')
// (2, 13, 'sp4_h_r_33')
// (2, 14, 'neigh_op_bnl_2')
// (3, 13, 'sp4_h_r_44')
// (4, 13, 'sp4_h_l_44')

reg n96 = 0;
// (0, 12, 'neigh_op_tnr_3')
// (0, 13, 'neigh_op_rgt_3')
// (0, 14, 'neigh_op_bnr_3')
// (1, 11, 'sp4_r_v_b_47')
// (1, 12, 'neigh_op_top_3')
// (1, 12, 'sp4_r_v_b_34')
// (1, 13, 'local_g1_3')
// (1, 13, 'lutff_0/in_2')
// (1, 13, 'lutff_1/in_3')
// (1, 13, 'lutff_3/in_3')
// (1, 13, 'lutff_3/out')
// (1, 13, 'sp4_r_v_b_23')
// (1, 14, 'neigh_op_bot_3')
// (1, 14, 'sp4_r_v_b_10')
// (2, 10, 'sp4_v_t_47')
// (2, 11, 'sp4_v_b_47')
// (2, 12, 'neigh_op_tnl_3')
// (2, 12, 'sp4_v_b_34')
// (2, 13, 'local_g1_7')
// (2, 13, 'lutff_1/in_3')
// (2, 13, 'neigh_op_lft_3')
// (2, 13, 'sp4_v_b_23')
// (2, 14, 'neigh_op_bnl_3')
// (2, 14, 'sp4_v_b_10')

wire n97;
// (0, 12, 'neigh_op_tnr_4')
// (0, 13, 'neigh_op_rgt_4')
// (0, 14, 'neigh_op_bnr_4')
// (1, 12, 'neigh_op_top_4')
// (1, 13, 'lutff_4/out')
// (1, 14, 'neigh_op_bot_4')
// (2, 12, 'neigh_op_tnl_4')
// (2, 13, 'local_g0_4')
// (2, 13, 'lutff_6/in_2')
// (2, 13, 'neigh_op_lft_4')
// (2, 14, 'neigh_op_bnl_4')

wire n98;
// (0, 12, 'neigh_op_tnr_5')
// (0, 13, 'neigh_op_rgt_5')
// (0, 14, 'neigh_op_bnr_5')
// (1, 12, 'neigh_op_top_5')
// (1, 13, 'lutff_5/out')
// (1, 13, 'sp4_r_v_b_43')
// (1, 14, 'neigh_op_bot_5')
// (1, 14, 'sp4_r_v_b_30')
// (1, 15, 'sp4_r_v_b_19')
// (1, 16, 'sp4_r_v_b_6')
// (2, 12, 'neigh_op_tnl_5')
// (2, 12, 'sp4_h_r_6')
// (2, 12, 'sp4_v_t_43')
// (2, 13, 'neigh_op_lft_5')
// (2, 13, 'sp4_v_b_43')
// (2, 14, 'neigh_op_bnl_5')
// (2, 14, 'sp4_v_b_30')
// (2, 15, 'sp4_v_b_19')
// (2, 16, 'sp4_v_b_6')
// (3, 12, 'local_g1_3')
// (3, 12, 'lutff_global/cen')
// (3, 12, 'sp4_h_r_19')
// (4, 12, 'sp4_h_r_30')
// (5, 12, 'sp4_h_r_43')
// (6, 12, 'sp4_h_l_43')

wire n99;
// (0, 12, 'neigh_op_tnr_6')
// (0, 13, 'neigh_op_rgt_6')
// (0, 14, 'neigh_op_bnr_6')
// (1, 12, 'neigh_op_top_6')
// (1, 13, 'local_g3_6')
// (1, 13, 'lutff_1/in_0')
// (1, 13, 'lutff_2/in_1')
// (1, 13, 'lutff_3/in_0')
// (1, 13, 'lutff_6/out')
// (1, 14, 'local_g0_6')
// (1, 14, 'lutff_0/in_0')
// (1, 14, 'lutff_3/in_1')
// (1, 14, 'lutff_6/in_2')
// (1, 14, 'neigh_op_bot_6')
// (2, 12, 'neigh_op_tnl_6')
// (2, 13, 'neigh_op_lft_6')
// (2, 14, 'neigh_op_bnl_6')

wire n100;
// (0, 12, 'neigh_op_tnr_7')
// (0, 13, 'neigh_op_rgt_7')
// (0, 14, 'neigh_op_bnr_7')
// (1, 12, 'neigh_op_top_7')
// (1, 13, 'lutff_7/out')
// (1, 14, 'neigh_op_bot_7')
// (2, 12, 'local_g3_7')
// (2, 12, 'lutff_2/in_0')
// (2, 12, 'neigh_op_tnl_7')
// (2, 13, 'local_g0_7')
// (2, 13, 'lutff_0/in_1')
// (2, 13, 'neigh_op_lft_7')
// (2, 14, 'neigh_op_bnl_7')

reg n101 = 0;
// (0, 12, 'sp4_h_r_2')
// (1, 11, 'neigh_op_tnr_5')
// (1, 12, 'neigh_op_rgt_5')
// (1, 12, 'sp4_h_r_15')
// (1, 13, 'neigh_op_bnr_5')
// (2, 11, 'neigh_op_top_5')
// (2, 12, 'local_g3_5')
// (2, 12, 'lutff_5/in_1')
// (2, 12, 'lutff_5/out')
// (2, 12, 'sp4_h_r_26')
// (2, 13, 'neigh_op_bot_5')
// (3, 5, 'sp4_r_v_b_45')
// (3, 6, 'sp4_r_v_b_32')
// (3, 7, 'sp4_r_v_b_21')
// (3, 8, 'sp4_r_v_b_8')
// (3, 9, 'sp4_r_v_b_45')
// (3, 10, 'sp4_r_v_b_32')
// (3, 11, 'neigh_op_tnl_5')
// (3, 11, 'sp4_r_v_b_21')
// (3, 12, 'neigh_op_lft_5')
// (3, 12, 'sp4_h_r_39')
// (3, 12, 'sp4_r_v_b_8')
// (3, 13, 'neigh_op_bnl_5')
// (4, 4, 'sp4_v_t_45')
// (4, 5, 'local_g2_5')
// (4, 5, 'lutff_4/in_1')
// (4, 5, 'sp4_v_b_45')
// (4, 6, 'sp4_v_b_32')
// (4, 7, 'sp4_v_b_21')
// (4, 8, 'sp4_v_b_8')
// (4, 8, 'sp4_v_t_45')
// (4, 9, 'sp4_v_b_45')
// (4, 10, 'sp4_v_b_32')
// (4, 11, 'sp4_v_b_21')
// (4, 12, 'sp4_h_l_39')
// (4, 12, 'sp4_v_b_8')

wire n102;
// (0, 12, 'sp4_h_r_22')
// (1, 12, 'local_g3_3')
// (1, 12, 'lutff_6/in_2')
// (1, 12, 'sp4_h_r_35')
// (2, 9, 'sp4_r_v_b_46')
// (2, 10, 'neigh_op_tnr_3')
// (2, 10, 'sp4_r_v_b_35')
// (2, 11, 'neigh_op_rgt_3')
// (2, 11, 'sp4_r_v_b_22')
// (2, 12, 'neigh_op_bnr_3')
// (2, 12, 'sp4_h_r_46')
// (2, 12, 'sp4_r_v_b_11')
// (3, 8, 'sp4_v_t_46')
// (3, 9, 'sp4_v_b_46')
// (3, 10, 'neigh_op_top_3')
// (3, 10, 'sp4_v_b_35')
// (3, 11, 'lutff_3/out')
// (3, 11, 'sp4_h_r_6')
// (3, 11, 'sp4_v_b_22')
// (3, 12, 'neigh_op_bot_3')
// (3, 12, 'sp4_h_l_46')
// (3, 12, 'sp4_v_b_11')
// (4, 10, 'neigh_op_tnl_3')
// (4, 11, 'neigh_op_lft_3')
// (4, 11, 'sp4_h_r_19')
// (4, 12, 'neigh_op_bnl_3')
// (5, 11, 'sp4_h_r_30')
// (6, 11, 'sp4_h_r_43')
// (7, 11, 'sp4_h_l_43')
// (7, 11, 'sp4_h_r_6')
// (8, 11, 'sp4_h_r_19')
// (9, 11, 'sp4_h_r_30')
// (10, 11, 'sp4_h_r_43')
// (10, 12, 'sp4_r_v_b_43')
// (10, 13, 'sp4_r_v_b_30')
// (10, 14, 'sp4_r_v_b_19')
// (10, 15, 'sp4_r_v_b_6')
// (11, 11, 'sp4_h_l_43')
// (11, 11, 'sp4_v_t_43')
// (11, 12, 'local_g3_3')
// (11, 12, 'lutff_global/cen')
// (11, 12, 'sp4_v_b_43')
// (11, 13, 'sp4_v_b_30')
// (11, 14, 'sp4_v_b_19')
// (11, 15, 'sp4_v_b_6')

reg n103 = 0;
// (0, 12, 'sp4_h_r_4')
// (1, 11, 'neigh_op_tnr_6')
// (1, 11, 'sp4_r_v_b_41')
// (1, 12, 'neigh_op_rgt_6')
// (1, 12, 'sp4_h_r_17')
// (1, 12, 'sp4_r_v_b_28')
// (1, 12, 'sp4_r_v_b_44')
// (1, 13, 'neigh_op_bnr_6')
// (1, 13, 'sp4_r_v_b_17')
// (1, 13, 'sp4_r_v_b_33')
// (1, 14, 'sp4_r_v_b_20')
// (1, 14, 'sp4_r_v_b_4')
// (1, 15, 'sp4_r_v_b_9')
// (2, 10, 'sp4_v_t_41')
// (2, 11, 'neigh_op_top_6')
// (2, 11, 'sp4_r_v_b_40')
// (2, 11, 'sp4_v_b_41')
// (2, 11, 'sp4_v_t_44')
// (2, 12, 'local_g3_6')
// (2, 12, 'lutff_2/in_1')
// (2, 12, 'lutff_6/in_3')
// (2, 12, 'lutff_6/out')
// (2, 12, 'sp4_h_r_28')
// (2, 12, 'sp4_r_v_b_29')
// (2, 12, 'sp4_v_b_28')
// (2, 12, 'sp4_v_b_44')
// (2, 13, 'neigh_op_bot_6')
// (2, 13, 'sp4_r_v_b_16')
// (2, 13, 'sp4_v_b_17')
// (2, 13, 'sp4_v_b_33')
// (2, 14, 'local_g1_4')
// (2, 14, 'lutff_6/in_1')
// (2, 14, 'sp4_h_r_4')
// (2, 14, 'sp4_r_v_b_5')
// (2, 14, 'sp4_v_b_20')
// (2, 14, 'sp4_v_b_4')
// (2, 15, 'sp4_v_b_9')
// (3, 10, 'sp4_v_t_40')
// (3, 11, 'neigh_op_tnl_6')
// (3, 11, 'sp4_v_b_40')
// (3, 12, 'neigh_op_lft_6')
// (3, 12, 'sp4_h_r_41')
// (3, 12, 'sp4_v_b_29')
// (3, 13, 'neigh_op_bnl_6')
// (3, 13, 'sp4_v_b_16')
// (3, 14, 'local_g0_5')
// (3, 14, 'lutff_4/in_3')
// (3, 14, 'sp4_h_r_17')
// (3, 14, 'sp4_v_b_5')
// (4, 12, 'sp4_h_l_41')
// (4, 12, 'sp4_h_r_0')
// (4, 14, 'local_g2_4')
// (4, 14, 'lutff_1/in_1')
// (4, 14, 'sp4_h_r_28')
// (5, 12, 'local_g0_5')
// (5, 12, 'lutff_2/in_3')
// (5, 12, 'sp4_h_r_13')
// (5, 14, 'sp4_h_r_41')
// (6, 12, 'sp4_h_r_24')
// (6, 14, 'sp4_h_l_41')
// (7, 12, 'sp4_h_r_37')
// (8, 12, 'sp4_h_l_37')

wire n104;
// (0, 12, 'sp4_r_v_b_38')
// (0, 13, 'sp4_r_v_b_27')
// (0, 14, 'sp4_r_v_b_14')
// (0, 15, 'sp4_r_v_b_3')
// (1, 11, 'sp4_h_r_3')
// (1, 11, 'sp4_v_t_38')
// (1, 12, 'local_g3_6')
// (1, 12, 'lutff_5/in_2')
// (1, 12, 'sp4_v_b_38')
// (1, 13, 'sp4_v_b_27')
// (1, 14, 'sp4_v_b_14')
// (1, 15, 'sp4_v_b_3')
// (2, 11, 'sp4_h_r_14')
// (3, 10, 'neigh_op_tnr_3')
// (3, 11, 'neigh_op_rgt_3')
// (3, 11, 'sp4_h_r_27')
// (3, 12, 'neigh_op_bnr_3')
// (4, 10, 'neigh_op_top_3')
// (4, 11, 'lutff_3/out')
// (4, 11, 'sp4_h_r_38')
// (4, 12, 'neigh_op_bot_3')
// (5, 10, 'neigh_op_tnl_3')
// (5, 11, 'neigh_op_lft_3')
// (5, 11, 'sp4_h_l_38')
// (5, 12, 'neigh_op_bnl_3')

wire n105;
// (0, 13, 'neigh_op_tnr_0')
// (0, 14, 'neigh_op_rgt_0')
// (0, 15, 'neigh_op_bnr_0')
// (1, 2, 'sp12_v_t_23')
// (1, 3, 'sp12_v_b_23')
// (1, 4, 'sp12_v_b_20')
// (1, 5, 'sp12_v_b_19')
// (1, 6, 'sp12_v_b_16')
// (1, 7, 'sp12_v_b_15')
// (1, 8, 'sp12_v_b_12')
// (1, 9, 'sp12_v_b_11')
// (1, 10, 'sp12_v_b_8')
// (1, 11, 'sp12_v_b_7')
// (1, 12, 'sp12_v_b_4')
// (1, 13, 'local_g3_3')
// (1, 13, 'lutff_global/cen')
// (1, 13, 'neigh_op_top_0')
// (1, 13, 'sp12_v_b_3')
// (1, 14, 'lutff_0/out')
// (1, 14, 'sp12_v_b_0')
// (1, 15, 'neigh_op_bot_0')
// (2, 13, 'neigh_op_tnl_0')
// (2, 14, 'neigh_op_lft_0')
// (2, 15, 'neigh_op_bnl_0')

wire n106;
// (0, 13, 'neigh_op_tnr_1')
// (0, 14, 'neigh_op_rgt_1')
// (0, 14, 'sp4_h_r_23')
// (0, 15, 'neigh_op_bnr_1')
// (1, 8, 'sp4_r_v_b_43')
// (1, 9, 'sp4_r_v_b_30')
// (1, 10, 'sp4_r_v_b_19')
// (1, 11, 'sp4_r_v_b_6')
// (1, 12, 'sp4_r_v_b_43')
// (1, 13, 'local_g0_1')
// (1, 13, 'lutff_5/in_2')
// (1, 13, 'neigh_op_top_1')
// (1, 13, 'sp4_r_v_b_30')
// (1, 14, 'lutff_1/out')
// (1, 14, 'sp4_h_r_34')
// (1, 14, 'sp4_r_v_b_19')
// (1, 15, 'neigh_op_bot_1')
// (1, 15, 'sp4_r_v_b_6')
// (2, 7, 'sp4_r_v_b_42')
// (2, 7, 'sp4_v_t_43')
// (2, 8, 'sp4_r_v_b_31')
// (2, 8, 'sp4_v_b_43')
// (2, 9, 'local_g3_6')
// (2, 9, 'lutff_4/in_1')
// (2, 9, 'lutff_7/in_0')
// (2, 9, 'sp4_r_v_b_18')
// (2, 9, 'sp4_v_b_30')
// (2, 10, 'local_g0_3')
// (2, 10, 'lutff_0/in_3')
// (2, 10, 'lutff_2/in_3')
// (2, 10, 'sp4_r_v_b_7')
// (2, 10, 'sp4_v_b_19')
// (2, 11, 'sp4_r_v_b_41')
// (2, 11, 'sp4_v_b_6')
// (2, 11, 'sp4_v_t_43')
// (2, 12, 'sp4_r_v_b_28')
// (2, 12, 'sp4_v_b_43')
// (2, 13, 'neigh_op_tnl_1')
// (2, 13, 'sp4_r_v_b_17')
// (2, 13, 'sp4_v_b_30')
// (2, 14, 'neigh_op_lft_1')
// (2, 14, 'sp4_h_r_47')
// (2, 14, 'sp4_r_v_b_4')
// (2, 14, 'sp4_v_b_19')
// (2, 15, 'neigh_op_bnl_1')
// (2, 15, 'sp4_v_b_6')
// (3, 6, 'sp4_v_t_42')
// (3, 7, 'sp4_v_b_42')
// (3, 8, 'sp4_v_b_31')
// (3, 9, 'local_g0_2')
// (3, 9, 'lutff_7/in_1')
// (3, 9, 'sp4_v_b_18')
// (3, 10, 'sp4_v_b_7')
// (3, 10, 'sp4_v_t_41')
// (3, 11, 'sp4_v_b_41')
// (3, 12, 'sp4_v_b_28')
// (3, 13, 'sp4_v_b_17')
// (3, 14, 'local_g1_6')
// (3, 14, 'lutff_5/in_2')
// (3, 14, 'sp4_h_l_47')
// (3, 14, 'sp4_h_r_6')
// (3, 14, 'sp4_v_b_4')
// (4, 14, 'sp4_h_r_19')
// (5, 14, 'sp4_h_r_30')
// (6, 14, 'sp4_h_r_43')
// (7, 14, 'sp4_h_l_43')

reg n107 = 0;
// (0, 13, 'neigh_op_tnr_3')
// (0, 14, 'neigh_op_rgt_3')
// (0, 15, 'neigh_op_bnr_3')
// (1, 13, 'neigh_op_top_3')
// (1, 14, 'local_g2_3')
// (1, 14, 'lutff_0/in_3')
// (1, 14, 'lutff_3/in_0')
// (1, 14, 'lutff_3/out')
// (1, 15, 'neigh_op_bot_3')
// (2, 13, 'neigh_op_tnl_3')
// (2, 14, 'neigh_op_lft_3')
// (2, 15, 'neigh_op_bnl_3')

reg n108 = 0;
// (0, 13, 'neigh_op_tnr_4')
// (0, 14, 'neigh_op_rgt_4')
// (0, 15, 'neigh_op_bnr_4')
// (1, 13, 'neigh_op_top_4')
// (1, 14, 'local_g3_4')
// (1, 14, 'lutff_4/in_1')
// (1, 14, 'lutff_4/out')
// (1, 15, 'local_g0_4')
// (1, 15, 'lutff_2/in_2')
// (1, 15, 'neigh_op_bot_4')
// (2, 13, 'neigh_op_tnl_4')
// (2, 14, 'neigh_op_lft_4')
// (2, 15, 'neigh_op_bnl_4')

wire n109;
// (0, 13, 'neigh_op_tnr_5')
// (0, 14, 'neigh_op_rgt_5')
// (0, 15, 'neigh_op_bnr_5')
// (1, 13, 'neigh_op_top_5')
// (1, 14, 'local_g3_5')
// (1, 14, 'lutff_3/in_3')
// (1, 14, 'lutff_5/out')
// (1, 15, 'neigh_op_bot_5')
// (2, 13, 'neigh_op_tnl_5')
// (2, 14, 'neigh_op_lft_5')
// (2, 15, 'neigh_op_bnl_5')

reg n110 = 0;
// (0, 13, 'neigh_op_tnr_6')
// (0, 13, 'sp4_r_v_b_41')
// (0, 14, 'neigh_op_rgt_6')
// (0, 14, 'sp4_r_v_b_28')
// (0, 15, 'neigh_op_bnr_6')
// (0, 15, 'sp4_r_v_b_17')
// (0, 16, 'sp4_r_v_b_4')
// (1, 12, 'local_g0_4')
// (1, 12, 'lutff_0/in_2')
// (1, 12, 'sp4_h_r_4')
// (1, 12, 'sp4_v_t_41')
// (1, 13, 'local_g1_6')
// (1, 13, 'lutff_7/in_2')
// (1, 13, 'neigh_op_top_6')
// (1, 13, 'sp4_v_b_41')
// (1, 14, 'local_g3_6')
// (1, 14, 'lutff_5/in_2')
// (1, 14, 'lutff_6/in_3')
// (1, 14, 'lutff_6/out')
// (1, 14, 'sp4_v_b_28')
// (1, 15, 'neigh_op_bot_6')
// (1, 15, 'sp4_v_b_17')
// (1, 16, 'sp4_v_b_4')
// (2, 12, 'sp4_h_r_17')
// (2, 13, 'neigh_op_tnl_6')
// (2, 14, 'neigh_op_lft_6')
// (2, 15, 'neigh_op_bnl_6')
// (3, 12, 'sp4_h_r_28')
// (4, 12, 'sp4_h_r_41')
// (5, 12, 'sp4_h_l_41')

wire n111;
// (0, 13, 'neigh_op_tnr_7')
// (0, 14, 'neigh_op_rgt_7')
// (0, 14, 'sp4_h_r_3')
// (0, 14, 'sp4_r_v_b_46')
// (0, 15, 'neigh_op_bnr_7')
// (0, 15, 'sp4_r_v_b_35')
// (0, 16, 'sp4_r_v_b_22')
// (0, 17, 'sp4_r_v_b_11')
// (1, 13, 'neigh_op_top_7')
// (1, 13, 'sp4_r_v_b_42')
// (1, 13, 'sp4_v_t_46')
// (1, 14, 'lutff_7/out')
// (1, 14, 'sp4_h_r_14')
// (1, 14, 'sp4_r_v_b_31')
// (1, 14, 'sp4_v_b_46')
// (1, 15, 'neigh_op_bot_7')
// (1, 15, 'sp4_r_v_b_18')
// (1, 15, 'sp4_v_b_35')
// (1, 16, 'sp4_r_v_b_7')
// (1, 16, 'sp4_v_b_22')
// (1, 17, 'sp4_h_r_5')
// (1, 17, 'sp4_r_v_b_47')
// (1, 17, 'sp4_v_b_11')
// (1, 18, 'sp4_r_v_b_34')
// (1, 19, 'local_g3_7')
// (1, 19, 'lutff_3/in_1')
// (1, 19, 'sp4_r_v_b_23')
// (1, 20, 'sp4_r_v_b_10')
// (2, 12, 'sp4_v_t_42')
// (2, 13, 'neigh_op_tnl_7')
// (2, 13, 'sp4_v_b_42')
// (2, 14, 'neigh_op_lft_7')
// (2, 14, 'sp4_h_r_27')
// (2, 14, 'sp4_v_b_31')
// (2, 15, 'neigh_op_bnl_7')
// (2, 15, 'sp4_v_b_18')
// (2, 16, 'sp4_h_r_7')
// (2, 16, 'sp4_v_b_7')
// (2, 16, 'sp4_v_t_47')
// (2, 17, 'sp4_h_r_16')
// (2, 17, 'sp4_v_b_47')
// (2, 18, 'sp4_v_b_34')
// (2, 19, 'sp4_v_b_23')
// (2, 20, 'sp4_v_b_10')
// (3, 14, 'sp4_h_r_38')
// (3, 15, 'sp4_r_v_b_45')
// (3, 16, 'local_g1_2')
// (3, 16, 'lutff_7/in_0')
// (3, 16, 'sp4_h_r_18')
// (3, 16, 'sp4_r_v_b_32')
// (3, 17, 'sp4_h_r_29')
// (3, 17, 'sp4_r_v_b_21')
// (3, 18, 'sp4_r_v_b_8')
// (4, 14, 'sp4_h_l_38')
// (4, 14, 'sp4_v_t_45')
// (4, 15, 'sp4_v_b_45')
// (4, 16, 'sp4_h_r_31')
// (4, 16, 'sp4_v_b_32')
// (4, 17, 'local_g1_5')
// (4, 17, 'local_g3_0')
// (4, 17, 'lutff_0/in_3')
// (4, 17, 'lutff_5/in_3')
// (4, 17, 'lutff_7/in_1')
// (4, 17, 'sp4_h_r_40')
// (4, 17, 'sp4_v_b_21')
// (4, 18, 'sp4_v_b_8')
// (5, 16, 'sp4_h_r_42')
// (5, 17, 'sp4_h_l_40')
// (6, 16, 'sp4_h_l_42')

wire n112;
// (0, 13, 'sp4_h_r_11')
// (1, 13, 'sp4_h_r_22')
// (2, 12, 'local_g2_7')
// (2, 12, 'lutff_1/in_0')
// (2, 12, 'sp4_r_v_b_39')
// (2, 13, 'local_g2_3')
// (2, 13, 'lutff_2/in_3')
// (2, 13, 'sp4_h_r_35')
// (2, 13, 'sp4_r_v_b_26')
// (2, 14, 'sp4_r_v_b_15')
// (2, 15, 'sp4_r_v_b_2')
// (2, 16, 'local_g2_5')
// (2, 16, 'lutff_6/in_1')
// (2, 16, 'neigh_op_tnr_5')
// (2, 16, 'sp4_r_v_b_39')
// (2, 17, 'neigh_op_rgt_5')
// (2, 17, 'sp4_r_v_b_26')
// (2, 18, 'local_g0_5')
// (2, 18, 'lutff_0/in_3')
// (2, 18, 'lutff_1/in_2')
// (2, 18, 'lutff_3/in_2')
// (2, 18, 'lutff_5/in_0')
// (2, 18, 'neigh_op_bnr_5')
// (2, 18, 'sp4_r_v_b_15')
// (2, 19, 'sp4_r_v_b_2')
// (2, 20, 'sp4_r_v_b_39')
// (2, 21, 'local_g1_2')
// (2, 21, 'lutff_7/in_2')
// (2, 21, 'sp4_r_v_b_26')
// (2, 22, 'sp4_r_v_b_15')
// (2, 23, 'sp4_r_v_b_2')
// (3, 11, 'sp4_v_t_39')
// (3, 12, 'sp4_v_b_39')
// (3, 13, 'sp4_h_r_46')
// (3, 13, 'sp4_v_b_26')
// (3, 14, 'sp4_r_v_b_46')
// (3, 14, 'sp4_v_b_15')
// (3, 15, 'sp4_r_v_b_35')
// (3, 15, 'sp4_v_b_2')
// (3, 15, 'sp4_v_t_39')
// (3, 16, 'local_g1_5')
// (3, 16, 'lutff_4/in_0')
// (3, 16, 'neigh_op_top_5')
// (3, 16, 'sp4_r_v_b_22')
// (3, 16, 'sp4_v_b_39')
// (3, 17, 'lutff_5/out')
// (3, 17, 'sp4_r_v_b_11')
// (3, 17, 'sp4_v_b_26')
// (3, 18, 'local_g0_5')
// (3, 18, 'lutff_3/in_2')
// (3, 18, 'neigh_op_bot_5')
// (3, 18, 'sp4_v_b_15')
// (3, 19, 'sp4_v_b_2')
// (3, 19, 'sp4_v_t_39')
// (3, 20, 'sp4_v_b_39')
// (3, 21, 'sp4_v_b_26')
// (3, 22, 'sp4_v_b_15')
// (3, 23, 'sp4_v_b_2')
// (4, 13, 'sp4_h_l_46')
// (4, 13, 'sp4_v_t_46')
// (4, 14, 'sp4_v_b_46')
// (4, 15, 'sp4_v_b_35')
// (4, 16, 'neigh_op_tnl_5')
// (4, 16, 'sp4_v_b_22')
// (4, 17, 'neigh_op_lft_5')
// (4, 17, 'sp4_v_b_11')
// (4, 18, 'neigh_op_bnl_5')

reg n113 = 0;
// (0, 13, 'sp4_h_r_2')
// (1, 12, 'local_g2_5')
// (1, 12, 'lutff_6/in_3')
// (1, 12, 'neigh_op_tnr_5')
// (1, 13, 'neigh_op_rgt_5')
// (1, 13, 'sp4_h_r_15')
// (1, 14, 'neigh_op_bnr_5')
// (1, 14, 'sp4_r_v_b_41')
// (1, 15, 'sp4_r_v_b_28')
// (1, 16, 'sp4_r_v_b_17')
// (1, 17, 'local_g1_4')
// (1, 17, 'lutff_5/in_0')
// (1, 17, 'sp4_r_v_b_4')
// (2, 10, 'sp4_r_v_b_46')
// (2, 11, 'sp4_r_v_b_35')
// (2, 12, 'neigh_op_top_5')
// (2, 12, 'sp4_r_v_b_22')
// (2, 13, 'local_g3_5')
// (2, 13, 'lutff_5/in_1')
// (2, 13, 'lutff_5/out')
// (2, 13, 'sp4_h_r_10')
// (2, 13, 'sp4_h_r_26')
// (2, 13, 'sp4_r_v_b_11')
// (2, 13, 'sp4_v_t_41')
// (2, 14, 'local_g1_5')
// (2, 14, 'lutff_2/in_0')
// (2, 14, 'neigh_op_bot_5')
// (2, 14, 'sp4_v_b_41')
// (2, 15, 'sp4_v_b_28')
// (2, 16, 'sp4_v_b_17')
// (2, 17, 'sp4_v_b_4')
// (3, 9, 'sp4_v_t_46')
// (3, 10, 'sp4_r_v_b_45')
// (3, 10, 'sp4_v_b_46')
// (3, 11, 'local_g3_3')
// (3, 11, 'lutff_6/in_0')
// (3, 11, 'sp4_r_v_b_32')
// (3, 11, 'sp4_v_b_35')
// (3, 12, 'local_g3_5')
// (3, 12, 'lutff_0/in_0')
// (3, 12, 'neigh_op_tnl_5')
// (3, 12, 'sp4_r_v_b_21')
// (3, 12, 'sp4_v_b_22')
// (3, 13, 'neigh_op_lft_5')
// (3, 13, 'sp4_h_r_23')
// (3, 13, 'sp4_h_r_39')
// (3, 13, 'sp4_r_v_b_8')
// (3, 13, 'sp4_v_b_11')
// (3, 14, 'local_g3_5')
// (3, 14, 'lutff_7/in_1')
// (3, 14, 'neigh_op_bnl_5')
// (4, 9, 'sp4_v_t_45')
// (4, 10, 'sp4_v_b_45')
// (4, 11, 'sp4_v_b_32')
// (4, 12, 'local_g1_5')
// (4, 12, 'lutff_1/in_1')
// (4, 12, 'sp4_v_b_21')
// (4, 13, 'sp4_h_l_39')
// (4, 13, 'sp4_h_r_34')
// (4, 13, 'sp4_v_b_8')
// (5, 10, 'sp4_r_v_b_41')
// (5, 11, 'sp4_r_v_b_28')
// (5, 12, 'local_g3_1')
// (5, 12, 'lutff_5/in_3')
// (5, 12, 'sp4_r_v_b_17')
// (5, 13, 'local_g2_7')
// (5, 13, 'lutff_3/in_0')
// (5, 13, 'lutff_4/in_1')
// (5, 13, 'lutff_7/in_0')
// (5, 13, 'sp4_h_r_47')
// (5, 13, 'sp4_r_v_b_4')
// (6, 9, 'sp4_v_t_41')
// (6, 10, 'sp4_v_b_41')
// (6, 11, 'sp4_v_b_28')
// (6, 12, 'sp4_v_b_17')
// (6, 13, 'sp4_h_l_47')
// (6, 13, 'sp4_v_b_4')

reg n114 = 0;
// (0, 14, 'neigh_op_tnr_2')
// (0, 15, 'neigh_op_rgt_2')
// (0, 16, 'neigh_op_bnr_2')
// (1, 4, 'sp4_r_v_b_36')
// (1, 5, 'sp4_r_v_b_25')
// (1, 6, 'sp4_r_v_b_12')
// (1, 7, 'sp4_r_v_b_1')
// (1, 8, 'sp4_r_v_b_40')
// (1, 9, 'sp4_r_v_b_29')
// (1, 10, 'sp4_r_v_b_16')
// (1, 11, 'sp4_r_v_b_5')
// (1, 12, 'sp4_r_v_b_40')
// (1, 13, 'sp4_r_v_b_29')
// (1, 14, 'neigh_op_top_2')
// (1, 14, 'sp4_r_v_b_16')
// (1, 15, 'lutff_2/out')
// (1, 15, 'sp4_r_v_b_37')
// (1, 15, 'sp4_r_v_b_5')
// (1, 16, 'neigh_op_bot_2')
// (1, 16, 'sp4_r_v_b_24')
// (1, 17, 'sp4_r_v_b_13')
// (1, 18, 'sp4_r_v_b_0')
// (2, 3, 'sp4_v_t_36')
// (2, 4, 'sp4_v_b_36')
// (2, 5, 'sp4_v_b_25')
// (2, 6, 'sp4_v_b_12')
// (2, 7, 'local_g1_1')
// (2, 7, 'lutff_7/in_1')
// (2, 7, 'sp4_v_b_1')
// (2, 7, 'sp4_v_t_40')
// (2, 8, 'sp4_v_b_40')
// (2, 9, 'sp4_v_b_29')
// (2, 10, 'sp4_v_b_16')
// (2, 11, 'sp4_v_b_5')
// (2, 11, 'sp4_v_t_40')
// (2, 12, 'sp4_v_b_40')
// (2, 13, 'sp4_v_b_29')
// (2, 14, 'neigh_op_tnl_2')
// (2, 14, 'sp4_v_b_16')
// (2, 14, 'sp4_v_t_37')
// (2, 15, 'neigh_op_lft_2')
// (2, 15, 'sp4_v_b_37')
// (2, 15, 'sp4_v_b_5')
// (2, 16, 'neigh_op_bnl_2')
// (2, 16, 'sp4_v_b_24')
// (2, 17, 'local_g0_5')
// (2, 17, 'lutff_7/in_0')
// (2, 17, 'sp4_v_b_13')
// (2, 18, 'sp4_v_b_0')

wire n115;
// (0, 14, 'neigh_op_tnr_3')
// (0, 15, 'neigh_op_rgt_3')
// (0, 16, 'neigh_op_bnr_3')
// (1, 14, 'local_g1_3')
// (1, 14, 'lutff_4/in_0')
// (1, 14, 'neigh_op_top_3')
// (1, 15, 'local_g3_3')
// (1, 15, 'lutff_3/out')
// (1, 15, 'lutff_global/cen')
// (1, 16, 'neigh_op_bot_3')
// (2, 14, 'neigh_op_tnl_3')
// (2, 15, 'neigh_op_lft_3')
// (2, 16, 'neigh_op_bnl_3')

wire n116;
// (0, 14, 'sp4_h_r_19')
// (1, 14, 'local_g2_6')
// (1, 14, 'lutff_1/in_1')
// (1, 14, 'sp4_h_r_30')
// (2, 7, 'sp4_r_v_b_36')
// (2, 8, 'neigh_op_tnr_6')
// (2, 8, 'sp4_r_v_b_25')
// (2, 9, 'neigh_op_rgt_6')
// (2, 9, 'sp4_r_v_b_12')
// (2, 10, 'neigh_op_bnr_6')
// (2, 10, 'sp4_r_v_b_1')
// (2, 11, 'sp4_r_v_b_36')
// (2, 12, 'sp4_r_v_b_25')
// (2, 13, 'sp4_r_v_b_12')
// (2, 14, 'sp4_h_r_43')
// (2, 14, 'sp4_r_v_b_1')
// (3, 6, 'sp4_v_t_36')
// (3, 7, 'sp4_v_b_36')
// (3, 8, 'neigh_op_top_6')
// (3, 8, 'sp4_v_b_25')
// (3, 9, 'lutff_6/out')
// (3, 9, 'sp4_v_b_12')
// (3, 10, 'neigh_op_bot_6')
// (3, 10, 'sp4_v_b_1')
// (3, 10, 'sp4_v_t_36')
// (3, 11, 'sp4_v_b_36')
// (3, 12, 'sp4_v_b_25')
// (3, 13, 'sp4_v_b_12')
// (3, 14, 'sp4_h_l_43')
// (3, 14, 'sp4_v_b_1')
// (4, 8, 'neigh_op_tnl_6')
// (4, 9, 'neigh_op_lft_6')
// (4, 10, 'neigh_op_bnl_6')

wire n117;
// (0, 14, 'sp4_h_r_4')
// (1, 12, 'local_g2_4')
// (1, 12, 'lutff_0/in_0')
// (1, 12, 'sp4_r_v_b_36')
// (1, 13, 'neigh_op_tnr_6')
// (1, 13, 'sp4_r_v_b_25')
// (1, 14, 'neigh_op_rgt_6')
// (1, 14, 'sp4_h_r_17')
// (1, 14, 'sp4_r_v_b_12')
// (1, 15, 'neigh_op_bnr_6')
// (1, 15, 'sp4_r_v_b_1')
// (2, 11, 'local_g1_6')
// (2, 11, 'lutff_5/in_0')
// (2, 11, 'sp4_h_r_6')
// (2, 11, 'sp4_v_t_36')
// (2, 12, 'local_g2_4')
// (2, 12, 'lutff_4/in_0')
// (2, 12, 'lutff_6/in_2')
// (2, 12, 'sp4_v_b_36')
// (2, 13, 'local_g1_6')
// (2, 13, 'lutff_0/in_3')
// (2, 13, 'neigh_op_top_6')
// (2, 13, 'sp4_v_b_25')
// (2, 14, 'local_g3_6')
// (2, 14, 'lutff_5/in_2')
// (2, 14, 'lutff_6/out')
// (2, 14, 'sp4_h_r_28')
// (2, 14, 'sp4_v_b_12')
// (2, 15, 'local_g1_6')
// (2, 15, 'lutff_3/in_0')
// (2, 15, 'neigh_op_bot_6')
// (2, 15, 'sp4_v_b_1')
// (3, 11, 'sp4_h_r_19')
// (3, 13, 'neigh_op_tnl_6')
// (3, 14, 'neigh_op_lft_6')
// (3, 14, 'sp4_h_r_41')
// (3, 15, 'neigh_op_bnl_6')
// (3, 15, 'sp4_r_v_b_44')
// (3, 16, 'sp4_r_v_b_33')
// (3, 17, 'sp4_r_v_b_20')
// (3, 18, 'sp4_r_v_b_9')
// (4, 11, 'sp4_h_r_30')
// (4, 14, 'sp4_h_l_41')
// (4, 14, 'sp4_v_t_44')
// (4, 15, 'sp4_v_b_44')
// (4, 16, 'local_g2_1')
// (4, 16, 'lutff_0/in_1')
// (4, 16, 'lutff_7/in_0')
// (4, 16, 'sp4_v_b_33')
// (4, 17, 'sp4_v_b_20')
// (4, 18, 'sp4_v_b_9')
// (5, 11, 'sp4_h_r_43')
// (6, 11, 'sp4_h_l_43')

wire n118;
// (0, 14, 'sp4_r_v_b_38')
// (0, 15, 'sp4_r_v_b_27')
// (0, 16, 'sp4_r_v_b_14')
// (0, 17, 'neigh_op_tnr_5')
// (0, 17, 'sp4_r_v_b_3')
// (0, 18, 'neigh_op_rgt_5')
// (0, 18, 'sp4_r_v_b_42')
// (0, 19, 'neigh_op_bnr_5')
// (0, 19, 'sp4_r_v_b_31')
// (0, 20, 'sp4_r_v_b_18')
// (0, 21, 'sp4_r_v_b_7')
// (1, 13, 'sp4_v_t_38')
// (1, 14, 'sp4_v_b_38')
// (1, 15, 'sp4_v_b_27')
// (1, 16, 'sp4_v_b_14')
// (1, 17, 'local_g1_3')
// (1, 17, 'lutff_global/cen')
// (1, 17, 'neigh_op_top_5')
// (1, 17, 'sp4_v_b_3')
// (1, 17, 'sp4_v_t_42')
// (1, 18, 'lutff_5/out')
// (1, 18, 'sp4_v_b_42')
// (1, 19, 'neigh_op_bot_5')
// (1, 19, 'sp4_v_b_31')
// (1, 20, 'sp4_v_b_18')
// (1, 21, 'sp4_v_b_7')
// (2, 17, 'neigh_op_tnl_5')
// (2, 18, 'neigh_op_lft_5')
// (2, 19, 'neigh_op_bnl_5')

reg n119 = 0;
// (0, 15, 'neigh_op_tnr_1')
// (0, 16, 'neigh_op_rgt_1')
// (0, 17, 'neigh_op_bnr_1')
// (1, 15, 'neigh_op_top_1')
// (1, 16, 'local_g2_1')
// (1, 16, 'lutff_1/in_2')
// (1, 16, 'lutff_1/out')
// (1, 17, 'neigh_op_bot_1')
// (2, 15, 'neigh_op_tnl_1')
// (2, 16, 'local_g0_1')
// (2, 16, 'lutff_1/in_2')
// (2, 16, 'neigh_op_lft_1')
// (2, 17, 'neigh_op_bnl_1')

reg n120 = 0;
// (0, 15, 'neigh_op_tnr_2')
// (0, 16, 'neigh_op_rgt_2')
// (0, 17, 'neigh_op_bnr_2')
// (1, 15, 'neigh_op_top_2')
// (1, 16, 'local_g0_2')
// (1, 16, 'lutff_2/in_0')
// (1, 16, 'lutff_2/out')
// (1, 17, 'neigh_op_bot_2')
// (2, 15, 'neigh_op_tnl_2')
// (2, 16, 'local_g0_2')
// (2, 16, 'lutff_1/in_3')
// (2, 16, 'neigh_op_lft_2')
// (2, 17, 'neigh_op_bnl_2')

wire n121;
// (0, 15, 'sp4_h_r_6')
// (1, 14, 'neigh_op_tnr_7')
// (1, 15, 'neigh_op_rgt_7')
// (1, 15, 'sp4_h_r_19')
// (1, 16, 'neigh_op_bnr_7')
// (2, 14, 'neigh_op_top_7')
// (2, 15, 'lutff_7/out')
// (2, 15, 'sp4_h_r_30')
// (2, 16, 'neigh_op_bot_7')
// (3, 12, 'sp4_r_v_b_37')
// (3, 13, 'sp4_r_v_b_24')
// (3, 14, 'neigh_op_tnl_7')
// (3, 14, 'sp4_r_v_b_13')
// (3, 15, 'neigh_op_lft_7')
// (3, 15, 'sp4_h_r_43')
// (3, 15, 'sp4_r_v_b_0')
// (3, 16, 'neigh_op_bnl_7')
// (4, 11, 'sp4_v_t_37')
// (4, 12, 'sp4_v_b_37')
// (4, 13, 'local_g3_0')
// (4, 13, 'lutff_7/in_2')
// (4, 13, 'sp4_v_b_24')
// (4, 14, 'sp4_v_b_13')
// (4, 15, 'sp4_h_l_43')
// (4, 15, 'sp4_v_b_0')

reg n122 = 0;
// (0, 16, 'neigh_op_tnr_2')
// (0, 17, 'neigh_op_rgt_2')
// (0, 18, 'neigh_op_bnr_2')
// (1, 16, 'neigh_op_top_2')
// (1, 17, 'local_g0_2')
// (1, 17, 'lutff_2/in_2')
// (1, 17, 'lutff_2/out')
// (1, 17, 'lutff_6/in_0')
// (1, 18, 'neigh_op_bot_2')
// (2, 16, 'neigh_op_tnl_2')
// (2, 17, 'local_g0_2')
// (2, 17, 'lutff_6/in_2')
// (2, 17, 'neigh_op_lft_2')
// (2, 18, 'neigh_op_bnl_2')

reg n123 = 0;
// (0, 16, 'neigh_op_tnr_4')
// (0, 17, 'neigh_op_rgt_4')
// (0, 18, 'neigh_op_bnr_4')
// (1, 16, 'neigh_op_top_4')
// (1, 17, 'local_g3_4')
// (1, 17, 'lutff_1/in_2')
// (1, 17, 'lutff_4/in_3')
// (1, 17, 'lutff_4/out')
// (1, 17, 'lutff_6/in_3')
// (1, 18, 'neigh_op_bot_4')
// (2, 16, 'neigh_op_tnl_4')
// (2, 17, 'local_g0_4')
// (2, 17, 'lutff_6/in_0')
// (2, 17, 'neigh_op_lft_4')
// (2, 18, 'neigh_op_bnl_4')

wire n124;
// (0, 16, 'neigh_op_tnr_5')
// (0, 17, 'neigh_op_rgt_5')
// (0, 18, 'neigh_op_bnr_5')
// (1, 16, 'neigh_op_top_5')
// (1, 17, 'lutff_5/out')
// (1, 17, 'sp4_h_r_10')
// (1, 18, 'neigh_op_bot_5')
// (2, 16, 'neigh_op_tnl_5')
// (2, 17, 'local_g1_7')
// (2, 17, 'lutff_5/in_3')
// (2, 17, 'neigh_op_lft_5')
// (2, 17, 'sp4_h_r_23')
// (2, 18, 'neigh_op_bnl_5')
// (3, 17, 'sp4_h_r_34')
// (4, 17, 'sp4_h_r_47')
// (5, 17, 'sp4_h_l_47')

wire n125;
// (0, 16, 'neigh_op_tnr_6')
// (0, 17, 'neigh_op_rgt_6')
// (0, 17, 'sp4_h_r_17')
// (0, 18, 'neigh_op_bnr_6')
// (1, 16, 'neigh_op_top_6')
// (1, 17, 'lutff_6/out')
// (1, 17, 'sp4_h_r_28')
// (1, 18, 'neigh_op_bot_6')
// (2, 10, 'sp4_r_v_b_43')
// (2, 11, 'sp4_r_v_b_30')
// (2, 12, 'sp4_r_v_b_19')
// (2, 13, 'sp4_r_v_b_6')
// (2, 14, 'sp4_r_v_b_47')
// (2, 15, 'sp4_r_v_b_34')
// (2, 16, 'neigh_op_tnl_6')
// (2, 16, 'sp4_r_v_b_23')
// (2, 17, 'neigh_op_lft_6')
// (2, 17, 'sp4_h_r_41')
// (2, 17, 'sp4_r_v_b_10')
// (2, 18, 'neigh_op_bnl_6')
// (3, 9, 'sp4_v_t_43')
// (3, 10, 'sp4_v_b_43')
// (3, 11, 'sp4_v_b_30')
// (3, 12, 'local_g0_3')
// (3, 12, 'lutff_5/in_2')
// (3, 12, 'sp4_v_b_19')
// (3, 13, 'sp4_v_b_6')
// (3, 13, 'sp4_v_t_47')
// (3, 14, 'sp4_v_b_47')
// (3, 15, 'sp4_v_b_34')
// (3, 16, 'sp4_v_b_23')
// (3, 17, 'sp4_h_l_41')
// (3, 17, 'sp4_v_b_10')

reg n126 = 0;
// (0, 16, 'neigh_op_tnr_7')
// (0, 17, 'neigh_op_rgt_7')
// (0, 18, 'neigh_op_bnr_7')
// (1, 16, 'neigh_op_top_7')
// (1, 17, 'local_g2_7')
// (1, 17, 'lutff_0/in_1')
// (1, 17, 'lutff_4/in_1')
// (1, 17, 'lutff_7/in_0')
// (1, 17, 'lutff_7/out')
// (1, 18, 'neigh_op_bot_7')
// (2, 16, 'neigh_op_tnl_7')
// (2, 17, 'local_g0_7')
// (2, 17, 'lutff_6/in_3')
// (2, 17, 'neigh_op_lft_7')
// (2, 18, 'neigh_op_bnl_7')

wire n127;
// (0, 16, 'sp4_h_r_2')
// (1, 13, 'sp4_r_v_b_47')
// (1, 14, 'sp4_r_v_b_34')
// (1, 15, 'neigh_op_tnr_5')
// (1, 15, 'sp4_r_v_b_23')
// (1, 16, 'local_g2_2')
// (1, 16, 'lutff_global/cen')
// (1, 16, 'neigh_op_rgt_5')
// (1, 16, 'sp4_h_r_15')
// (1, 16, 'sp4_r_v_b_10')
// (1, 17, 'neigh_op_bnr_5')
// (2, 12, 'sp4_v_t_47')
// (2, 13, 'sp4_v_b_47')
// (2, 14, 'sp4_v_b_34')
// (2, 15, 'neigh_op_top_5')
// (2, 15, 'sp4_v_b_23')
// (2, 16, 'local_g2_2')
// (2, 16, 'lutff_5/out')
// (2, 16, 'lutff_global/cen')
// (2, 16, 'sp4_h_r_26')
// (2, 16, 'sp4_v_b_10')
// (2, 17, 'neigh_op_bot_5')
// (3, 15, 'neigh_op_tnl_5')
// (3, 16, 'neigh_op_lft_5')
// (3, 16, 'sp4_h_r_39')
// (3, 17, 'neigh_op_bnl_5')
// (4, 16, 'sp4_h_l_39')

wire n128;
// (0, 16, 'sp4_h_r_3')
// (1, 16, 'sp4_h_r_14')
// (2, 9, 'sp4_r_v_b_44')
// (2, 10, 'local_g0_2')
// (2, 10, 'lutff_1/in_1')
// (2, 10, 'sp4_r_v_b_33')
// (2, 11, 'local_g3_4')
// (2, 11, 'lutff_7/in_2')
// (2, 11, 'sp4_r_v_b_20')
// (2, 12, 'sp4_r_v_b_46')
// (2, 12, 'sp4_r_v_b_9')
// (2, 13, 'sp4_r_v_b_35')
// (2, 13, 'sp4_r_v_b_43')
// (2, 14, 'local_g1_6')
// (2, 14, 'lutff_4/in_3')
// (2, 14, 'lutff_5/in_0')
// (2, 14, 'sp4_r_v_b_22')
// (2, 14, 'sp4_r_v_b_30')
// (2, 15, 'neigh_op_tnr_3')
// (2, 15, 'sp4_r_v_b_11')
// (2, 15, 'sp4_r_v_b_19')
// (2, 16, 'neigh_op_rgt_3')
// (2, 16, 'sp4_h_r_11')
// (2, 16, 'sp4_h_r_27')
// (2, 16, 'sp4_r_v_b_38')
// (2, 16, 'sp4_r_v_b_6')
// (2, 17, 'neigh_op_bnr_3')
// (2, 17, 'sp4_r_v_b_27')
// (2, 18, 'sp4_r_v_b_14')
// (2, 19, 'sp4_r_v_b_3')
// (3, 8, 'sp4_v_t_44')
// (3, 9, 'sp4_r_v_b_40')
// (3, 9, 'sp4_v_b_44')
// (3, 10, 'sp4_r_v_b_29')
// (3, 10, 'sp4_v_b_33')
// (3, 11, 'local_g0_4')
// (3, 11, 'lutff_0/in_0')
// (3, 11, 'lutff_3/in_3')
// (3, 11, 'sp4_h_r_11')
// (3, 11, 'sp4_r_v_b_16')
// (3, 11, 'sp4_v_b_20')
// (3, 11, 'sp4_v_t_46')
// (3, 12, 'local_g1_1')
// (3, 12, 'lutff_2/in_2')
// (3, 12, 'sp4_h_r_11')
// (3, 12, 'sp4_r_v_b_5')
// (3, 12, 'sp4_v_b_46')
// (3, 12, 'sp4_v_b_9')
// (3, 12, 'sp4_v_t_43')
// (3, 13, 'sp4_r_v_b_44')
// (3, 13, 'sp4_v_b_35')
// (3, 13, 'sp4_v_b_43')
// (3, 14, 'sp4_r_v_b_33')
// (3, 14, 'sp4_r_v_b_47')
// (3, 14, 'sp4_v_b_22')
// (3, 14, 'sp4_v_b_30')
// (3, 15, 'neigh_op_top_3')
// (3, 15, 'sp4_r_v_b_20')
// (3, 15, 'sp4_r_v_b_34')
// (3, 15, 'sp4_v_b_11')
// (3, 15, 'sp4_v_b_19')
// (3, 15, 'sp4_v_t_38')
// (3, 16, 'local_g0_3')
// (3, 16, 'lutff_3/out')
// (3, 16, 'lutff_4/in_1')
// (3, 16, 'sp4_h_r_22')
// (3, 16, 'sp4_h_r_38')
// (3, 16, 'sp4_r_v_b_23')
// (3, 16, 'sp4_r_v_b_9')
// (3, 16, 'sp4_v_b_38')
// (3, 16, 'sp4_v_b_6')
// (3, 17, 'neigh_op_bot_3')
// (3, 17, 'sp4_r_v_b_10')
// (3, 17, 'sp4_v_b_27')
// (3, 18, 'sp4_v_b_14')
// (3, 19, 'sp4_v_b_3')
// (4, 8, 'sp4_v_t_40')
// (4, 9, 'sp4_v_b_40')
// (4, 10, 'sp4_v_b_29')
// (4, 11, 'local_g1_0')
// (4, 11, 'lutff_3/in_2')
// (4, 11, 'sp4_h_r_22')
// (4, 11, 'sp4_v_b_16')
// (4, 12, 'sp4_h_r_22')
// (4, 12, 'sp4_v_b_5')
// (4, 12, 'sp4_v_t_44')
// (4, 13, 'sp4_v_b_44')
// (4, 13, 'sp4_v_t_47')
// (4, 14, 'local_g2_7')
// (4, 14, 'lutff_0/in_3')
// (4, 14, 'lutff_6/in_1')
// (4, 14, 'sp4_v_b_33')
// (4, 14, 'sp4_v_b_47')
// (4, 15, 'neigh_op_tnl_3')
// (4, 15, 'sp4_v_b_20')
// (4, 15, 'sp4_v_b_34')
// (4, 16, 'local_g0_3')
// (4, 16, 'lutff_3/in_2')
// (4, 16, 'neigh_op_lft_3')
// (4, 16, 'sp4_h_l_38')
// (4, 16, 'sp4_h_r_35')
// (4, 16, 'sp4_v_b_23')
// (4, 16, 'sp4_v_b_9')
// (4, 17, 'neigh_op_bnl_3')
// (4, 17, 'sp4_v_b_10')
// (5, 11, 'local_g3_3')
// (5, 11, 'lutff_global/cen')
// (5, 11, 'sp4_h_r_35')
// (5, 12, 'local_g2_3')
// (5, 12, 'lutff_1/in_0')
// (5, 12, 'lutff_6/in_3')
// (5, 12, 'sp4_h_r_35')
// (5, 13, 'local_g3_0')
// (5, 13, 'lutff_0/in_3')
// (5, 13, 'lutff_7/in_2')
// (5, 13, 'sp4_r_v_b_40')
// (5, 14, 'local_g0_5')
// (5, 14, 'lutff_3/in_0')
// (5, 14, 'lutff_4/in_3')
// (5, 14, 'lutff_5/in_0')
// (5, 14, 'lutff_6/in_3')
// (5, 14, 'sp4_r_v_b_29')
// (5, 15, 'sp4_r_v_b_16')
// (5, 16, 'sp4_h_r_46')
// (5, 16, 'sp4_r_v_b_5')
// (6, 11, 'sp4_h_r_46')
// (6, 12, 'sp4_h_r_46')
// (6, 12, 'sp4_v_t_40')
// (6, 13, 'sp4_v_b_40')
// (6, 14, 'sp4_v_b_29')
// (6, 15, 'sp4_v_b_16')
// (6, 16, 'sp4_h_l_46')
// (6, 16, 'sp4_v_b_5')
// (7, 11, 'sp4_h_l_46')
// (7, 12, 'sp4_h_l_46')

wire n129;
// (0, 16, 'sp4_h_r_4')
// (1, 15, 'neigh_op_tnr_6')
// (1, 16, 'local_g3_6')
// (1, 16, 'lutff_1/in_0')
// (1, 16, 'lutff_2/in_1')
// (1, 16, 'neigh_op_rgt_6')
// (1, 16, 'sp4_h_r_17')
// (1, 17, 'neigh_op_bnr_6')
// (2, 15, 'neigh_op_top_6')
// (2, 16, 'local_g3_6')
// (2, 16, 'lutff_3/in_0')
// (2, 16, 'lutff_5/in_2')
// (2, 16, 'lutff_6/out')
// (2, 16, 'sp4_h_r_28')
// (2, 17, 'neigh_op_bot_6')
// (3, 15, 'neigh_op_tnl_6')
// (3, 16, 'neigh_op_lft_6')
// (3, 16, 'sp4_h_r_41')
// (3, 17, 'neigh_op_bnl_6')
// (4, 16, 'local_g1_0')
// (4, 16, 'lutff_6/in_3')
// (4, 16, 'sp4_h_l_41')
// (4, 16, 'sp4_h_r_0')
// (5, 16, 'sp4_h_r_13')
// (6, 16, 'sp4_h_r_24')
// (7, 16, 'sp4_h_r_37')
// (8, 16, 'sp4_h_l_37')

wire n130;
// (0, 17, 'neigh_op_tnr_0')
// (0, 18, 'neigh_op_rgt_0')
// (0, 19, 'neigh_op_bnr_0')
// (1, 17, 'neigh_op_top_0')
// (1, 18, 'local_g3_0')
// (1, 18, 'lutff_0/out')
// (1, 18, 'lutff_5/in_2')
// (1, 18, 'sp4_h_r_0')
// (1, 19, 'neigh_op_bot_0')
// (2, 17, 'neigh_op_tnl_0')
// (2, 18, 'neigh_op_lft_0')
// (2, 18, 'sp4_h_r_13')
// (2, 19, 'neigh_op_bnl_0')
// (3, 18, 'local_g3_0')
// (3, 18, 'lutff_7/in_2')
// (3, 18, 'sp4_h_r_24')
// (4, 18, 'sp4_h_r_37')
// (5, 18, 'sp4_h_l_37')

wire n131;
// (0, 17, 'sp12_h_r_5')
// (1, 17, 'sp12_h_r_6')
// (2, 16, 'neigh_op_tnr_1')
// (2, 17, 'neigh_op_rgt_1')
// (2, 17, 'sp12_h_r_9')
// (2, 18, 'neigh_op_bnr_1')
// (3, 16, 'neigh_op_top_1')
// (3, 17, 'lutff_1/out')
// (3, 17, 'sp12_h_r_10')
// (3, 18, 'neigh_op_bot_1')
// (4, 16, 'neigh_op_tnl_1')
// (4, 17, 'neigh_op_lft_1')
// (4, 17, 'sp12_h_r_13')
// (4, 18, 'neigh_op_bnl_1')
// (5, 17, 'sp12_h_r_14')
// (6, 17, 'sp12_h_r_17')
// (7, 17, 'local_g1_2')
// (7, 17, 'lutff_2/in_1')
// (7, 17, 'sp12_h_r_18')
// (8, 17, 'sp12_h_r_21')
// (9, 17, 'sp12_h_r_22')
// (10, 17, 'sp12_h_l_22')

reg n132 = 0;
// (0, 17, 'sp4_h_r_0')
// (1, 16, 'neigh_op_tnr_4')
// (1, 17, 'local_g2_4')
// (1, 17, 'lutff_6/in_2')
// (1, 17, 'neigh_op_rgt_4')
// (1, 17, 'sp4_h_r_13')
// (1, 18, 'local_g1_4')
// (1, 18, 'lutff_0/in_1')
// (1, 18, 'neigh_op_bnr_4')
// (2, 10, 'sp4_r_v_b_40')
// (2, 11, 'local_g0_5')
// (2, 11, 'lutff_4/in_1')
// (2, 11, 'sp4_r_v_b_29')
// (2, 12, 'sp4_r_v_b_16')
// (2, 13, 'sp4_r_v_b_5')
// (2, 14, 'sp4_r_v_b_44')
// (2, 15, 'sp4_r_v_b_33')
// (2, 16, 'neigh_op_top_4')
// (2, 16, 'sp4_r_v_b_20')
// (2, 16, 'sp4_r_v_b_36')
// (2, 17, 'local_g2_0')
// (2, 17, 'lutff_4/in_2')
// (2, 17, 'lutff_4/out')
// (2, 17, 'sp4_h_r_24')
// (2, 17, 'sp4_r_v_b_25')
// (2, 17, 'sp4_r_v_b_9')
// (2, 18, 'local_g1_4')
// (2, 18, 'lutff_7/in_2')
// (2, 18, 'neigh_op_bot_4')
// (2, 18, 'sp4_r_v_b_12')
// (2, 19, 'sp4_r_v_b_1')
// (3, 9, 'sp4_v_t_40')
// (3, 10, 'sp4_v_b_40')
// (3, 11, 'sp4_v_b_29')
// (3, 12, 'local_g0_0')
// (3, 12, 'lutff_6/in_2')
// (3, 12, 'sp4_v_b_16')
// (3, 13, 'sp4_v_b_5')
// (3, 13, 'sp4_v_t_44')
// (3, 14, 'sp4_r_v_b_37')
// (3, 14, 'sp4_v_b_44')
// (3, 15, 'local_g3_1')
// (3, 15, 'lutff_3/in_1')
// (3, 15, 'sp4_h_r_1')
// (3, 15, 'sp4_r_v_b_24')
// (3, 15, 'sp4_v_b_33')
// (3, 15, 'sp4_v_t_36')
// (3, 16, 'neigh_op_tnl_4')
// (3, 16, 'sp4_r_v_b_13')
// (3, 16, 'sp4_v_b_20')
// (3, 16, 'sp4_v_b_36')
// (3, 17, 'neigh_op_lft_4')
// (3, 17, 'sp4_h_r_37')
// (3, 17, 'sp4_r_v_b_0')
// (3, 17, 'sp4_v_b_25')
// (3, 17, 'sp4_v_b_9')
// (3, 18, 'local_g2_4')
// (3, 18, 'lutff_4/in_0')
// (3, 18, 'neigh_op_bnl_4')
// (3, 18, 'sp4_v_b_12')
// (3, 19, 'sp4_v_b_1')
// (4, 13, 'sp4_v_t_37')
// (4, 14, 'local_g2_5')
// (4, 14, 'lutff_3/in_2')
// (4, 14, 'sp4_v_b_37')
// (4, 15, 'local_g0_4')
// (4, 15, 'lutff_2/in_0')
// (4, 15, 'lutff_6/in_0')
// (4, 15, 'sp4_h_r_12')
// (4, 15, 'sp4_v_b_24')
// (4, 16, 'sp4_v_b_13')
// (4, 17, 'sp4_h_l_37')
// (4, 17, 'sp4_v_b_0')
// (5, 15, 'sp4_h_r_25')
// (6, 15, 'sp4_h_r_36')
// (7, 15, 'sp4_h_l_36')

wire n133;
// (0, 17, 'sp4_h_r_1')
// (1, 17, 'sp4_h_r_12')
// (2, 16, 'neigh_op_tnr_2')
// (2, 17, 'neigh_op_rgt_2')
// (2, 17, 'sp4_h_r_25')
// (2, 18, 'neigh_op_bnr_2')
// (3, 16, 'neigh_op_top_2')
// (3, 17, 'lutff_2/out')
// (3, 17, 'sp4_h_r_36')
// (3, 18, 'neigh_op_bot_2')
// (4, 16, 'neigh_op_tnl_2')
// (4, 17, 'neigh_op_lft_2')
// (4, 17, 'sp4_h_l_36')
// (4, 17, 'sp4_h_r_4')
// (4, 18, 'neigh_op_bnl_2')
// (5, 17, 'sp4_h_r_17')
// (6, 17, 'sp4_h_r_28')
// (7, 17, 'local_g2_1')
// (7, 17, 'lutff_4/in_3')
// (7, 17, 'sp4_h_r_41')
// (8, 17, 'sp4_h_l_41')

wire n134;
// (0, 17, 'sp4_h_r_30')
// (1, 15, 'sp4_h_r_3')
// (1, 17, 'local_g3_3')
// (1, 17, 'lutff_5/in_3')
// (1, 17, 'sp4_h_r_43')
// (1, 18, 'neigh_op_tnr_7')
// (1, 18, 'sp4_r_v_b_43')
// (1, 19, 'neigh_op_rgt_7')
// (1, 19, 'sp4_h_r_3')
// (1, 19, 'sp4_r_v_b_30')
// (1, 20, 'neigh_op_bnr_7')
// (1, 20, 'sp4_r_v_b_19')
// (1, 21, 'sp4_r_v_b_6')
// (2, 15, 'sp4_h_r_14')
// (2, 17, 'sp4_h_l_43')
// (2, 17, 'sp4_v_t_43')
// (2, 18, 'neigh_op_top_7')
// (2, 18, 'sp4_v_b_43')
// (2, 19, 'lutff_7/out')
// (2, 19, 'sp4_h_r_14')
// (2, 19, 'sp4_v_b_30')
// (2, 20, 'local_g0_7')
// (2, 20, 'lutff_4/in_3')
// (2, 20, 'neigh_op_bot_7')
// (2, 20, 'sp4_v_b_19')
// (2, 21, 'sp4_v_b_6')
// (3, 15, 'sp4_h_r_27')
// (3, 18, 'neigh_op_tnl_7')
// (3, 19, 'neigh_op_lft_7')
// (3, 19, 'sp4_h_r_27')
// (3, 20, 'neigh_op_bnl_7')
// (4, 15, 'local_g3_6')
// (4, 15, 'lutff_2/in_1')
// (4, 15, 'sp4_h_r_38')
// (4, 16, 'sp4_r_v_b_44')
// (4, 17, 'sp4_r_v_b_33')
// (4, 18, 'sp4_r_v_b_20')
// (4, 19, 'sp4_h_r_38')
// (4, 19, 'sp4_r_v_b_9')
// (5, 15, 'sp4_h_l_38')
// (5, 15, 'sp4_v_t_44')
// (5, 16, 'sp4_v_b_44')
// (5, 17, 'sp4_v_b_33')
// (5, 18, 'sp4_v_b_20')
// (5, 19, 'sp4_h_l_38')
// (5, 19, 'sp4_v_b_9')

reg n135 = 0;
// (0, 18, 'neigh_op_tnr_1')
// (0, 19, 'neigh_op_rgt_1')
// (0, 20, 'neigh_op_bnr_1')
// (1, 18, 'neigh_op_top_1')
// (1, 19, 'local_g3_1')
// (1, 19, 'lutff_1/in_1')
// (1, 19, 'lutff_1/out')
// (1, 19, 'lutff_4/in_2')
// (1, 19, 'lutff_5/in_3')
// (1, 20, 'neigh_op_bot_1')
// (2, 18, 'neigh_op_tnl_1')
// (2, 19, 'neigh_op_lft_1')
// (2, 20, 'neigh_op_bnl_1')

reg n136 = 0;
// (0, 18, 'neigh_op_tnr_2')
// (0, 19, 'neigh_op_rgt_2')
// (0, 20, 'neigh_op_bnr_2')
// (1, 18, 'neigh_op_top_2')
// (1, 19, 'local_g0_2')
// (1, 19, 'lutff_2/in_2')
// (1, 19, 'lutff_2/out')
// (1, 19, 'lutff_4/in_0')
// (1, 19, 'lutff_5/in_1')
// (1, 20, 'neigh_op_bot_2')
// (2, 18, 'neigh_op_tnl_2')
// (2, 19, 'neigh_op_lft_2')
// (2, 20, 'neigh_op_bnl_2')

wire n137;
// (0, 18, 'neigh_op_tnr_3')
// (0, 19, 'neigh_op_rgt_3')
// (0, 20, 'neigh_op_bnr_3')
// (1, 18, 'neigh_op_top_3')
// (1, 19, 'lutff_3/out')
// (1, 20, 'local_g1_3')
// (1, 20, 'lutff_4/in_0')
// (1, 20, 'lutff_6/in_2')
// (1, 20, 'lutff_7/in_1')
// (1, 20, 'neigh_op_bot_3')
// (2, 18, 'neigh_op_tnl_3')
// (2, 19, 'neigh_op_lft_3')
// (2, 20, 'neigh_op_bnl_3')

wire n138;
// (0, 18, 'neigh_op_tnr_4')
// (0, 19, 'neigh_op_rgt_4')
// (0, 19, 'sp4_h_r_13')
// (0, 20, 'neigh_op_bnr_4')
// (1, 18, 'neigh_op_top_4')
// (1, 19, 'lutff_4/out')
// (1, 19, 'sp4_h_r_24')
// (1, 20, 'neigh_op_bot_4')
// (2, 12, 'sp4_r_v_b_37')
// (2, 13, 'sp4_r_v_b_24')
// (2, 14, 'sp4_r_v_b_13')
// (2, 15, 'sp4_r_v_b_0')
// (2, 16, 'sp4_r_v_b_37')
// (2, 17, 'sp4_r_v_b_24')
// (2, 18, 'neigh_op_tnl_4')
// (2, 18, 'sp4_r_v_b_13')
// (2, 19, 'neigh_op_lft_4')
// (2, 19, 'sp4_h_r_37')
// (2, 19, 'sp4_r_v_b_0')
// (2, 20, 'neigh_op_bnl_4')
// (3, 11, 'sp4_v_t_37')
// (3, 12, 'local_g2_5')
// (3, 12, 'lutff_4/in_1')
// (3, 12, 'sp4_v_b_37')
// (3, 13, 'sp4_v_b_24')
// (3, 14, 'sp4_v_b_13')
// (3, 15, 'sp4_v_b_0')
// (3, 15, 'sp4_v_t_37')
// (3, 16, 'sp4_v_b_37')
// (3, 17, 'sp4_v_b_24')
// (3, 18, 'sp4_v_b_13')
// (3, 19, 'sp4_h_l_37')
// (3, 19, 'sp4_v_b_0')

wire n139;
// (0, 18, 'neigh_op_tnr_5')
// (0, 19, 'neigh_op_rgt_5')
// (0, 20, 'neigh_op_bnr_5')
// (1, 18, 'neigh_op_top_5')
// (1, 19, 'local_g2_5')
// (1, 19, 'lutff_5/out')
// (1, 19, 'lutff_6/in_1')
// (1, 19, 'sp4_h_r_10')
// (1, 20, 'neigh_op_bot_5')
// (2, 18, 'local_g2_5')
// (2, 18, 'local_g3_5')
// (2, 18, 'lutff_2/in_1')
// (2, 18, 'lutff_4/in_2')
// (2, 18, 'lutff_6/in_2')
// (2, 18, 'neigh_op_tnl_5')
// (2, 19, 'local_g0_7')
// (2, 19, 'lutff_4/in_1')
// (2, 19, 'neigh_op_lft_5')
// (2, 19, 'sp4_h_r_23')
// (2, 20, 'neigh_op_bnl_5')
// (3, 19, 'local_g3_2')
// (3, 19, 'lutff_7/in_2')
// (3, 19, 'sp4_h_r_34')
// (4, 16, 'sp4_r_v_b_41')
// (4, 17, 'sp4_r_v_b_28')
// (4, 18, 'sp4_r_v_b_17')
// (4, 19, 'sp4_h_r_47')
// (4, 19, 'sp4_r_v_b_4')
// (5, 15, 'sp4_v_t_41')
// (5, 16, 'sp4_v_b_41')
// (5, 17, 'local_g3_4')
// (5, 17, 'lutff_5/in_2')
// (5, 17, 'sp4_v_b_28')
// (5, 18, 'sp4_v_b_17')
// (5, 19, 'sp4_h_l_47')
// (5, 19, 'sp4_v_b_4')

wire n140;
// (0, 18, 'neigh_op_tnr_6')
// (0, 19, 'neigh_op_rgt_6')
// (0, 19, 'sp4_h_r_33')
// (0, 20, 'neigh_op_bnr_6')
// (1, 16, 'sp4_r_v_b_38')
// (1, 17, 'sp4_r_v_b_27')
// (1, 18, 'neigh_op_top_6')
// (1, 18, 'sp4_r_v_b_14')
// (1, 19, 'local_g1_3')
// (1, 19, 'lutff_6/out')
// (1, 19, 'lutff_global/cen')
// (1, 19, 'sp4_h_r_44')
// (1, 19, 'sp4_r_v_b_3')
// (1, 20, 'neigh_op_bot_6')
// (2, 15, 'sp4_v_t_38')
// (2, 16, 'sp4_v_b_38')
// (2, 17, 'sp4_v_b_27')
// (2, 18, 'neigh_op_tnl_6')
// (2, 18, 'sp4_v_b_14')
// (2, 19, 'neigh_op_lft_6')
// (2, 19, 'sp4_h_l_44')
// (2, 19, 'sp4_v_b_3')
// (2, 20, 'neigh_op_bnl_6')

reg n141 = 0;
// (0, 18, 'neigh_op_tnr_7')
// (0, 19, 'neigh_op_rgt_7')
// (0, 20, 'neigh_op_bnr_7')
// (1, 18, 'neigh_op_top_7')
// (1, 19, 'local_g1_7')
// (1, 19, 'local_g2_7')
// (1, 19, 'lutff_0/in_1')
// (1, 19, 'lutff_1/in_3')
// (1, 19, 'lutff_5/in_0')
// (1, 19, 'lutff_7/in_0')
// (1, 19, 'lutff_7/out')
// (1, 20, 'neigh_op_bot_7')
// (2, 18, 'neigh_op_tnl_7')
// (2, 19, 'neigh_op_lft_7')
// (2, 20, 'neigh_op_bnl_7')

reg n142 = 0;
// (0, 18, 'sp4_r_v_b_37')
// (0, 19, 'sp4_r_v_b_24')
// (0, 20, 'sp4_r_v_b_13')
// (0, 21, 'sp4_r_v_b_0')
// (1, 17, 'sp4_h_r_6')
// (1, 17, 'sp4_v_t_37')
// (1, 18, 'sp4_v_b_37')
// (1, 19, 'local_g2_0')
// (1, 19, 'lutff_3/in_3')
// (1, 19, 'lutff_6/in_2')
// (1, 19, 'sp4_v_b_24')
// (1, 20, 'sp4_v_b_13')
// (1, 21, 'sp4_v_b_0')
// (2, 7, 'sp4_r_v_b_43')
// (2, 8, 'sp4_r_v_b_30')
// (2, 9, 'sp4_r_v_b_19')
// (2, 10, 'local_g1_6')
// (2, 10, 'lutff_7/in_0')
// (2, 10, 'sp4_r_v_b_6')
// (2, 11, 'local_g3_3')
// (2, 11, 'lutff_4/in_0')
// (2, 11, 'sp4_r_v_b_38')
// (2, 11, 'sp4_r_v_b_43')
// (2, 12, 'local_g0_3')
// (2, 12, 'lutff_4/in_1')
// (2, 12, 'sp4_r_v_b_27')
// (2, 12, 'sp4_r_v_b_30')
// (2, 13, 'sp4_r_v_b_14')
// (2, 13, 'sp4_r_v_b_19')
// (2, 14, 'sp4_r_v_b_3')
// (2, 14, 'sp4_r_v_b_6')
// (2, 15, 'local_g2_6')
// (2, 15, 'lutff_0/in_0')
// (2, 15, 'sp4_r_v_b_38')
// (2, 16, 'neigh_op_tnr_7')
// (2, 16, 'sp4_r_v_b_27')
// (2, 17, 'neigh_op_rgt_7')
// (2, 17, 'sp4_h_r_19')
// (2, 17, 'sp4_r_v_b_14')
// (2, 17, 'sp4_r_v_b_46')
// (2, 18, 'local_g1_7')
// (2, 18, 'lutff_4/in_0')
// (2, 18, 'lutff_6/in_0')
// (2, 18, 'lutff_7/in_1')
// (2, 18, 'neigh_op_bnr_7')
// (2, 18, 'sp4_r_v_b_3')
// (2, 18, 'sp4_r_v_b_35')
// (2, 19, 'sp4_r_v_b_22')
// (2, 20, 'local_g2_3')
// (2, 20, 'lutff_2/in_3')
// (2, 20, 'sp4_r_v_b_11')
// (3, 6, 'sp4_v_t_43')
// (3, 7, 'sp4_v_b_43')
// (3, 8, 'sp4_v_b_30')
// (3, 9, 'sp4_v_b_19')
// (3, 10, 'sp4_v_b_6')
// (3, 10, 'sp4_v_t_38')
// (3, 10, 'sp4_v_t_43')
// (3, 11, 'sp4_r_v_b_40')
// (3, 11, 'sp4_v_b_38')
// (3, 11, 'sp4_v_b_43')
// (3, 12, 'sp4_r_v_b_29')
// (3, 12, 'sp4_v_b_27')
// (3, 12, 'sp4_v_b_30')
// (3, 13, 'sp4_r_v_b_16')
// (3, 13, 'sp4_v_b_14')
// (3, 13, 'sp4_v_b_19')
// (3, 14, 'sp4_r_v_b_5')
// (3, 14, 'sp4_v_b_3')
// (3, 14, 'sp4_v_b_6')
// (3, 14, 'sp4_v_t_38')
// (3, 15, 'local_g3_6')
// (3, 15, 'lutff_3/in_2')
// (3, 15, 'sp4_r_v_b_39')
// (3, 15, 'sp4_v_b_38')
// (3, 16, 'neigh_op_top_7')
// (3, 16, 'sp4_r_v_b_26')
// (3, 16, 'sp4_v_b_27')
// (3, 16, 'sp4_v_t_46')
// (3, 17, 'lutff_7/out')
// (3, 17, 'sp4_h_r_30')
// (3, 17, 'sp4_r_v_b_15')
// (3, 17, 'sp4_v_b_14')
// (3, 17, 'sp4_v_b_46')
// (3, 18, 'local_g1_7')
// (3, 18, 'lutff_7/in_3')
// (3, 18, 'neigh_op_bot_7')
// (3, 18, 'sp4_r_v_b_2')
// (3, 18, 'sp4_v_b_3')
// (3, 18, 'sp4_v_b_35')
// (3, 19, 'sp4_v_b_22')
// (3, 20, 'sp4_v_b_11')
// (4, 10, 'sp4_v_t_40')
// (4, 11, 'sp4_v_b_40')
// (4, 12, 'sp4_v_b_29')
// (4, 13, 'local_g0_0')
// (4, 13, 'lutff_6/in_2')
// (4, 13, 'sp4_v_b_16')
// (4, 14, 'local_g0_2')
// (4, 14, 'lutff_7/in_1')
// (4, 14, 'sp4_h_r_2')
// (4, 14, 'sp4_v_b_5')
// (4, 14, 'sp4_v_t_39')
// (4, 15, 'sp4_v_b_39')
// (4, 16, 'neigh_op_tnl_7')
// (4, 16, 'sp4_v_b_26')
// (4, 17, 'local_g0_7')
// (4, 17, 'lutff_2/in_3')
// (4, 17, 'neigh_op_lft_7')
// (4, 17, 'sp4_h_r_43')
// (4, 17, 'sp4_v_b_15')
// (4, 18, 'neigh_op_bnl_7')
// (4, 18, 'sp4_v_b_2')
// (5, 14, 'sp4_h_r_15')
// (5, 17, 'sp4_h_l_43')
// (6, 14, 'sp4_h_r_26')
// (7, 14, 'sp4_h_r_39')
// (8, 14, 'sp4_h_l_39')

wire n143;
// (0, 19, 'neigh_op_tnr_1')
// (0, 20, 'neigh_op_rgt_1')
// (0, 21, 'neigh_op_bnr_1')
// (1, 19, 'neigh_op_top_1')
// (1, 20, 'local_g1_1')
// (1, 20, 'lutff_1/out')
// (1, 20, 'lutff_4/in_2')
// (1, 21, 'neigh_op_bot_1')
// (2, 19, 'neigh_op_tnl_1')
// (2, 20, 'neigh_op_lft_1')
// (2, 21, 'neigh_op_bnl_1')

wire n144;
// (0, 19, 'neigh_op_tnr_2')
// (0, 20, 'neigh_op_rgt_2')
// (0, 21, 'neigh_op_bnr_2')
// (1, 19, 'neigh_op_top_2')
// (1, 20, 'local_g1_2')
// (1, 20, 'lutff_2/out')
// (1, 20, 'lutff_6/in_1')
// (1, 21, 'neigh_op_bot_2')
// (2, 19, 'neigh_op_tnl_2')
// (2, 20, 'neigh_op_lft_2')
// (2, 21, 'neigh_op_bnl_2')

wire n145;
// (0, 19, 'neigh_op_tnr_3')
// (0, 20, 'neigh_op_rgt_3')
// (0, 21, 'neigh_op_bnr_3')
// (1, 19, 'neigh_op_top_3')
// (1, 20, 'local_g3_3')
// (1, 20, 'lutff_3/out')
// (1, 20, 'lutff_5/in_3')
// (1, 21, 'neigh_op_bot_3')
// (2, 19, 'neigh_op_tnl_3')
// (2, 20, 'neigh_op_lft_3')
// (2, 21, 'neigh_op_bnl_3')

reg n146 = 0;
// (0, 19, 'neigh_op_tnr_4')
// (0, 20, 'neigh_op_rgt_4')
// (0, 21, 'neigh_op_bnr_4')
// (1, 19, 'neigh_op_top_4')
// (1, 20, 'local_g0_4')
// (1, 20, 'lutff_1/in_1')
// (1, 20, 'lutff_3/in_3')
// (1, 20, 'lutff_4/out')
// (1, 21, 'neigh_op_bot_4')
// (2, 19, 'neigh_op_tnl_4')
// (2, 20, 'local_g0_4')
// (2, 20, 'lutff_7/in_1')
// (2, 20, 'neigh_op_lft_4')
// (2, 21, 'neigh_op_bnl_4')

wire n147;
// (0, 19, 'neigh_op_tnr_5')
// (0, 20, 'neigh_op_rgt_5')
// (0, 21, 'neigh_op_bnr_5')
// (1, 19, 'neigh_op_top_5')
// (1, 20, 'local_g0_2')
// (1, 20, 'lutff_5/out')
// (1, 20, 'lutff_global/cen')
// (1, 20, 'sp4_h_r_10')
// (1, 21, 'neigh_op_bot_5')
// (2, 19, 'neigh_op_tnl_5')
// (2, 20, 'neigh_op_lft_5')
// (2, 20, 'sp4_h_r_23')
// (2, 21, 'neigh_op_bnl_5')
// (3, 20, 'sp4_h_r_34')
// (4, 20, 'sp4_h_r_47')
// (5, 20, 'sp4_h_l_47')

reg n148 = 0;
// (0, 19, 'neigh_op_tnr_6')
// (0, 20, 'neigh_op_rgt_6')
// (0, 21, 'neigh_op_bnr_6')
// (1, 19, 'neigh_op_top_6')
// (1, 20, 'local_g0_6')
// (1, 20, 'lutff_2/in_2')
// (1, 20, 'lutff_3/in_1')
// (1, 20, 'lutff_6/out')
// (1, 21, 'neigh_op_bot_6')
// (2, 19, 'neigh_op_tnl_6')
// (2, 20, 'local_g0_6')
// (2, 20, 'lutff_7/in_3')
// (2, 20, 'neigh_op_lft_6')
// (2, 21, 'neigh_op_bnl_6')

reg n149 = 0;
// (0, 19, 'neigh_op_tnr_7')
// (0, 20, 'neigh_op_rgt_7')
// (0, 21, 'neigh_op_bnr_7')
// (1, 19, 'neigh_op_top_7')
// (1, 19, 'sp4_r_v_b_42')
// (1, 20, 'local_g0_7')
// (1, 20, 'local_g1_7')
// (1, 20, 'lutff_0/in_2')
// (1, 20, 'lutff_1/in_3')
// (1, 20, 'lutff_7/in_0')
// (1, 20, 'lutff_7/out')
// (1, 20, 'sp4_r_v_b_31')
// (1, 21, 'neigh_op_bot_7')
// (1, 21, 'sp4_r_v_b_18')
// (1, 22, 'sp4_r_v_b_7')
// (2, 18, 'sp4_v_t_42')
// (2, 19, 'neigh_op_tnl_7')
// (2, 19, 'sp4_v_b_42')
// (2, 20, 'local_g2_7')
// (2, 20, 'lutff_7/in_0')
// (2, 20, 'neigh_op_lft_7')
// (2, 20, 'sp4_v_b_31')
// (2, 21, 'neigh_op_bnl_7')
// (2, 21, 'sp4_v_b_18')
// (2, 22, 'sp4_v_b_7')

wire n150;
// (0, 19, 'sp4_h_r_12')
// (1, 19, 'local_g2_1')
// (1, 19, 'local_g2_6')
// (1, 19, 'lutff_1/in_0')
// (1, 19, 'lutff_2/in_0')
// (1, 19, 'lutff_6/in_0')
// (1, 19, 'lutff_7/in_3')
// (1, 19, 'sp4_h_r_25')
// (1, 19, 'sp4_r_v_b_38')
// (1, 20, 'local_g2_7')
// (1, 20, 'lutff_4/in_1')
// (1, 20, 'lutff_5/in_0')
// (1, 20, 'lutff_6/in_3')
// (1, 20, 'lutff_7/in_2')
// (1, 20, 'neigh_op_tnr_7')
// (1, 20, 'sp4_r_v_b_27')
// (1, 21, 'neigh_op_rgt_7')
// (1, 21, 'sp4_r_v_b_14')
// (1, 22, 'neigh_op_bnr_7')
// (1, 22, 'sp4_r_v_b_3')
// (2, 18, 'sp4_v_t_38')
// (2, 19, 'sp4_h_r_36')
// (2, 19, 'sp4_v_b_38')
// (2, 20, 'local_g1_7')
// (2, 20, 'lutff_0/in_0')
// (2, 20, 'lutff_1/in_3')
// (2, 20, 'lutff_3/in_3')
// (2, 20, 'neigh_op_top_7')
// (2, 20, 'sp4_r_v_b_42')
// (2, 20, 'sp4_v_b_27')
// (2, 21, 'local_g0_7')
// (2, 21, 'local_g3_7')
// (2, 21, 'lutff_1/in_0')
// (2, 21, 'lutff_2/in_2')
// (2, 21, 'lutff_3/in_2')
// (2, 21, 'lutff_7/out')
// (2, 21, 'sp4_r_v_b_31')
// (2, 21, 'sp4_v_b_14')
// (2, 22, 'neigh_op_bot_7')
// (2, 22, 'sp4_r_v_b_18')
// (2, 22, 'sp4_v_b_3')
// (2, 23, 'sp4_r_v_b_7')
// (3, 19, 'sp4_h_l_36')
// (3, 19, 'sp4_v_t_42')
// (3, 20, 'neigh_op_tnl_7')
// (3, 20, 'sp4_v_b_42')
// (3, 21, 'neigh_op_lft_7')
// (3, 21, 'sp4_v_b_31')
// (3, 22, 'neigh_op_bnl_7')
// (3, 22, 'sp4_v_b_18')
// (3, 23, 'sp4_v_b_7')

reg n151 = 0;
// (0, 19, 'sp4_h_r_21')
// (1, 19, 'local_g3_0')
// (1, 19, 'lutff_4/in_1')
// (1, 19, 'sp4_h_r_32')
// (2, 10, 'sp4_r_v_b_38')
// (2, 11, 'sp4_r_v_b_27')
// (2, 12, 'local_g2_6')
// (2, 12, 'lutff_3/in_3')
// (2, 12, 'sp4_r_v_b_14')
// (2, 13, 'sp4_r_v_b_3')
// (2, 14, 'local_g3_2')
// (2, 14, 'lutff_7/in_2')
// (2, 14, 'sp4_r_v_b_42')
// (2, 15, 'local_g0_7')
// (2, 15, 'lutff_0/in_1')
// (2, 15, 'sp4_r_v_b_31')
// (2, 16, 'sp4_r_v_b_18')
// (2, 16, 'sp4_r_v_b_40')
// (2, 17, 'sp4_r_v_b_29')
// (2, 17, 'sp4_r_v_b_7')
// (2, 18, 'local_g3_0')
// (2, 18, 'lutff_4/in_1')
// (2, 18, 'sp4_r_v_b_16')
// (2, 18, 'sp4_r_v_b_46')
// (2, 19, 'sp4_h_r_45')
// (2, 19, 'sp4_r_v_b_35')
// (2, 19, 'sp4_r_v_b_5')
// (2, 20, 'local_g3_6')
// (2, 20, 'lutff_7/in_2')
// (2, 20, 'sp4_r_v_b_22')
// (2, 21, 'sp4_r_v_b_11')
// (3, 9, 'sp4_v_t_38')
// (3, 10, 'sp4_v_b_38')
// (3, 11, 'sp4_v_b_27')
// (3, 12, 'sp4_v_b_14')
// (3, 13, 'sp4_v_b_3')
// (3, 13, 'sp4_v_t_42')
// (3, 14, 'sp4_v_b_42')
// (3, 15, 'sp4_v_b_31')
// (3, 15, 'sp4_v_t_40')
// (3, 16, 'sp4_v_b_18')
// (3, 16, 'sp4_v_b_40')
// (3, 17, 'sp4_h_r_2')
// (3, 17, 'sp4_v_b_29')
// (3, 17, 'sp4_v_b_7')
// (3, 17, 'sp4_v_t_46')
// (3, 18, 'sp4_r_v_b_47')
// (3, 18, 'sp4_v_b_16')
// (3, 18, 'sp4_v_b_46')
// (3, 19, 'local_g0_1')
// (3, 19, 'lutff_7/in_0')
// (3, 19, 'sp4_h_l_45')
// (3, 19, 'sp4_h_r_0')
// (3, 19, 'sp4_r_v_b_34')
// (3, 19, 'sp4_v_b_35')
// (3, 19, 'sp4_v_b_5')
// (3, 20, 'sp4_r_v_b_23')
// (3, 20, 'sp4_v_b_22')
// (3, 21, 'sp4_h_r_11')
// (3, 21, 'sp4_r_v_b_10')
// (3, 21, 'sp4_v_b_11')
// (4, 14, 'local_g3_0')
// (4, 14, 'lutff_7/in_2')
// (4, 14, 'sp4_r_v_b_40')
// (4, 15, 'sp4_r_v_b_29')
// (4, 16, 'sp4_r_v_b_16')
// (4, 17, 'sp4_h_r_15')
// (4, 17, 'sp4_r_v_b_5')
// (4, 17, 'sp4_v_t_47')
// (4, 18, 'sp4_r_v_b_40')
// (4, 18, 'sp4_v_b_47')
// (4, 19, 'sp4_h_r_13')
// (4, 19, 'sp4_r_v_b_29')
// (4, 19, 'sp4_v_b_34')
// (4, 20, 'sp4_r_v_b_16')
// (4, 20, 'sp4_v_b_23')
// (4, 21, 'sp4_h_r_22')
// (4, 21, 'sp4_h_r_5')
// (4, 21, 'sp4_r_v_b_5')
// (4, 21, 'sp4_v_b_10')
// (5, 13, 'sp4_v_t_40')
// (5, 14, 'sp4_v_b_40')
// (5, 15, 'sp4_v_b_29')
// (5, 16, 'local_g0_0')
// (5, 16, 'lutff_7/in_1')
// (5, 16, 'sp4_v_b_16')
// (5, 17, 'sp4_h_r_26')
// (5, 17, 'sp4_v_b_5')
// (5, 17, 'sp4_v_t_40')
// (5, 18, 'sp4_v_b_40')
// (5, 19, 'sp4_h_r_24')
// (5, 19, 'sp4_v_b_29')
// (5, 20, 'sp4_v_b_16')
// (5, 21, 'sp4_h_r_0')
// (5, 21, 'sp4_h_r_16')
// (5, 21, 'sp4_h_r_35')
// (5, 21, 'sp4_v_b_5')
// (6, 17, 'sp4_h_r_39')
// (6, 18, 'sp4_r_v_b_45')
// (6, 19, 'sp4_h_r_37')
// (6, 19, 'sp4_r_v_b_32')
// (6, 20, 'neigh_op_tnr_4')
// (6, 20, 'sp4_r_v_b_21')
// (6, 20, 'sp4_r_v_b_37')
// (6, 21, 'neigh_op_rgt_4')
// (6, 21, 'sp4_h_r_13')
// (6, 21, 'sp4_h_r_29')
// (6, 21, 'sp4_h_r_46')
// (6, 21, 'sp4_r_v_b_24')
// (6, 21, 'sp4_r_v_b_8')
// (6, 22, 'neigh_op_bnr_4')
// (6, 22, 'sp4_r_v_b_13')
// (6, 23, 'sp4_r_v_b_0')
// (7, 17, 'sp4_h_l_39')
// (7, 17, 'sp4_v_t_45')
// (7, 18, 'sp4_r_v_b_44')
// (7, 18, 'sp4_v_b_45')
// (7, 19, 'sp4_h_l_37')
// (7, 19, 'sp4_r_v_b_33')
// (7, 19, 'sp4_v_b_32')
// (7, 19, 'sp4_v_t_37')
// (7, 20, 'neigh_op_top_4')
// (7, 20, 'sp4_r_v_b_20')
// (7, 20, 'sp4_v_b_21')
// (7, 20, 'sp4_v_b_37')
// (7, 21, 'local_g2_4')
// (7, 21, 'lutff_4/in_0')
// (7, 21, 'lutff_4/out')
// (7, 21, 'sp4_h_l_46')
// (7, 21, 'sp4_h_r_24')
// (7, 21, 'sp4_h_r_40')
// (7, 21, 'sp4_h_r_8')
// (7, 21, 'sp4_r_v_b_9')
// (7, 21, 'sp4_v_b_24')
// (7, 21, 'sp4_v_b_8')
// (7, 22, 'neigh_op_bot_4')
// (7, 22, 'sp4_v_b_13')
// (7, 23, 'sp4_v_b_0')
// (8, 17, 'sp4_h_r_9')
// (8, 17, 'sp4_v_t_44')
// (8, 18, 'sp4_v_b_44')
// (8, 19, 'sp4_v_b_33')
// (8, 20, 'neigh_op_tnl_4')
// (8, 20, 'sp4_v_b_20')
// (8, 21, 'neigh_op_lft_4')
// (8, 21, 'sp4_h_l_40')
// (8, 21, 'sp4_h_r_21')
// (8, 21, 'sp4_h_r_37')
// (8, 21, 'sp4_v_b_9')
// (8, 22, 'neigh_op_bnl_4')
// (9, 17, 'sp4_h_r_20')
// (9, 21, 'sp4_h_l_37')
// (9, 21, 'sp4_h_r_32')
// (10, 17, 'sp4_h_r_33')
// (10, 18, 'sp4_r_v_b_39')
// (10, 19, 'sp4_r_v_b_26')
// (10, 20, 'sp4_r_v_b_15')
// (10, 21, 'sp4_h_r_45')
// (10, 21, 'sp4_r_v_b_2')
// (11, 17, 'local_g3_4')
// (11, 17, 'lutff_2/in_3')
// (11, 17, 'sp4_h_r_44')
// (11, 17, 'sp4_v_t_39')
// (11, 18, 'local_g3_7')
// (11, 18, 'lutff_6/in_2')
// (11, 18, 'sp4_v_b_39')
// (11, 19, 'sp4_v_b_26')
// (11, 20, 'sp4_v_b_15')
// (11, 21, 'sp4_h_l_45')
// (11, 21, 'sp4_v_b_2')
// (12, 17, 'sp4_h_l_44')

reg n152 = 0;
// (0, 20, 'neigh_op_tnr_1')
// (0, 21, 'neigh_op_rgt_1')
// (0, 22, 'neigh_op_bnr_1')
// (1, 20, 'neigh_op_top_1')
// (1, 21, 'local_g1_1')
// (1, 21, 'lutff_1/in_1')
// (1, 21, 'lutff_1/out')
// (1, 21, 'lutff_5/in_1')
// (1, 21, 'lutff_7/in_3')
// (1, 22, 'neigh_op_bot_1')
// (2, 20, 'neigh_op_tnl_1')
// (2, 21, 'neigh_op_lft_1')
// (2, 22, 'neigh_op_bnl_1')

reg n153 = 0;
// (0, 20, 'neigh_op_tnr_2')
// (0, 21, 'neigh_op_rgt_2')
// (0, 22, 'neigh_op_bnr_2')
// (1, 20, 'neigh_op_top_2')
// (1, 21, 'local_g2_2')
// (1, 21, 'local_g3_2')
// (1, 21, 'lutff_2/in_1')
// (1, 21, 'lutff_2/out')
// (1, 21, 'lutff_5/in_0')
// (1, 21, 'lutff_7/in_1')
// (1, 22, 'neigh_op_bot_2')
// (2, 20, 'neigh_op_tnl_2')
// (2, 21, 'neigh_op_lft_2')
// (2, 22, 'neigh_op_bnl_2')

reg n154 = 0;
// (0, 20, 'neigh_op_tnr_3')
// (0, 21, 'neigh_op_rgt_3')
// (0, 22, 'neigh_op_bnr_3')
// (1, 20, 'neigh_op_top_3')
// (1, 21, 'local_g0_3')
// (1, 21, 'lutff_3/in_0')
// (1, 21, 'lutff_3/out')
// (1, 21, 'lutff_5/in_2')
// (1, 21, 'lutff_7/in_2')
// (1, 22, 'neigh_op_bot_3')
// (2, 20, 'neigh_op_tnl_3')
// (2, 21, 'neigh_op_lft_3')
// (2, 22, 'neigh_op_bnl_3')

wire n155;
// (0, 20, 'neigh_op_tnr_5')
// (0, 21, 'neigh_op_rgt_5')
// (0, 22, 'neigh_op_bnr_5')
// (1, 20, 'neigh_op_top_5')
// (1, 21, 'lutff_5/out')
// (1, 22, 'neigh_op_bot_5')
// (2, 20, 'neigh_op_tnl_5')
// (2, 21, 'local_g1_5')
// (2, 21, 'lutff_6/in_2')
// (2, 21, 'neigh_op_lft_5')
// (2, 22, 'neigh_op_bnl_5')

reg n156 = 0;
// (0, 20, 'neigh_op_tnr_6')
// (0, 21, 'neigh_op_rgt_6')
// (0, 22, 'neigh_op_bnr_6')
// (1, 20, 'neigh_op_top_6')
// (1, 21, 'local_g0_6')
// (1, 21, 'lutff_0/in_2')
// (1, 21, 'lutff_1/in_3')
// (1, 21, 'lutff_5/in_3')
// (1, 21, 'lutff_6/in_2')
// (1, 21, 'lutff_6/out')
// (1, 22, 'neigh_op_bot_6')
// (2, 20, 'neigh_op_tnl_6')
// (2, 21, 'neigh_op_lft_6')
// (2, 22, 'neigh_op_bnl_6')

wire n157;
// (0, 20, 'neigh_op_tnr_7')
// (0, 21, 'neigh_op_rgt_7')
// (0, 22, 'neigh_op_bnr_7')
// (1, 20, 'neigh_op_top_7')
// (1, 21, 'local_g1_7')
// (1, 21, 'local_g2_7')
// (1, 21, 'lutff_1/in_0')
// (1, 21, 'lutff_2/in_0')
// (1, 21, 'lutff_3/in_2')
// (1, 21, 'lutff_6/in_3')
// (1, 21, 'lutff_7/out')
// (1, 22, 'neigh_op_bot_7')
// (2, 20, 'neigh_op_tnl_7')
// (2, 21, 'neigh_op_lft_7')
// (2, 22, 'neigh_op_bnl_7')

wire n158;
// (0, 20, 'sp4_h_r_0')
// (1, 17, 'sp4_r_v_b_45')
// (1, 18, 'sp4_r_v_b_32')
// (1, 19, 'neigh_op_tnr_4')
// (1, 19, 'sp4_r_v_b_21')
// (1, 20, 'neigh_op_rgt_4')
// (1, 20, 'sp4_h_r_13')
// (1, 20, 'sp4_r_v_b_8')
// (1, 21, 'neigh_op_bnr_4')
// (2, 16, 'sp4_v_t_45')
// (2, 17, 'local_g3_5')
// (2, 17, 'lutff_4/in_0')
// (2, 17, 'sp4_v_b_45')
// (2, 18, 'local_g2_0')
// (2, 18, 'lutff_5/in_1')
// (2, 18, 'sp4_v_b_32')
// (2, 19, 'neigh_op_top_4')
// (2, 19, 'sp4_v_b_21')
// (2, 20, 'lutff_4/out')
// (2, 20, 'sp4_h_r_24')
// (2, 20, 'sp4_v_b_8')
// (2, 21, 'neigh_op_bot_4')
// (3, 17, 'sp4_r_v_b_43')
// (3, 18, 'sp4_r_v_b_30')
// (3, 19, 'neigh_op_tnl_4')
// (3, 19, 'sp4_r_v_b_19')
// (3, 20, 'neigh_op_lft_4')
// (3, 20, 'sp4_h_r_37')
// (3, 20, 'sp4_r_v_b_6')
// (3, 21, 'neigh_op_bnl_4')
// (4, 16, 'sp4_v_t_43')
// (4, 17, 'local_g2_3')
// (4, 17, 'lutff_4/in_1')
// (4, 17, 'sp4_v_b_43')
// (4, 18, 'sp4_v_b_30')
// (4, 19, 'sp4_v_b_19')
// (4, 20, 'sp4_h_l_37')
// (4, 20, 'sp4_h_r_3')
// (4, 20, 'sp4_v_b_6')
// (5, 20, 'sp4_h_r_14')
// (6, 20, 'sp4_h_r_27')
// (7, 20, 'sp4_h_r_38')
// (7, 21, 'sp4_r_v_b_38')
// (7, 22, 'sp4_r_v_b_27')
// (7, 23, 'sp4_r_v_b_14')
// (7, 24, 'sp4_r_v_b_3')
// (8, 20, 'sp4_h_l_38')
// (8, 20, 'sp4_v_t_38')
// (8, 21, 'local_g3_6')
// (8, 21, 'lutff_4/in_3')
// (8, 21, 'sp4_v_b_38')
// (8, 22, 'sp4_v_b_27')
// (8, 23, 'sp4_v_b_14')
// (8, 24, 'sp4_v_b_3')

wire n159;
// (0, 20, 'sp4_h_r_2')
// (1, 15, 'sp4_r_v_b_40')
// (1, 15, 'sp4_r_v_b_47')
// (1, 16, 'sp4_r_v_b_29')
// (1, 16, 'sp4_r_v_b_34')
// (1, 17, 'sp4_r_v_b_16')
// (1, 17, 'sp4_r_v_b_23')
// (1, 18, 'sp4_r_v_b_10')
// (1, 18, 'sp4_r_v_b_5')
// (1, 19, 'neigh_op_tnr_5')
// (1, 19, 'sp4_r_v_b_39')
// (1, 20, 'neigh_op_rgt_5')
// (1, 20, 'sp4_h_r_15')
// (1, 20, 'sp4_r_v_b_26')
// (1, 21, 'neigh_op_bnr_5')
// (1, 21, 'sp4_r_v_b_15')
// (1, 22, 'sp4_r_v_b_2')
// (2, 14, 'local_g1_2')
// (2, 14, 'lutff_1/in_0')
// (2, 14, 'lutff_4/in_1')
// (2, 14, 'sp4_h_r_10')
// (2, 14, 'sp4_v_t_40')
// (2, 14, 'sp4_v_t_47')
// (2, 15, 'local_g3_0')
// (2, 15, 'lutff_1/in_2')
// (2, 15, 'sp4_r_v_b_46')
// (2, 15, 'sp4_v_b_40')
// (2, 15, 'sp4_v_b_47')
// (2, 16, 'sp4_r_v_b_35')
// (2, 16, 'sp4_v_b_29')
// (2, 16, 'sp4_v_b_34')
// (2, 17, 'sp4_r_v_b_22')
// (2, 17, 'sp4_v_b_16')
// (2, 17, 'sp4_v_b_23')
// (2, 18, 'sp4_h_r_7')
// (2, 18, 'sp4_r_v_b_11')
// (2, 18, 'sp4_v_b_10')
// (2, 18, 'sp4_v_b_5')
// (2, 18, 'sp4_v_t_39')
// (2, 19, 'neigh_op_top_5')
// (2, 19, 'sp4_r_v_b_38')
// (2, 19, 'sp4_v_b_39')
// (2, 20, 'lutff_5/out')
// (2, 20, 'sp4_h_r_26')
// (2, 20, 'sp4_r_v_b_27')
// (2, 20, 'sp4_v_b_26')
// (2, 21, 'local_g0_5')
// (2, 21, 'lutff_7/in_0')
// (2, 21, 'neigh_op_bot_5')
// (2, 21, 'sp4_r_v_b_14')
// (2, 21, 'sp4_v_b_15')
// (2, 22, 'sp4_r_v_b_3')
// (2, 22, 'sp4_v_b_2')
// (3, 14, 'sp4_h_r_23')
// (3, 14, 'sp4_v_t_46')
// (3, 15, 'sp4_v_b_46')
// (3, 16, 'local_g2_3')
// (3, 16, 'lutff_6/in_1')
// (3, 16, 'sp4_v_b_35')
// (3, 17, 'local_g1_6')
// (3, 17, 'lutff_7/in_0')
// (3, 17, 'sp4_r_v_b_39')
// (3, 17, 'sp4_v_b_22')
// (3, 18, 'sp4_h_r_18')
// (3, 18, 'sp4_r_v_b_26')
// (3, 18, 'sp4_v_b_11')
// (3, 18, 'sp4_v_t_38')
// (3, 19, 'neigh_op_tnl_5')
// (3, 19, 'sp4_r_v_b_15')
// (3, 19, 'sp4_v_b_38')
// (3, 20, 'neigh_op_lft_5')
// (3, 20, 'sp4_h_r_39')
// (3, 20, 'sp4_r_v_b_2')
// (3, 20, 'sp4_v_b_27')
// (3, 21, 'neigh_op_bnl_5')
// (3, 21, 'sp4_v_b_14')
// (3, 22, 'sp4_h_r_3')
// (3, 22, 'sp4_v_b_3')
// (4, 14, 'sp4_h_r_34')
// (4, 16, 'sp4_h_r_2')
// (4, 16, 'sp4_v_t_39')
// (4, 17, 'local_g2_7')
// (4, 17, 'lutff_4/in_3')
// (4, 17, 'sp4_v_b_39')
// (4, 18, 'sp4_h_r_31')
// (4, 18, 'sp4_v_b_26')
// (4, 19, 'sp4_v_b_15')
// (4, 20, 'sp4_h_l_39')
// (4, 20, 'sp4_v_b_2')
// (4, 22, 'sp4_h_r_14')
// (5, 14, 'sp4_h_r_47')
// (5, 15, 'sp4_r_v_b_42')
// (5, 16, 'sp4_h_r_15')
// (5, 16, 'sp4_r_v_b_31')
// (5, 17, 'local_g3_2')
// (5, 17, 'lutff_0/in_3')
// (5, 17, 'sp4_r_v_b_18')
// (5, 18, 'sp4_h_r_42')
// (5, 18, 'sp4_r_v_b_7')
// (5, 22, 'sp4_h_r_27')
// (6, 14, 'sp4_h_l_47')
// (6, 14, 'sp4_v_t_42')
// (6, 15, 'sp4_v_b_42')
// (6, 16, 'sp4_h_r_26')
// (6, 16, 'sp4_v_b_31')
// (6, 17, 'sp4_v_b_18')
// (6, 18, 'sp4_h_l_42')
// (6, 18, 'sp4_v_b_7')
// (6, 19, 'sp4_r_v_b_44')
// (6, 20, 'sp4_r_v_b_33')
// (6, 21, 'sp4_r_v_b_20')
// (6, 22, 'sp4_h_r_38')
// (6, 22, 'sp4_r_v_b_9')
// (7, 16, 'sp4_h_r_39')
// (7, 18, 'sp4_v_t_44')
// (7, 19, 'sp4_v_b_44')
// (7, 20, 'sp4_v_b_33')
// (7, 21, 'local_g0_4')
// (7, 21, 'lutff_5/in_1')
// (7, 21, 'sp4_v_b_20')
// (7, 22, 'sp4_h_l_38')
// (7, 22, 'sp4_v_b_9')
// (8, 16, 'sp4_h_l_39')
// (8, 16, 'sp4_h_r_2')
// (9, 16, 'sp4_h_r_15')
// (10, 16, 'sp4_h_r_26')
// (11, 16, 'local_g2_7')
// (11, 16, 'lutff_5/in_0')
// (11, 16, 'sp4_h_r_39')
// (12, 16, 'sp4_h_l_39')

wire n160;
// (0, 21, 'sp4_h_r_19')
// (1, 19, 'neigh_op_tnr_1')
// (1, 20, 'neigh_op_rgt_1')
// (1, 21, 'neigh_op_bnr_1')
// (1, 21, 'sp4_h_r_30')
// (2, 18, 'sp4_r_v_b_43')
// (2, 19, 'neigh_op_top_1')
// (2, 19, 'sp4_r_v_b_30')
// (2, 20, 'lutff_1/out')
// (2, 20, 'sp4_r_v_b_19')
// (2, 21, 'local_g3_3')
// (2, 21, 'lutff_global/cen')
// (2, 21, 'neigh_op_bot_1')
// (2, 21, 'sp4_h_r_43')
// (2, 21, 'sp4_r_v_b_6')
// (3, 17, 'sp4_v_t_43')
// (3, 18, 'sp4_v_b_43')
// (3, 19, 'neigh_op_tnl_1')
// (3, 19, 'sp4_v_b_30')
// (3, 20, 'neigh_op_lft_1')
// (3, 20, 'sp4_v_b_19')
// (3, 21, 'neigh_op_bnl_1')
// (3, 21, 'sp4_h_l_43')
// (3, 21, 'sp4_v_b_6')

reg n161 = 0;
// (1, 0, 'logic_op_tnr_0')
// (1, 1, 'neigh_op_rgt_0')
// (1, 2, 'neigh_op_bnr_0')
// (2, 0, 'logic_op_top_0')
// (2, 1, 'local_g1_0')
// (2, 1, 'lutff_0/out')
// (2, 1, 'lutff_4/in_3')
// (2, 2, 'neigh_op_bot_0')
// (3, 0, 'logic_op_tnl_0')
// (3, 1, 'neigh_op_lft_0')
// (3, 2, 'neigh_op_bnl_0')

reg n162 = 0;
// (1, 0, 'logic_op_tnr_2')
// (1, 1, 'neigh_op_rgt_2')
// (1, 2, 'neigh_op_bnr_2')
// (2, 0, 'logic_op_top_2')
// (2, 1, 'local_g0_2')
// (2, 1, 'lutff_2/out')
// (2, 1, 'lutff_6/in_2')
// (2, 2, 'neigh_op_bot_2')
// (3, 0, 'logic_op_tnl_2')
// (3, 1, 'neigh_op_lft_2')
// (3, 2, 'neigh_op_bnl_2')

wire n163;
// (1, 0, 'logic_op_tnr_4')
// (1, 1, 'neigh_op_rgt_4')
// (1, 2, 'neigh_op_bnr_4')
// (2, 0, 'logic_op_top_4')
// (2, 1, 'lutff_4/out')
// (2, 2, 'local_g0_4')
// (2, 2, 'lutff_1/in_3')
// (2, 2, 'neigh_op_bot_4')
// (3, 0, 'logic_op_tnl_4')
// (3, 1, 'neigh_op_lft_4')
// (3, 2, 'neigh_op_bnl_4')

reg n164 = 0;
// (1, 0, 'logic_op_tnr_5')
// (1, 1, 'neigh_op_rgt_5')
// (1, 2, 'neigh_op_bnr_5')
// (2, 0, 'logic_op_top_5')
// (2, 1, 'local_g0_5')
// (2, 1, 'lutff_4/in_1')
// (2, 1, 'lutff_5/out')
// (2, 2, 'neigh_op_bot_5')
// (3, 0, 'logic_op_tnl_5')
// (3, 1, 'neigh_op_lft_5')
// (3, 2, 'neigh_op_bnl_5')

wire n165;
// (1, 0, 'logic_op_tnr_6')
// (1, 1, 'neigh_op_rgt_6')
// (1, 2, 'neigh_op_bnr_6')
// (2, 0, 'logic_op_top_6')
// (2, 1, 'lutff_6/out')
// (2, 2, 'local_g0_6')
// (2, 2, 'lutff_2/in_2')
// (2, 2, 'neigh_op_bot_6')
// (3, 0, 'logic_op_tnl_6')
// (3, 1, 'neigh_op_lft_6')
// (3, 2, 'neigh_op_bnl_6')

reg n166 = 0;
// (1, 0, 'logic_op_tnr_7')
// (1, 1, 'neigh_op_rgt_7')
// (1, 2, 'neigh_op_bnr_7')
// (2, 0, 'logic_op_top_7')
// (2, 1, 'local_g2_7')
// (2, 1, 'lutff_6/in_3')
// (2, 1, 'lutff_7/out')
// (2, 2, 'neigh_op_bot_7')
// (3, 0, 'logic_op_tnl_7')
// (3, 1, 'neigh_op_lft_7')
// (3, 2, 'neigh_op_bnl_7')

wire n167;
// (1, 1, 'neigh_op_tnr_0')
// (1, 2, 'neigh_op_rgt_0')
// (1, 3, 'neigh_op_bnr_0')
// (2, 1, 'neigh_op_top_0')
// (2, 2, 'local_g1_0')
// (2, 2, 'lutff_0/out')
// (2, 2, 'lutff_1/in_2')
// (2, 3, 'neigh_op_bot_0')
// (3, 1, 'neigh_op_tnl_0')
// (3, 2, 'neigh_op_lft_0')
// (3, 3, 'neigh_op_bnl_0')

wire n168;
// (1, 1, 'neigh_op_tnr_1')
// (1, 2, 'neigh_op_rgt_1')
// (1, 3, 'neigh_op_bnr_1')
// (2, 1, 'neigh_op_top_1')
// (2, 2, 'lutff_1/out')
// (2, 3, 'neigh_op_bot_1')
// (3, 1, 'neigh_op_tnl_1')
// (3, 2, 'local_g0_1')
// (3, 2, 'lutff_7/in_0')
// (3, 2, 'neigh_op_lft_1')
// (3, 3, 'neigh_op_bnl_1')

wire n169;
// (1, 1, 'neigh_op_tnr_2')
// (1, 2, 'neigh_op_rgt_2')
// (1, 3, 'neigh_op_bnr_2')
// (2, 1, 'neigh_op_top_2')
// (2, 2, 'local_g2_2')
// (2, 2, 'lutff_1/in_1')
// (2, 2, 'lutff_2/out')
// (2, 3, 'neigh_op_bot_2')
// (3, 1, 'neigh_op_tnl_2')
// (3, 2, 'neigh_op_lft_2')
// (3, 3, 'neigh_op_bnl_2')

reg n170 = 0;
// (1, 1, 'neigh_op_tnr_3')
// (1, 2, 'neigh_op_rgt_3')
// (1, 3, 'neigh_op_bnr_3')
// (2, 1, 'neigh_op_top_3')
// (2, 2, 'local_g2_3')
// (2, 2, 'lutff_0/in_3')
// (2, 2, 'lutff_3/out')
// (2, 3, 'neigh_op_bot_3')
// (3, 1, 'neigh_op_tnl_3')
// (3, 2, 'neigh_op_lft_3')
// (3, 3, 'neigh_op_bnl_3')

reg n171 = 0;
// (1, 1, 'neigh_op_tnr_4')
// (1, 2, 'neigh_op_rgt_4')
// (1, 3, 'neigh_op_bnr_4')
// (2, 1, 'neigh_op_top_4')
// (2, 2, 'local_g2_4')
// (2, 2, 'lutff_4/out')
// (2, 2, 'lutff_5/in_1')
// (2, 3, 'neigh_op_bot_4')
// (3, 1, 'neigh_op_tnl_4')
// (3, 2, 'neigh_op_lft_4')
// (3, 3, 'neigh_op_bnl_4')

wire n172;
// (1, 1, 'neigh_op_tnr_5')
// (1, 2, 'neigh_op_rgt_5')
// (1, 3, 'neigh_op_bnr_5')
// (2, 1, 'neigh_op_top_5')
// (2, 2, 'local_g0_5')
// (2, 2, 'lutff_2/in_1')
// (2, 2, 'lutff_5/out')
// (2, 3, 'neigh_op_bot_5')
// (3, 1, 'neigh_op_tnl_5')
// (3, 2, 'neigh_op_lft_5')
// (3, 3, 'neigh_op_bnl_5')

reg n173 = 0;
// (1, 1, 'neigh_op_tnr_6')
// (1, 2, 'neigh_op_rgt_6')
// (1, 3, 'neigh_op_bnr_6')
// (2, 1, 'neigh_op_top_6')
// (2, 2, 'local_g1_6')
// (2, 2, 'lutff_5/in_2')
// (2, 2, 'lutff_6/out')
// (2, 3, 'neigh_op_bot_6')
// (3, 1, 'neigh_op_tnl_6')
// (3, 2, 'neigh_op_lft_6')
// (3, 3, 'neigh_op_bnl_6')

reg n174 = 0;
// (1, 1, 'neigh_op_tnr_7')
// (1, 2, 'neigh_op_rgt_7')
// (1, 3, 'neigh_op_bnr_7')
// (2, 1, 'neigh_op_top_7')
// (2, 2, 'local_g1_7')
// (2, 2, 'lutff_0/in_0')
// (2, 2, 'lutff_7/out')
// (2, 3, 'neigh_op_bot_7')
// (3, 1, 'neigh_op_tnl_7')
// (3, 2, 'neigh_op_lft_7')
// (3, 3, 'neigh_op_bnl_7')

reg n175 = 0;
// (1, 1, 'sp4_h_r_2')
// (2, 1, 'local_g1_7')
// (2, 1, 'lutff_0/in_2')
// (2, 1, 'sp4_h_r_15')
// (3, 1, 'local_g2_2')
// (3, 1, 'lutff_6/in_0')
// (3, 1, 'sp4_h_r_26')
// (4, 1, 'sp4_h_r_39')
// (4, 2, 'local_g3_5')
// (4, 2, 'lutff_5/in_3')
// (4, 2, 'sp4_r_v_b_36')
// (4, 2, 'sp4_r_v_b_45')
// (4, 3, 'sp4_r_v_b_25')
// (4, 3, 'sp4_r_v_b_32')
// (4, 4, 'sp4_r_v_b_12')
// (4, 4, 'sp4_r_v_b_21')
// (4, 5, 'sp4_r_v_b_1')
// (4, 5, 'sp4_r_v_b_8')
// (4, 7, 'sp4_r_v_b_41')
// (4, 8, 'sp4_r_v_b_28')
// (4, 9, 'sp4_r_v_b_17')
// (4, 10, 'local_g1_4')
// (4, 10, 'lutff_1/in_0')
// (4, 10, 'sp4_r_v_b_4')
// (4, 13, 'sp4_r_v_b_38')
// (4, 14, 'sp4_r_v_b_27')
// (4, 15, 'sp4_r_v_b_14')
// (4, 16, 'sp4_r_v_b_3')
// (4, 17, 'sp4_r_v_b_46')
// (4, 18, 'sp4_r_v_b_35')
// (4, 19, 'sp4_r_v_b_22')
// (4, 20, 'local_g2_3')
// (4, 20, 'lutff_5/in_2')
// (4, 20, 'sp4_r_v_b_11')
// (5, 1, 'local_g0_3')
// (5, 1, 'lutff_4/in_3')
// (5, 1, 'sp4_h_l_39')
// (5, 1, 'sp4_h_r_11')
// (5, 1, 'sp4_v_t_36')
// (5, 1, 'sp4_v_t_45')
// (5, 2, 'sp4_v_b_36')
// (5, 2, 'sp4_v_b_45')
// (5, 3, 'local_g3_1')
// (5, 3, 'lutff_1/in_1')
// (5, 3, 'sp4_v_b_25')
// (5, 3, 'sp4_v_b_32')
// (5, 4, 'sp4_v_b_12')
// (5, 4, 'sp4_v_b_21')
// (5, 5, 'local_g0_0')
// (5, 5, 'lutff_2/in_2')
// (5, 5, 'sp4_h_r_3')
// (5, 5, 'sp4_h_r_8')
// (5, 5, 'sp4_v_b_1')
// (5, 5, 'sp4_v_b_8')
// (5, 6, 'sp4_r_v_b_42')
// (5, 6, 'sp4_v_t_41')
// (5, 7, 'local_g0_7')
// (5, 7, 'lutff_0/in_1')
// (5, 7, 'sp4_r_v_b_31')
// (5, 7, 'sp4_v_b_41')
// (5, 8, 'sp4_r_v_b_18')
// (5, 8, 'sp4_v_b_28')
// (5, 9, 'sp4_r_v_b_7')
// (5, 9, 'sp4_v_b_17')
// (5, 10, 'sp4_h_r_4')
// (5, 10, 'sp4_v_b_4')
// (5, 12, 'sp4_h_r_9')
// (5, 12, 'sp4_v_t_38')
// (5, 13, 'sp4_v_b_38')
// (5, 14, 'sp4_v_b_27')
// (5, 15, 'sp4_v_b_14')
// (5, 16, 'sp4_v_b_3')
// (5, 16, 'sp4_v_t_46')
// (5, 17, 'sp4_v_b_46')
// (5, 18, 'sp4_v_b_35')
// (5, 19, 'sp4_v_b_22')
// (5, 20, 'sp4_v_b_11')
// (6, 1, 'sp4_h_r_22')
// (6, 5, 'sp4_h_r_14')
// (6, 5, 'sp4_h_r_21')
// (6, 5, 'sp4_v_t_42')
// (6, 6, 'sp4_v_b_42')
// (6, 7, 'sp4_v_b_31')
// (6, 8, 'sp4_v_b_18')
// (6, 9, 'sp4_h_r_7')
// (6, 9, 'sp4_v_b_7')
// (6, 10, 'sp4_h_r_17')
// (6, 12, 'sp4_h_r_20')
// (7, 1, 'sp4_h_r_35')
// (7, 2, 'sp4_r_v_b_44')
// (7, 3, 'sp4_r_v_b_33')
// (7, 4, 'local_g3_4')
// (7, 4, 'lutff_4/in_1')
// (7, 4, 'sp4_r_v_b_20')
// (7, 5, 'sp4_h_r_27')
// (7, 5, 'sp4_h_r_32')
// (7, 5, 'sp4_r_v_b_9')
// (7, 9, 'sp4_h_r_18')
// (7, 10, 'sp4_h_r_28')
// (7, 10, 'sp4_r_v_b_46')
// (7, 11, 'sp4_r_v_b_35')
// (7, 12, 'sp4_h_r_33')
// (7, 12, 'sp4_r_v_b_22')
// (7, 13, 'sp4_r_v_b_11')
// (8, 1, 'sp4_h_r_46')
// (8, 1, 'sp4_v_t_44')
// (8, 2, 'sp4_v_b_44')
// (8, 3, 'sp4_v_b_33')
// (8, 4, 'sp4_v_b_20')
// (8, 5, 'local_g3_5')
// (8, 5, 'lutff_0/in_0')
// (8, 5, 'sp4_h_r_38')
// (8, 5, 'sp4_h_r_4')
// (8, 5, 'sp4_h_r_45')
// (8, 5, 'sp4_v_b_9')
// (8, 9, 'sp4_h_r_31')
// (8, 9, 'sp4_h_r_5')
// (8, 9, 'sp4_v_t_46')
// (8, 10, 'sp4_h_r_41')
// (8, 10, 'sp4_v_b_46')
// (8, 11, 'sp4_v_b_35')
// (8, 12, 'local_g1_6')
// (8, 12, 'lutff_2/in_3')
// (8, 12, 'sp4_h_r_44')
// (8, 12, 'sp4_v_b_22')
// (8, 13, 'sp4_v_b_11')
// (9, 1, 'sp4_h_l_46')
// (9, 1, 'sp4_h_r_3')
// (9, 2, 'sp4_r_v_b_40')
// (9, 2, 'sp4_r_v_b_44')
// (9, 3, 'sp4_r_v_b_29')
// (9, 3, 'sp4_r_v_b_33')
// (9, 4, 'sp4_r_v_b_16')
// (9, 4, 'sp4_r_v_b_20')
// (9, 5, 'local_g2_1')
// (9, 5, 'lutff_6/in_1')
// (9, 5, 'sp4_h_l_38')
// (9, 5, 'sp4_h_l_45')
// (9, 5, 'sp4_h_r_0')
// (9, 5, 'sp4_h_r_17')
// (9, 5, 'sp4_r_v_b_5')
// (9, 5, 'sp4_r_v_b_9')
// (9, 6, 'sp4_r_v_b_44')
// (9, 7, 'local_g2_1')
// (9, 7, 'lutff_5/in_2')
// (9, 7, 'sp4_r_v_b_33')
// (9, 8, 'sp4_r_v_b_20')
// (9, 9, 'sp4_h_r_16')
// (9, 9, 'sp4_h_r_42')
// (9, 9, 'sp4_r_v_b_9')
// (9, 10, 'sp4_h_l_41')
// (9, 10, 'sp4_h_r_1')
// (9, 12, 'sp4_h_l_44')
// (9, 12, 'sp4_h_r_1')
// (9, 14, 'local_g1_2')
// (9, 14, 'lutff_2/in_1')
// (9, 14, 'sp4_h_r_2')
// (9, 14, 'sp4_r_v_b_36')
// (9, 14, 'sp4_r_v_b_41')
// (9, 15, 'sp4_r_v_b_25')
// (9, 15, 'sp4_r_v_b_28')
// (9, 16, 'sp4_r_v_b_12')
// (9, 16, 'sp4_r_v_b_17')
// (9, 17, 'sp4_r_v_b_1')
// (9, 17, 'sp4_r_v_b_4')
// (9, 18, 'sp4_r_v_b_36')
// (9, 18, 'sp4_r_v_b_41')
// (9, 19, 'sp4_r_v_b_25')
// (9, 19, 'sp4_r_v_b_28')
// (9, 20, 'sp4_r_v_b_12')
// (9, 20, 'sp4_r_v_b_17')
// (9, 21, 'local_g1_1')
// (9, 21, 'lutff_5/in_1')
// (9, 21, 'sp4_r_v_b_1')
// (9, 21, 'sp4_r_v_b_4')
// (10, 1, 'sp4_h_r_14')
// (10, 1, 'sp4_v_t_40')
// (10, 1, 'sp4_v_t_44')
// (10, 2, 'local_g2_4')
// (10, 2, 'lutff_7/in_1')
// (10, 2, 'sp4_v_b_40')
// (10, 2, 'sp4_v_b_44')
// (10, 3, 'local_g3_5')
// (10, 3, 'lutff_5/in_3')
// (10, 3, 'sp4_v_b_29')
// (10, 3, 'sp4_v_b_33')
// (10, 4, 'sp4_v_b_16')
// (10, 4, 'sp4_v_b_20')
// (10, 5, 'sp4_h_r_13')
// (10, 5, 'sp4_h_r_28')
// (10, 5, 'sp4_h_r_7')
// (10, 5, 'sp4_v_b_5')
// (10, 5, 'sp4_v_b_9')
// (10, 5, 'sp4_v_t_44')
// (10, 6, 'sp4_v_b_44')
// (10, 7, 'sp4_v_b_33')
// (10, 8, 'sp4_v_b_20')
// (10, 9, 'sp4_h_l_42')
// (10, 9, 'sp4_h_r_29')
// (10, 9, 'sp4_h_r_4')
// (10, 9, 'sp4_v_b_9')
// (10, 10, 'sp4_h_r_12')
// (10, 12, 'sp4_h_r_12')
// (10, 13, 'sp4_h_r_10')
// (10, 13, 'sp4_h_r_7')
// (10, 13, 'sp4_v_t_36')
// (10, 13, 'sp4_v_t_41')
// (10, 14, 'sp4_h_r_15')
// (10, 14, 'sp4_v_b_36')
// (10, 14, 'sp4_v_b_41')
// (10, 15, 'sp4_v_b_25')
// (10, 15, 'sp4_v_b_28')
// (10, 16, 'sp4_v_b_12')
// (10, 16, 'sp4_v_b_17')
// (10, 17, 'sp4_v_b_1')
// (10, 17, 'sp4_v_b_4')
// (10, 17, 'sp4_v_t_36')
// (10, 17, 'sp4_v_t_41')
// (10, 18, 'local_g3_1')
// (10, 18, 'lutff_7/in_1')
// (10, 18, 'sp4_v_b_36')
// (10, 18, 'sp4_v_b_41')
// (10, 19, 'sp4_v_b_25')
// (10, 19, 'sp4_v_b_28')
// (10, 20, 'local_g0_1')
// (10, 20, 'lutff_6/in_1')
// (10, 20, 'sp4_v_b_12')
// (10, 20, 'sp4_v_b_17')
// (10, 21, 'sp4_v_b_1')
// (10, 21, 'sp4_v_b_4')
// (11, 1, 'sp4_h_r_27')
// (11, 2, 'local_g3_1')
// (11, 2, 'lutff_5/in_1')
// (11, 2, 'sp4_r_v_b_41')
// (11, 3, 'sp4_r_v_b_28')
// (11, 4, 'sp4_r_v_b_17')
// (11, 5, 'local_g3_0')
// (11, 5, 'lutff_3/in_0')
// (11, 5, 'sp4_h_r_18')
// (11, 5, 'sp4_h_r_24')
// (11, 5, 'sp4_h_r_41')
// (11, 5, 'sp4_r_v_b_4')
// (11, 9, 'sp4_h_r_17')
// (11, 9, 'sp4_h_r_40')
// (11, 10, 'sp4_h_r_25')
// (11, 12, 'sp4_h_r_25')
// (11, 13, 'sp4_h_r_18')
// (11, 13, 'sp4_h_r_23')
// (11, 14, 'sp4_h_r_26')
// (12, 1, 'sp4_h_r_38')
// (12, 1, 'sp4_v_t_41')
// (12, 2, 'sp4_v_b_41')
// (12, 3, 'sp4_v_b_28')
// (12, 4, 'sp4_v_b_17')
// (12, 5, 'local_g3_7')
// (12, 5, 'lutff_1/in_1')
// (12, 5, 'sp4_h_l_41')
// (12, 5, 'sp4_h_r_31')
// (12, 5, 'sp4_h_r_37')
// (12, 5, 'sp4_h_r_4')
// (12, 5, 'sp4_v_b_4')
// (12, 7, 'sp4_r_v_b_42')
// (12, 8, 'sp4_r_v_b_31')
// (12, 9, 'sp4_h_l_40')
// (12, 9, 'sp4_h_r_28')
// (12, 9, 'sp4_h_r_5')
// (12, 9, 'sp4_r_v_b_18')
// (12, 10, 'local_g1_7')
// (12, 10, 'lutff_4/in_2')
// (12, 10, 'sp4_h_r_36')
// (12, 10, 'sp4_r_v_b_7')
// (12, 12, 'sp4_h_r_36')
// (12, 13, 'sp4_h_r_31')
// (12, 13, 'sp4_h_r_34')
// (12, 14, 'sp4_h_r_39')
// (13, 1, 'sp4_h_l_38')
// (13, 1, 'sp4_h_r_7')
// (13, 2, 'sp4_h_r_11')
// (13, 2, 'sp4_r_v_b_44')
// (13, 3, 'sp4_r_v_b_33')
// (13, 4, 'sp4_r_v_b_20')
// (13, 5, 'sp4_h_l_37')
// (13, 5, 'sp4_h_r_17')
// (13, 5, 'sp4_h_r_4')
// (13, 5, 'sp4_h_r_42')
// (13, 5, 'sp4_r_v_b_9')
// (13, 6, 'local_g2_4')
// (13, 6, 'lutff_7/in_3')
// (13, 6, 'sp4_r_v_b_36')
// (13, 6, 'sp4_r_v_b_39')
// (13, 6, 'sp4_v_t_42')
// (13, 7, 'sp4_r_v_b_25')
// (13, 7, 'sp4_r_v_b_26')
// (13, 7, 'sp4_v_b_42')
// (13, 8, 'local_g2_7')
// (13, 8, 'lutff_0/in_3')
// (13, 8, 'sp4_r_v_b_12')
// (13, 8, 'sp4_r_v_b_15')
// (13, 8, 'sp4_v_b_31')
// (13, 9, 'sp4_h_r_16')
// (13, 9, 'sp4_h_r_41')
// (13, 9, 'sp4_r_v_b_1')
// (13, 9, 'sp4_r_v_b_2')
// (13, 9, 'sp4_v_b_18')
// (13, 10, 'sp4_h_l_36')
// (13, 10, 'sp4_h_r_2')
// (13, 10, 'sp4_h_r_5')
// (13, 10, 'sp4_v_b_7')
// (13, 12, 'sp4_h_l_36')
// (13, 12, 'sp4_h_r_1')
// (13, 13, 'sp4_h_r_42')
// (13, 13, 'sp4_h_r_47')
// (13, 14, 'sp4_h_l_39')
// (13, 14, 'sp4_h_r_2')
// (14, 1, 'sp4_h_r_18')
// (14, 1, 'sp4_v_t_44')
// (14, 2, 'sp4_h_r_22')
// (14, 2, 'sp4_v_b_44')
// (14, 3, 'local_g2_1')
// (14, 3, 'lutff_6/in_3')
// (14, 3, 'sp4_v_b_33')
// (14, 4, 'sp4_v_b_20')
// (14, 5, 'sp4_h_l_42')
// (14, 5, 'sp4_h_r_17')
// (14, 5, 'sp4_h_r_28')
// (14, 5, 'sp4_v_b_9')
// (14, 5, 'sp4_v_t_36')
// (14, 5, 'sp4_v_t_39')
// (14, 6, 'sp4_v_b_36')
// (14, 6, 'sp4_v_b_39')
// (14, 7, 'sp4_v_b_25')
// (14, 7, 'sp4_v_b_26')
// (14, 8, 'sp4_v_b_12')
// (14, 8, 'sp4_v_b_15')
// (14, 9, 'sp4_h_l_41')
// (14, 9, 'sp4_h_r_1')
// (14, 9, 'sp4_h_r_29')
// (14, 9, 'sp4_h_r_9')
// (14, 9, 'sp4_v_b_1')
// (14, 9, 'sp4_v_b_2')
// (14, 10, 'sp4_h_r_15')
// (14, 10, 'sp4_h_r_16')
// (14, 12, 'sp4_h_r_12')
// (14, 13, 'sp4_h_l_42')
// (14, 13, 'sp4_h_l_47')
// (14, 13, 'sp4_h_r_7')
// (14, 14, 'sp4_h_r_15')
// (15, 1, 'sp4_h_r_31')
// (15, 2, 'local_g2_3')
// (15, 2, 'lutff_0/in_1')
// (15, 2, 'sp4_h_r_35')
// (15, 2, 'sp4_r_v_b_40')
// (15, 3, 'local_g1_5')
// (15, 3, 'lutff_1/in_3')
// (15, 3, 'sp4_r_v_b_29')
// (15, 4, 'sp4_r_v_b_16')
// (15, 5, 'local_g3_4')
// (15, 5, 'lutff_0/in_1')
// (15, 5, 'sp4_h_r_28')
// (15, 5, 'sp4_h_r_41')
// (15, 5, 'sp4_r_v_b_5')
// (15, 6, 'sp4_r_v_b_40')
// (15, 7, 'sp4_r_v_b_29')
// (15, 8, 'sp4_r_v_b_16')
// (15, 9, 'sp4_h_r_12')
// (15, 9, 'sp4_h_r_20')
// (15, 9, 'sp4_h_r_40')
// (15, 9, 'sp4_r_v_b_5')
// (15, 10, 'sp4_h_r_26')
// (15, 10, 'sp4_h_r_29')
// (15, 12, 'sp4_h_r_25')
// (15, 13, 'sp4_h_r_18')
// (15, 14, 'sp4_h_r_26')
// (16, 1, 'sp4_h_r_42')
// (16, 1, 'sp4_v_t_40')
// (16, 2, 'sp4_h_r_46')
// (16, 2, 'sp4_v_b_40')
// (16, 3, 'sp4_v_b_29')
// (16, 4, 'sp4_v_b_16')
// (16, 5, 'sp4_h_l_41')
// (16, 5, 'sp4_h_r_41')
// (16, 5, 'sp4_h_r_8')
// (16, 5, 'sp4_v_b_5')
// (16, 5, 'sp4_v_t_40')
// (16, 6, 'sp4_v_b_40')
// (16, 7, 'sp4_v_b_29')
// (16, 8, 'sp4_v_b_16')
// (16, 9, 'sp4_h_l_40')
// (16, 9, 'sp4_h_r_25')
// (16, 9, 'sp4_h_r_33')
// (16, 9, 'sp4_h_r_5')
// (16, 9, 'sp4_v_b_5')
// (16, 10, 'sp4_h_r_39')
// (16, 10, 'sp4_h_r_40')
// (16, 11, 'sp4_r_v_b_39')
// (16, 12, 'sp4_h_r_36')
// (16, 12, 'sp4_r_v_b_26')
// (16, 13, 'sp4_h_r_31')
// (16, 13, 'sp4_r_v_b_15')
// (16, 14, 'sp4_h_r_39')
// (16, 14, 'sp4_r_v_b_2')
// (17, 1, 'sp4_h_l_42')
// (17, 1, 'sp4_h_r_4')
// (17, 2, 'sp4_h_l_46')
// (17, 2, 'sp4_h_r_11')
// (17, 5, 'sp4_h_l_41')
// (17, 5, 'sp4_h_r_21')
// (17, 5, 'sp4_h_r_4')
// (17, 9, 'sp4_h_r_16')
// (17, 9, 'sp4_h_r_36')
// (17, 9, 'sp4_h_r_44')
// (17, 10, 'sp4_h_l_39')
// (17, 10, 'sp4_h_l_40')
// (17, 10, 'sp4_h_r_2')
// (17, 10, 'sp4_r_v_b_42')
// (17, 10, 'sp4_v_t_39')
// (17, 11, 'sp4_r_v_b_31')
// (17, 11, 'sp4_v_b_39')
// (17, 12, 'sp4_h_l_36')
// (17, 12, 'sp4_h_r_1')
// (17, 12, 'sp4_r_v_b_18')
// (17, 12, 'sp4_v_b_26')
// (17, 13, 'sp4_h_r_42')
// (17, 13, 'sp4_r_v_b_7')
// (17, 13, 'sp4_v_b_15')
// (17, 14, 'sp4_h_l_39')
// (17, 14, 'sp4_v_b_2')
// (18, 1, 'sp4_h_r_17')
// (18, 2, 'sp4_h_r_22')
// (18, 5, 'sp4_h_r_17')
// (18, 5, 'sp4_h_r_32')
// (18, 9, 'sp4_h_l_36')
// (18, 9, 'sp4_h_l_44')
// (18, 9, 'sp4_h_r_1')
// (18, 9, 'sp4_h_r_29')
// (18, 9, 'sp4_v_t_42')
// (18, 10, 'sp4_h_r_15')
// (18, 10, 'sp4_v_b_42')
// (18, 11, 'sp4_v_b_31')
// (18, 12, 'sp4_h_r_12')
// (18, 12, 'sp4_v_b_18')
// (18, 13, 'sp4_h_l_42')
// (18, 13, 'sp4_v_b_7')
// (19, 1, 'sp4_h_r_28')
// (19, 2, 'sp4_h_r_35')
// (19, 5, 'sp4_h_r_28')
// (19, 5, 'sp4_h_r_45')
// (19, 6, 'sp4_r_v_b_39')
// (19, 7, 'sp4_r_v_b_26')
// (19, 8, 'sp4_r_v_b_15')
// (19, 9, 'sp4_h_r_12')
// (19, 9, 'sp4_h_r_40')
// (19, 9, 'sp4_r_v_b_2')
// (19, 10, 'sp4_h_r_26')
// (19, 12, 'sp4_h_r_25')
// (20, 1, 'sp4_h_r_41')
// (20, 2, 'sp4_h_r_46')
// (20, 2, 'sp4_r_v_b_41')
// (20, 3, 'sp4_r_v_b_28')
// (20, 3, 'sp4_r_v_b_40')
// (20, 4, 'sp4_r_v_b_17')
// (20, 4, 'sp4_r_v_b_29')
// (20, 5, 'sp4_h_l_45')
// (20, 5, 'sp4_h_r_41')
// (20, 5, 'sp4_r_v_b_16')
// (20, 5, 'sp4_r_v_b_4')
// (20, 5, 'sp4_v_t_39')
// (20, 6, 'sp4_r_v_b_41')
// (20, 6, 'sp4_r_v_b_5')
// (20, 6, 'sp4_v_b_39')
// (20, 7, 'sp4_r_v_b_28')
// (20, 7, 'sp4_r_v_b_44')
// (20, 7, 'sp4_v_b_26')
// (20, 8, 'neigh_op_tnr_2')
// (20, 8, 'sp4_r_v_b_17')
// (20, 8, 'sp4_r_v_b_33')
// (20, 8, 'sp4_v_b_15')
// (20, 9, 'neigh_op_rgt_2')
// (20, 9, 'sp4_h_l_40')
// (20, 9, 'sp4_h_r_25')
// (20, 9, 'sp4_h_r_9')
// (20, 9, 'sp4_r_v_b_20')
// (20, 9, 'sp4_r_v_b_36')
// (20, 9, 'sp4_r_v_b_4')
// (20, 9, 'sp4_v_b_2')
// (20, 10, 'neigh_op_bnr_2')
// (20, 10, 'sp4_h_r_39')
// (20, 10, 'sp4_r_v_b_25')
// (20, 10, 'sp4_r_v_b_9')
// (20, 11, 'sp4_r_v_b_12')
// (20, 12, 'sp4_h_r_36')
// (20, 12, 'sp4_r_v_b_1')
// (21, 1, 'sp4_h_l_41')
// (21, 1, 'sp4_v_t_41')
// (21, 2, 'sp4_h_l_46')
// (21, 2, 'sp4_v_b_41')
// (21, 2, 'sp4_v_t_40')
// (21, 3, 'sp4_v_b_28')
// (21, 3, 'sp4_v_b_40')
// (21, 4, 'sp4_v_b_17')
// (21, 4, 'sp4_v_b_29')
// (21, 5, 'sp4_h_l_41')
// (21, 5, 'sp4_v_b_16')
// (21, 5, 'sp4_v_b_4')
// (21, 5, 'sp4_v_t_41')
// (21, 6, 'sp4_v_b_41')
// (21, 6, 'sp4_v_b_5')
// (21, 6, 'sp4_v_t_44')
// (21, 7, 'sp4_v_b_28')
// (21, 7, 'sp4_v_b_44')
// (21, 8, 'neigh_op_top_2')
// (21, 8, 'sp4_v_b_17')
// (21, 8, 'sp4_v_b_33')
// (21, 8, 'sp4_v_t_36')
// (21, 9, 'lutff_2/out')
// (21, 9, 'sp4_h_r_20')
// (21, 9, 'sp4_h_r_36')
// (21, 9, 'sp4_v_b_20')
// (21, 9, 'sp4_v_b_36')
// (21, 9, 'sp4_v_b_4')
// (21, 10, 'neigh_op_bot_2')
// (21, 10, 'sp4_h_l_39')
// (21, 10, 'sp4_v_b_25')
// (21, 10, 'sp4_v_b_9')
// (21, 11, 'sp4_v_b_12')
// (21, 12, 'sp4_h_l_36')
// (21, 12, 'sp4_v_b_1')
// (22, 8, 'neigh_op_tnl_2')
// (22, 9, 'neigh_op_lft_2')
// (22, 9, 'sp4_h_l_36')
// (22, 9, 'sp4_h_r_33')
// (22, 10, 'neigh_op_bnl_2')
// (23, 9, 'sp4_h_r_44')
// (24, 9, 'sp4_h_l_44')

reg n176 = 0;
// (1, 1, 'sp4_r_v_b_17')
// (1, 2, 'sp4_r_v_b_4')
// (1, 3, 'sp4_r_v_b_41')
// (1, 4, 'sp4_r_v_b_28')
// (1, 4, 'sp4_r_v_b_44')
// (1, 5, 'neigh_op_tnr_2')
// (1, 5, 'sp4_r_v_b_17')
// (1, 5, 'sp4_r_v_b_33')
// (1, 6, 'neigh_op_rgt_2')
// (1, 6, 'sp4_h_r_9')
// (1, 6, 'sp4_r_v_b_20')
// (1, 6, 'sp4_r_v_b_4')
// (1, 7, 'neigh_op_bnr_2')
// (1, 7, 'sp4_r_v_b_9')
// (2, 0, 'span4_vert_17')
// (2, 1, 'local_g1_1')
// (2, 1, 'lutff_4/in_2')
// (2, 1, 'sp4_v_b_17')
// (2, 2, 'local_g1_1')
// (2, 2, 'lutff_0/in_2')
// (2, 2, 'lutff_2/in_0')
// (2, 2, 'sp4_h_r_9')
// (2, 2, 'sp4_v_b_4')
// (2, 2, 'sp4_v_t_41')
// (2, 3, 'sp4_h_r_2')
// (2, 3, 'sp4_r_v_b_40')
// (2, 3, 'sp4_v_b_41')
// (2, 3, 'sp4_v_t_44')
// (2, 4, 'sp4_r_v_b_29')
// (2, 4, 'sp4_r_v_b_45')
// (2, 4, 'sp4_v_b_28')
// (2, 4, 'sp4_v_b_44')
// (2, 5, 'local_g0_2')
// (2, 5, 'lutff_4/in_2')
// (2, 5, 'neigh_op_top_2')
// (2, 5, 'sp4_r_v_b_16')
// (2, 5, 'sp4_r_v_b_32')
// (2, 5, 'sp4_v_b_17')
// (2, 5, 'sp4_v_b_33')
// (2, 6, 'local_g2_2')
// (2, 6, 'lutff_2/in_2')
// (2, 6, 'lutff_2/out')
// (2, 6, 'lutff_7/in_1')
// (2, 6, 'sp4_h_r_20')
// (2, 6, 'sp4_h_r_4')
// (2, 6, 'sp4_r_v_b_21')
// (2, 6, 'sp4_r_v_b_5')
// (2, 6, 'sp4_v_b_20')
// (2, 6, 'sp4_v_b_4')
// (2, 7, 'local_g1_2')
// (2, 7, 'lutff_1/in_0')
// (2, 7, 'neigh_op_bot_2')
// (2, 7, 'sp4_r_v_b_8')
// (2, 7, 'sp4_v_b_9')
// (3, 2, 'sp4_h_r_10')
// (3, 2, 'sp4_h_r_20')
// (3, 2, 'sp4_v_t_40')
// (3, 3, 'sp4_h_r_1')
// (3, 3, 'sp4_h_r_15')
// (3, 3, 'sp4_v_b_40')
// (3, 3, 'sp4_v_t_45')
// (3, 4, 'local_g3_5')
// (3, 4, 'lutff_4/in_0')
// (3, 4, 'sp4_v_b_29')
// (3, 4, 'sp4_v_b_45')
// (3, 5, 'local_g3_2')
// (3, 5, 'lutff_4/in_1')
// (3, 5, 'neigh_op_tnl_2')
// (3, 5, 'sp4_v_b_16')
// (3, 5, 'sp4_v_b_32')
// (3, 6, 'local_g0_1')
// (3, 6, 'lutff_5/in_0')
// (3, 6, 'neigh_op_lft_2')
// (3, 6, 'sp4_h_r_17')
// (3, 6, 'sp4_h_r_33')
// (3, 6, 'sp4_v_b_21')
// (3, 6, 'sp4_v_b_5')
// (3, 7, 'neigh_op_bnl_2')
// (3, 7, 'sp4_h_r_8')
// (3, 7, 'sp4_v_b_8')
// (4, 1, 'local_g2_5')
// (4, 1, 'lutff_7/in_2')
// (4, 1, 'sp4_r_v_b_13')
// (4, 2, 'local_g0_7')
// (4, 2, 'lutff_1/in_0')
// (4, 2, 'sp4_h_r_23')
// (4, 2, 'sp4_h_r_33')
// (4, 2, 'sp4_r_v_b_0')
// (4, 3, 'local_g2_2')
// (4, 3, 'local_g3_2')
// (4, 3, 'lutff_0/in_3')
// (4, 3, 'lutff_2/in_3')
// (4, 3, 'lutff_3/in_3')
// (4, 3, 'sp4_h_r_12')
// (4, 3, 'sp4_h_r_26')
// (4, 3, 'sp4_r_v_b_44')
// (4, 4, 'local_g0_2')
// (4, 4, 'lutff_2/in_0')
// (4, 4, 'sp4_r_v_b_33')
// (4, 5, 'local_g3_4')
// (4, 5, 'lutff_2/in_1')
// (4, 5, 'sp4_r_v_b_20')
// (4, 6, 'sp4_h_r_28')
// (4, 6, 'sp4_h_r_44')
// (4, 6, 'sp4_r_v_b_9')
// (4, 7, 'local_g1_5')
// (4, 7, 'lutff_4/in_0')
// (4, 7, 'sp4_h_r_21')
// (5, 0, 'span4_vert_13')
// (5, 1, 'local_g3_4')
// (5, 1, 'lutff_2/in_1')
// (5, 1, 'sp4_r_v_b_20')
// (5, 1, 'sp4_v_b_13')
// (5, 2, 'sp4_h_r_34')
// (5, 2, 'sp4_h_r_44')
// (5, 2, 'sp4_r_v_b_9')
// (5, 2, 'sp4_v_b_0')
// (5, 2, 'sp4_v_t_44')
// (5, 3, 'sp4_h_r_25')
// (5, 3, 'sp4_h_r_39')
// (5, 3, 'sp4_v_b_44')
// (5, 4, 'local_g3_1')
// (5, 4, 'lutff_0/in_0')
// (5, 4, 'sp4_v_b_33')
// (5, 5, 'sp4_v_b_20')
// (5, 6, 'local_g3_1')
// (5, 6, 'lutff_7/in_3')
// (5, 6, 'sp4_h_l_44')
// (5, 6, 'sp4_h_r_41')
// (5, 6, 'sp4_v_b_9')
// (5, 7, 'local_g2_0')
// (5, 7, 'lutff_2/in_2')
// (5, 7, 'sp4_h_r_32')
// (6, 0, 'span4_vert_20')
// (6, 1, 'sp4_v_b_20')
// (6, 2, 'sp4_h_l_44')
// (6, 2, 'sp4_h_r_0')
// (6, 2, 'sp4_h_r_47')
// (6, 2, 'sp4_h_r_9')
// (6, 2, 'sp4_v_b_9')
// (6, 3, 'sp4_h_l_39')
// (6, 3, 'sp4_h_r_2')
// (6, 3, 'sp4_h_r_36')
// (6, 6, 'sp4_h_l_41')
// (6, 7, 'sp4_h_r_45')
// (7, 2, 'local_g0_5')
// (7, 2, 'lutff_0/in_1')
// (7, 2, 'sp4_h_l_47')
// (7, 2, 'sp4_h_r_10')
// (7, 2, 'sp4_h_r_13')
// (7, 2, 'sp4_h_r_20')
// (7, 3, 'sp4_h_l_36')
// (7, 3, 'sp4_h_r_15')
// (7, 3, 'sp4_h_r_4')
// (7, 7, 'sp4_h_l_45')
// (8, 2, 'local_g0_7')
// (8, 2, 'lutff_2/in_1')
// (8, 2, 'lutff_3/in_0')
// (8, 2, 'sp4_h_r_23')
// (8, 2, 'sp4_h_r_24')
// (8, 2, 'sp4_h_r_33')
// (8, 3, 'local_g0_1')
// (8, 3, 'local_g1_1')
// (8, 3, 'lutff_0/in_1')
// (8, 3, 'lutff_1/in_1')
// (8, 3, 'sp4_h_r_17')
// (8, 3, 'sp4_h_r_26')
// (9, 1, 'local_g2_6')
// (9, 1, 'lutff_1/in_1')
// (9, 1, 'lutff_6/in_2')
// (9, 1, 'sp4_r_v_b_14')
// (9, 2, 'local_g2_5')
// (9, 2, 'lutff_1/in_2')
// (9, 2, 'lutff_2/in_3')
// (9, 2, 'lutff_7/in_2')
// (9, 2, 'sp4_h_r_34')
// (9, 2, 'sp4_h_r_37')
// (9, 2, 'sp4_h_r_44')
// (9, 2, 'sp4_r_v_b_3')
// (9, 3, 'local_g3_7')
// (9, 3, 'lutff_1/in_3')
// (9, 3, 'sp4_h_r_28')
// (9, 3, 'sp4_h_r_39')
// (10, 0, 'span4_vert_14')
// (10, 1, 'sp4_v_b_14')
// (10, 2, 'sp4_h_l_37')
// (10, 2, 'sp4_h_l_44')
// (10, 2, 'sp4_h_r_47')
// (10, 2, 'sp4_v_b_3')
// (10, 3, 'sp4_h_l_39')
// (10, 3, 'sp4_h_r_41')
// (11, 2, 'sp4_h_l_47')
// (11, 3, 'sp4_h_l_41')

reg n177 = 0;
// (1, 1, 'sp4_r_v_b_25')
// (1, 2, 'sp4_r_v_b_12')
// (1, 3, 'sp4_r_v_b_1')
// (2, 0, 'span4_vert_25')
// (2, 1, 'sp4_v_b_25')
// (2, 2, 'local_g1_4')
// (2, 2, 'lutff_4/in_3')
// (2, 2, 'sp4_v_b_12')
// (2, 3, 'sp4_h_r_1')
// (2, 3, 'sp4_v_b_1')
// (3, 1, 'sp4_r_v_b_32')
// (3, 2, 'local_g3_5')
// (3, 2, 'lutff_3/in_3')
// (3, 2, 'sp4_r_v_b_21')
// (3, 3, 'sp4_h_r_12')
// (3, 3, 'sp4_r_v_b_8')
// (3, 4, 'sp4_r_v_b_39')
// (3, 5, 'sp4_r_v_b_26')
// (3, 6, 'local_g2_7')
// (3, 6, 'lutff_3/in_0')
// (3, 6, 'sp4_r_v_b_15')
// (3, 7, 'sp4_r_v_b_2')
// (3, 8, 'sp4_r_v_b_42')
// (3, 9, 'sp4_r_v_b_31')
// (3, 10, 'sp4_r_v_b_18')
// (3, 11, 'sp4_r_v_b_7')
// (3, 15, 'sp12_h_r_1')
// (3, 15, 'sp12_v_t_22')
// (3, 16, 'sp12_v_b_22')
// (3, 17, 'sp12_v_b_21')
// (3, 18, 'sp12_v_b_18')
// (3, 19, 'sp12_v_b_17')
// (3, 20, 'local_g2_6')
// (3, 20, 'lutff_5/in_1')
// (3, 20, 'sp12_v_b_14')
// (3, 21, 'sp12_v_b_13')
// (3, 22, 'sp12_v_b_10')
// (3, 23, 'sp12_v_b_9')
// (3, 24, 'sp12_v_b_6')
// (3, 25, 'sp12_v_b_5')
// (3, 26, 'sp12_v_b_2')
// (3, 27, 'sp12_v_b_1')
// (4, 0, 'span4_vert_32')
// (4, 1, 'sp4_v_b_32')
// (4, 2, 'sp4_v_b_21')
// (4, 3, 'sp4_h_r_25')
// (4, 3, 'sp4_h_r_8')
// (4, 3, 'sp4_v_b_8')
// (4, 3, 'sp4_v_t_39')
// (4, 4, 'sp4_v_b_39')
// (4, 5, 'sp4_h_r_10')
// (4, 5, 'sp4_v_b_26')
// (4, 6, 'sp4_v_b_15')
// (4, 7, 'local_g1_0')
// (4, 7, 'lutff_2/in_1')
// (4, 7, 'sp4_h_r_0')
// (4, 7, 'sp4_h_r_7')
// (4, 7, 'sp4_v_b_2')
// (4, 7, 'sp4_v_t_42')
// (4, 8, 'sp4_v_b_42')
// (4, 9, 'sp4_v_b_31')
// (4, 10, 'local_g0_2')
// (4, 10, 'lutff_5/in_1')
// (4, 10, 'sp4_v_b_18')
// (4, 11, 'sp4_v_b_7')
// (4, 15, 'sp12_h_r_2')
// (5, 1, 'local_g1_1')
// (5, 1, 'lutff_1/in_1')
// (5, 1, 'sp4_r_v_b_25')
// (5, 2, 'local_g2_4')
// (5, 2, 'lutff_4/in_2')
// (5, 2, 'sp4_r_v_b_12')
// (5, 3, 'local_g1_1')
// (5, 3, 'lutff_3/in_1')
// (5, 3, 'sp4_h_r_21')
// (5, 3, 'sp4_h_r_36')
// (5, 3, 'sp4_r_v_b_1')
// (5, 5, 'local_g0_7')
// (5, 5, 'lutff_4/in_3')
// (5, 5, 'sp4_h_r_23')
// (5, 7, 'sp4_h_r_13')
// (5, 7, 'sp4_h_r_18')
// (5, 15, 'sp12_h_r_5')
// (6, 0, 'span4_vert_25')
// (6, 1, 'sp4_v_b_25')
// (6, 2, 'sp4_v_b_12')
// (6, 3, 'sp4_h_l_36')
// (6, 3, 'sp4_h_r_1')
// (6, 3, 'sp4_h_r_32')
// (6, 3, 'sp4_v_b_1')
// (6, 5, 'sp4_h_r_34')
// (6, 7, 'sp4_h_r_24')
// (6, 7, 'sp4_h_r_31')
// (6, 15, 'sp12_h_r_6')
// (7, 3, 'sp4_h_r_12')
// (7, 3, 'sp4_h_r_45')
// (7, 4, 'sp4_r_v_b_42')
// (7, 5, 'sp4_h_r_47')
// (7, 5, 'sp4_r_v_b_31')
// (7, 6, 'sp4_r_v_b_18')
// (7, 7, 'sp4_h_r_37')
// (7, 7, 'sp4_h_r_42')
// (7, 7, 'sp4_r_v_b_7')
// (7, 15, 'sp12_h_r_9')
// (7, 18, 'sp4_r_v_b_40')
// (7, 19, 'sp4_r_v_b_29')
// (7, 20, 'sp4_r_v_b_16')
// (7, 21, 'local_g1_5')
// (7, 21, 'lutff_3/in_3')
// (7, 21, 'sp4_r_v_b_5')
// (8, 3, 'sp4_h_l_45')
// (8, 3, 'sp4_h_r_1')
// (8, 3, 'sp4_h_r_25')
// (8, 3, 'sp4_h_r_8')
// (8, 3, 'sp4_v_t_42')
// (8, 4, 'local_g1_6')
// (8, 4, 'lutff_4/in_3')
// (8, 4, 'sp4_h_r_6')
// (8, 4, 'sp4_v_b_42')
// (8, 5, 'sp4_h_l_47')
// (8, 5, 'sp4_h_r_2')
// (8, 5, 'sp4_v_b_31')
// (8, 6, 'sp4_v_b_18')
// (8, 7, 'sp4_h_l_37')
// (8, 7, 'sp4_h_l_42')
// (8, 7, 'sp4_v_b_7')
// (8, 12, 'local_g0_1')
// (8, 12, 'lutff_7/in_2')
// (8, 12, 'sp12_h_r_1')
// (8, 12, 'sp12_v_t_22')
// (8, 13, 'sp12_v_b_22')
// (8, 14, 'sp12_v_b_21')
// (8, 15, 'sp12_h_r_10')
// (8, 15, 'sp12_v_b_18')
// (8, 16, 'sp12_v_b_17')
// (8, 17, 'sp12_v_b_14')
// (8, 17, 'sp4_v_t_40')
// (8, 18, 'sp12_v_b_13')
// (8, 18, 'sp4_v_b_40')
// (8, 19, 'sp12_v_b_10')
// (8, 19, 'sp4_v_b_29')
// (8, 20, 'sp12_v_b_9')
// (8, 20, 'sp4_v_b_16')
// (8, 21, 'sp12_v_b_6')
// (8, 21, 'sp4_v_b_5')
// (8, 22, 'sp12_v_b_5')
// (8, 23, 'sp12_v_b_2')
// (8, 24, 'sp12_v_b_1')
// (9, 1, 'local_g0_3')
// (9, 1, 'lutff_7/in_0')
// (9, 1, 'sp4_r_v_b_27')
// (9, 2, 'sp4_r_v_b_14')
// (9, 3, 'sp4_h_r_12')
// (9, 3, 'sp4_h_r_21')
// (9, 3, 'sp4_h_r_36')
// (9, 3, 'sp4_r_v_b_3')
// (9, 4, 'local_g0_3')
// (9, 4, 'lutff_4/in_3')
// (9, 4, 'sp4_h_r_19')
// (9, 4, 'sp4_r_v_b_47')
// (9, 5, 'sp4_h_r_15')
// (9, 5, 'sp4_r_v_b_34')
// (9, 6, 'sp4_r_v_b_23')
// (9, 7, 'local_g2_2')
// (9, 7, 'lutff_6/in_0')
// (9, 7, 'sp4_r_v_b_10')
// (9, 8, 'sp4_r_v_b_38')
// (9, 9, 'sp4_r_v_b_27')
// (9, 10, 'sp4_r_v_b_14')
// (9, 11, 'sp4_r_v_b_3')
// (9, 12, 'sp12_h_r_2')
// (9, 12, 'sp4_r_v_b_38')
// (9, 13, 'sp4_r_v_b_27')
// (9, 14, 'local_g2_6')
// (9, 14, 'lutff_4/in_2')
// (9, 14, 'sp4_r_v_b_14')
// (9, 15, 'sp12_h_r_13')
// (9, 15, 'sp4_r_v_b_3')
// (9, 16, 'sp4_r_v_b_43')
// (9, 17, 'sp4_r_v_b_30')
// (9, 18, 'sp4_r_v_b_19')
// (9, 19, 'sp4_r_v_b_6')
// (10, 0, 'span4_vert_27')
// (10, 1, 'local_g3_3')
// (10, 1, 'lutff_1/in_1')
// (10, 1, 'sp4_v_b_27')
// (10, 2, 'sp4_v_b_14')
// (10, 3, 'sp4_h_l_36')
// (10, 3, 'sp4_h_r_10')
// (10, 3, 'sp4_h_r_25')
// (10, 3, 'sp4_h_r_32')
// (10, 3, 'sp4_v_b_3')
// (10, 3, 'sp4_v_t_47')
// (10, 4, 'local_g2_6')
// (10, 4, 'lutff_7/in_1')
// (10, 4, 'sp4_h_r_30')
// (10, 4, 'sp4_v_b_47')
// (10, 5, 'sp4_h_r_26')
// (10, 5, 'sp4_v_b_34')
// (10, 6, 'sp4_v_b_23')
// (10, 7, 'sp4_h_r_9')
// (10, 7, 'sp4_v_b_10')
// (10, 7, 'sp4_v_t_38')
// (10, 8, 'sp4_v_b_38')
// (10, 9, 'sp4_v_b_27')
// (10, 10, 'sp4_v_b_14')
// (10, 11, 'sp4_v_b_3')
// (10, 11, 'sp4_v_t_38')
// (10, 12, 'sp12_h_r_5')
// (10, 12, 'sp4_v_b_38')
// (10, 13, 'sp4_v_b_27')
// (10, 14, 'sp4_v_b_14')
// (10, 15, 'sp12_h_r_14')
// (10, 15, 'sp4_v_b_3')
// (10, 15, 'sp4_v_t_43')
// (10, 16, 'sp4_v_b_43')
// (10, 17, 'sp4_r_v_b_37')
// (10, 17, 'sp4_v_b_30')
// (10, 18, 'local_g0_3')
// (10, 18, 'lutff_6/in_1')
// (10, 18, 'sp4_r_v_b_24')
// (10, 18, 'sp4_v_b_19')
// (10, 19, 'sp4_r_v_b_13')
// (10, 19, 'sp4_v_b_6')
// (10, 20, 'local_g1_0')
// (10, 20, 'lutff_6/in_3')
// (10, 20, 'sp4_r_v_b_0')
// (11, 3, 'sp4_h_r_23')
// (11, 3, 'sp4_h_r_36')
// (11, 3, 'sp4_h_r_45')
// (11, 4, 'sp4_h_r_43')
// (11, 5, 'sp4_h_r_39')
// (11, 7, 'sp4_h_r_20')
// (11, 8, 'sp4_r_v_b_41')
// (11, 9, 'sp4_r_v_b_28')
// (11, 10, 'sp4_r_v_b_17')
// (11, 11, 'sp4_r_v_b_4')
// (11, 12, 'sp12_h_r_6')
// (11, 15, 'sp12_h_r_17')
// (11, 16, 'sp4_h_r_6')
// (11, 16, 'sp4_v_t_37')
// (11, 17, 'sp4_v_b_37')
// (11, 18, 'sp4_v_b_24')
// (11, 19, 'sp4_v_b_13')
// (11, 20, 'sp4_v_b_0')
// (12, 3, 'sp4_h_l_36')
// (12, 3, 'sp4_h_l_45')
// (12, 3, 'sp4_h_r_10')
// (12, 3, 'sp4_h_r_34')
// (12, 3, 'sp4_h_r_8')
// (12, 4, 'sp4_h_l_43')
// (12, 4, 'sp4_h_r_10')
// (12, 5, 'local_g1_6')
// (12, 5, 'lutff_0/in_3')
// (12, 5, 'sp4_h_l_39')
// (12, 5, 'sp4_h_r_6')
// (12, 7, 'sp4_h_r_33')
// (12, 7, 'sp4_h_r_4')
// (12, 7, 'sp4_v_t_41')
// (12, 8, 'sp4_v_b_41')
// (12, 9, 'sp4_v_b_28')
// (12, 10, 'local_g1_1')
// (12, 10, 'lutff_0/in_0')
// (12, 10, 'sp4_v_b_17')
// (12, 11, 'sp4_v_b_4')
// (12, 12, 'sp12_h_r_9')
// (12, 15, 'sp12_h_r_18')
// (12, 16, 'sp4_h_r_19')
// (13, 3, 'sp4_h_r_21')
// (13, 3, 'sp4_h_r_23')
// (13, 3, 'sp4_h_r_47')
// (13, 4, 'sp4_h_r_23')
// (13, 4, 'sp4_r_v_b_41')
// (13, 5, 'local_g1_3')
// (13, 5, 'lutff_1/in_1')
// (13, 5, 'sp4_h_r_19')
// (13, 5, 'sp4_r_v_b_28')
// (13, 6, 'sp4_r_v_b_17')
// (13, 7, 'sp4_h_r_17')
// (13, 7, 'sp4_h_r_44')
// (13, 7, 'sp4_r_v_b_4')
// (13, 12, 'sp12_h_r_10')
// (13, 15, 'sp12_h_r_21')
// (13, 16, 'sp4_h_r_30')
// (14, 3, 'local_g1_1')
// (14, 3, 'lutff_2/in_0')
// (14, 3, 'sp4_h_l_47')
// (14, 3, 'sp4_h_r_1')
// (14, 3, 'sp4_h_r_10')
// (14, 3, 'sp4_h_r_32')
// (14, 3, 'sp4_h_r_34')
// (14, 3, 'sp4_v_t_41')
// (14, 4, 'sp4_h_r_34')
// (14, 4, 'sp4_v_b_41')
// (14, 5, 'sp4_h_r_30')
// (14, 5, 'sp4_v_b_28')
// (14, 6, 'sp4_v_b_17')
// (14, 7, 'sp4_h_l_44')
// (14, 7, 'sp4_h_r_28')
// (14, 7, 'sp4_v_b_4')
// (14, 12, 'sp12_h_r_13')
// (14, 13, 'sp4_r_v_b_36')
// (14, 14, 'sp4_r_v_b_25')
// (14, 15, 'sp12_h_r_22')
// (14, 15, 'sp4_r_v_b_12')
// (14, 16, 'sp4_h_r_43')
// (14, 16, 'sp4_r_v_b_1')
// (15, 1, 'sp4_r_v_b_29')
// (15, 1, 'sp4_r_v_b_37')
// (15, 2, 'sp4_r_v_b_16')
// (15, 2, 'sp4_r_v_b_24')
// (15, 3, 'sp12_h_r_1')
// (15, 3, 'sp12_v_t_22')
// (15, 3, 'sp4_h_r_12')
// (15, 3, 'sp4_h_r_23')
// (15, 3, 'sp4_h_r_45')
// (15, 3, 'sp4_h_r_47')
// (15, 3, 'sp4_r_v_b_13')
// (15, 3, 'sp4_r_v_b_5')
// (15, 4, 'local_g1_0')
// (15, 4, 'lutff_1/in_0')
// (15, 4, 'sp12_v_b_22')
// (15, 4, 'sp4_h_r_47')
// (15, 4, 'sp4_r_v_b_0')
// (15, 4, 'sp4_r_v_b_46')
// (15, 5, 'local_g2_3')
// (15, 5, 'lutff_4/in_3')
// (15, 5, 'sp12_v_b_21')
// (15, 5, 'sp4_h_r_43')
// (15, 5, 'sp4_r_v_b_35')
// (15, 6, 'sp12_v_b_18')
// (15, 6, 'sp4_r_v_b_22')
// (15, 7, 'sp12_v_b_17')
// (15, 7, 'sp4_h_r_41')
// (15, 7, 'sp4_r_v_b_11')
// (15, 8, 'sp12_v_b_14')
// (15, 9, 'sp12_v_b_13')
// (15, 10, 'sp12_v_b_10')
// (15, 11, 'sp12_v_b_9')
// (15, 12, 'sp12_h_r_14')
// (15, 12, 'sp12_v_b_6')
// (15, 12, 'sp4_v_t_36')
// (15, 13, 'sp12_v_b_5')
// (15, 13, 'sp4_v_b_36')
// (15, 14, 'sp12_v_b_2')
// (15, 14, 'sp4_v_b_25')
// (15, 15, 'sp12_h_l_22')
// (15, 15, 'sp12_v_b_1')
// (15, 15, 'sp4_v_b_12')
// (15, 16, 'sp4_h_l_43')
// (15, 16, 'sp4_v_b_1')
// (16, 0, 'span4_vert_29')
// (16, 0, 'span4_vert_37')
// (16, 1, 'sp4_v_b_29')
// (16, 1, 'sp4_v_b_37')
// (16, 2, 'local_g1_0')
// (16, 2, 'lutff_1/in_0')
// (16, 2, 'sp4_v_b_16')
// (16, 2, 'sp4_v_b_24')
// (16, 3, 'sp12_h_r_2')
// (16, 3, 'sp4_h_l_45')
// (16, 3, 'sp4_h_l_47')
// (16, 3, 'sp4_h_r_10')
// (16, 3, 'sp4_h_r_25')
// (16, 3, 'sp4_h_r_34')
// (16, 3, 'sp4_h_r_5')
// (16, 3, 'sp4_v_b_13')
// (16, 3, 'sp4_v_b_5')
// (16, 3, 'sp4_v_t_46')
// (16, 4, 'sp4_h_l_47')
// (16, 4, 'sp4_h_r_7')
// (16, 4, 'sp4_v_b_0')
// (16, 4, 'sp4_v_b_46')
// (16, 5, 'sp4_h_l_43')
// (16, 5, 'sp4_h_r_3')
// (16, 5, 'sp4_v_b_35')
// (16, 6, 'local_g1_6')
// (16, 6, 'lutff_5/in_2')
// (16, 6, 'sp4_v_b_22')
// (16, 7, 'sp4_h_l_41')
// (16, 7, 'sp4_v_b_11')
// (16, 12, 'sp12_h_r_17')
// (17, 3, 'sp12_h_r_5')
// (17, 3, 'sp4_h_r_16')
// (17, 3, 'sp4_h_r_23')
// (17, 3, 'sp4_h_r_36')
// (17, 3, 'sp4_h_r_47')
// (17, 4, 'sp4_h_r_18')
// (17, 5, 'sp4_h_r_14')
// (17, 12, 'sp12_h_r_18')
// (18, 3, 'sp12_h_r_6')
// (18, 3, 'sp4_h_l_36')
// (18, 3, 'sp4_h_l_47')
// (18, 3, 'sp4_h_r_10')
// (18, 3, 'sp4_h_r_29')
// (18, 3, 'sp4_h_r_34')
// (18, 4, 'sp4_h_r_31')
// (18, 5, 'sp4_h_r_27')
// (18, 12, 'sp12_h_r_21')
// (19, 1, 'sp4_r_v_b_42')
// (19, 2, 'neigh_op_tnr_1')
// (19, 2, 'sp4_r_v_b_31')
// (19, 2, 'sp4_r_v_b_47')
// (19, 3, 'neigh_op_rgt_1')
// (19, 3, 'sp12_h_r_9')
// (19, 3, 'sp4_h_r_23')
// (19, 3, 'sp4_h_r_40')
// (19, 3, 'sp4_h_r_47')
// (19, 3, 'sp4_r_v_b_18')
// (19, 3, 'sp4_r_v_b_34')
// (19, 4, 'neigh_op_bnr_1')
// (19, 4, 'sp4_h_r_42')
// (19, 4, 'sp4_r_v_b_23')
// (19, 4, 'sp4_r_v_b_7')
// (19, 5, 'sp4_h_r_38')
// (19, 5, 'sp4_r_v_b_10')
// (19, 12, 'sp12_h_r_22')
// (20, 0, 'span12_vert_22')
// (20, 0, 'span4_vert_42')
// (20, 1, 'sp12_v_b_22')
// (20, 1, 'sp4_v_b_42')
// (20, 1, 'sp4_v_t_47')
// (20, 2, 'neigh_op_top_1')
// (20, 2, 'sp12_v_b_21')
// (20, 2, 'sp4_v_b_31')
// (20, 2, 'sp4_v_b_47')
// (20, 3, 'lutff_1/out')
// (20, 3, 'sp12_h_r_10')
// (20, 3, 'sp12_v_b_18')
// (20, 3, 'sp4_h_l_40')
// (20, 3, 'sp4_h_l_47')
// (20, 3, 'sp4_h_r_2')
// (20, 3, 'sp4_h_r_34')
// (20, 3, 'sp4_v_b_18')
// (20, 3, 'sp4_v_b_34')
// (20, 4, 'neigh_op_bot_1')
// (20, 4, 'sp12_v_b_17')
// (20, 4, 'sp4_h_l_42')
// (20, 4, 'sp4_v_b_23')
// (20, 4, 'sp4_v_b_7')
// (20, 5, 'sp12_v_b_14')
// (20, 5, 'sp4_h_l_38')
// (20, 5, 'sp4_v_b_10')
// (20, 6, 'sp12_v_b_13')
// (20, 7, 'sp12_v_b_10')
// (20, 8, 'sp12_v_b_9')
// (20, 9, 'sp12_v_b_6')
// (20, 10, 'sp12_v_b_5')
// (20, 11, 'sp12_v_b_2')
// (20, 12, 'sp12_h_l_22')
// (20, 12, 'sp12_v_b_1')
// (21, 2, 'neigh_op_tnl_1')
// (21, 3, 'neigh_op_lft_1')
// (21, 3, 'sp12_h_r_13')
// (21, 3, 'sp4_h_r_15')
// (21, 3, 'sp4_h_r_47')
// (21, 4, 'neigh_op_bnl_1')
// (22, 3, 'sp12_h_r_14')
// (22, 3, 'sp4_h_l_47')
// (22, 3, 'sp4_h_r_26')
// (23, 3, 'sp12_h_r_17')
// (23, 3, 'sp4_h_r_39')
// (24, 3, 'sp12_h_r_18')
// (24, 3, 'sp4_h_l_39')
// (25, 3, 'sp12_h_r_21')

wire n178;
// (1, 1, 'sp4_r_v_b_31')
// (1, 1, 'sp4_r_v_b_35')
// (1, 2, 'sp4_r_v_b_18')
// (1, 2, 'sp4_r_v_b_22')
// (1, 3, 'sp4_r_v_b_11')
// (1, 3, 'sp4_r_v_b_7')
// (2, 0, 'span4_vert_31')
// (2, 0, 'span4_vert_35')
// (2, 1, 'local_g3_3')
// (2, 1, 'lutff_global/cen')
// (2, 1, 'sp4_v_b_31')
// (2, 1, 'sp4_v_b_35')
// (2, 2, 'local_g0_2')
// (2, 2, 'lutff_global/cen')
// (2, 2, 'sp4_v_b_18')
// (2, 2, 'sp4_v_b_22')
// (2, 3, 'sp4_h_r_11')
// (2, 3, 'sp4_h_r_7')
// (2, 3, 'sp4_v_b_11')
// (2, 3, 'sp4_v_b_7')
// (3, 3, 'sp4_h_r_18')
// (3, 3, 'sp4_h_r_22')
// (4, 3, 'sp4_h_r_31')
// (4, 3, 'sp4_h_r_35')
// (5, 3, 'sp4_h_r_42')
// (5, 3, 'sp4_h_r_46')
// (6, 2, 'neigh_op_tnr_3')
// (6, 3, 'neigh_op_rgt_3')
// (6, 3, 'sp4_h_l_42')
// (6, 3, 'sp4_h_l_46')
// (6, 3, 'sp4_h_r_11')
// (6, 4, 'neigh_op_bnr_3')
// (7, 2, 'neigh_op_top_3')
// (7, 3, 'lutff_3/out')
// (7, 3, 'sp4_h_r_22')
// (7, 4, 'neigh_op_bot_3')
// (8, 2, 'neigh_op_tnl_3')
// (8, 3, 'neigh_op_lft_3')
// (8, 3, 'sp4_h_r_35')
// (8, 4, 'neigh_op_bnl_3')
// (9, 3, 'sp4_h_r_46')
// (10, 3, 'sp4_h_l_46')

reg n179 = 0;
// (1, 1, 'sp4_r_v_b_32')
// (1, 2, 'sp4_r_v_b_21')
// (1, 3, 'sp4_r_v_b_8')
// (2, 0, 'span4_vert_32')
// (2, 1, 'local_g2_0')
// (2, 1, 'lutff_2/in_0')
// (2, 1, 'sp4_v_b_32')
// (2, 2, 'sp4_v_b_21')
// (2, 3, 'sp4_h_r_8')
// (2, 3, 'sp4_v_b_8')
// (2, 7, 'sp4_h_r_4')
// (3, 1, 'local_g3_5')
// (3, 1, 'lutff_7/in_3')
// (3, 1, 'sp4_r_v_b_21')
// (3, 2, 'sp4_r_v_b_8')
// (3, 3, 'local_g3_1')
// (3, 3, 'lutff_2/in_2')
// (3, 3, 'sp4_h_r_21')
// (3, 3, 'sp4_r_v_b_41')
// (3, 4, 'sp4_r_v_b_28')
// (3, 5, 'sp4_r_v_b_17')
// (3, 6, 'sp4_r_v_b_4')
// (3, 7, 'local_g1_1')
// (3, 7, 'lutff_0/in_0')
// (3, 7, 'sp4_h_r_17')
// (3, 7, 'sp4_r_v_b_46')
// (3, 8, 'sp4_r_v_b_35')
// (3, 9, 'sp4_r_v_b_22')
// (3, 10, 'sp4_r_v_b_11')
// (3, 19, 'sp4_h_r_1')
// (4, 0, 'span4_vert_21')
// (4, 1, 'sp4_v_b_21')
// (4, 2, 'sp4_h_r_2')
// (4, 2, 'sp4_h_r_8')
// (4, 2, 'sp4_v_b_8')
// (4, 2, 'sp4_v_t_41')
// (4, 3, 'sp4_h_r_32')
// (4, 3, 'sp4_v_b_41')
// (4, 4, 'sp4_v_b_28')
// (4, 5, 'local_g0_1')
// (4, 5, 'lutff_7/in_0')
// (4, 5, 'sp4_v_b_17')
// (4, 6, 'sp4_h_r_11')
// (4, 6, 'sp4_v_b_4')
// (4, 6, 'sp4_v_t_46')
// (4, 7, 'local_g2_4')
// (4, 7, 'lutff_0/in_2')
// (4, 7, 'sp4_h_r_28')
// (4, 7, 'sp4_v_b_46')
// (4, 8, 'sp4_v_b_35')
// (4, 9, 'sp4_v_b_22')
// (4, 10, 'local_g0_3')
// (4, 10, 'lutff_2/in_1')
// (4, 10, 'sp4_v_b_11')
// (4, 19, 'sp4_h_r_12')
// (5, 2, 'local_g1_7')
// (5, 2, 'lutff_2/in_0')
// (5, 2, 'sp4_h_r_15')
// (5, 2, 'sp4_h_r_21')
// (5, 3, 'sp4_h_r_45')
// (5, 6, 'sp4_h_r_22')
// (5, 7, 'sp4_h_r_41')
// (5, 19, 'local_g3_1')
// (5, 19, 'lutff_2/in_0')
// (5, 19, 'sp4_h_r_25')
// (6, 2, 'sp4_h_r_26')
// (6, 2, 'sp4_h_r_32')
// (6, 3, 'sp4_h_l_45')
// (6, 3, 'sp4_h_r_5')
// (6, 6, 'sp4_h_r_35')
// (6, 7, 'sp4_h_l_41')
// (6, 7, 'sp4_h_r_8')
// (6, 19, 'sp4_h_r_36')
// (7, 1, 'sp4_r_v_b_22')
// (7, 2, 'sp4_h_r_39')
// (7, 2, 'sp4_h_r_45')
// (7, 2, 'sp4_r_v_b_11')
// (7, 3, 'local_g3_5')
// (7, 3, 'lutff_2/in_2')
// (7, 3, 'sp4_h_r_16')
// (7, 3, 'sp4_r_v_b_38')
// (7, 3, 'sp4_r_v_b_45')
// (7, 4, 'sp4_r_v_b_27')
// (7, 4, 'sp4_r_v_b_32')
// (7, 5, 'sp4_r_v_b_14')
// (7, 5, 'sp4_r_v_b_21')
// (7, 6, 'sp4_h_r_46')
// (7, 6, 'sp4_r_v_b_3')
// (7, 6, 'sp4_r_v_b_8')
// (7, 7, 'sp4_h_r_21')
// (7, 7, 'sp4_r_v_b_38')
// (7, 8, 'sp4_h_r_6')
// (7, 8, 'sp4_r_v_b_27')
// (7, 9, 'sp4_r_v_b_14')
// (7, 10, 'sp4_r_v_b_3')
// (7, 11, 'sp4_r_v_b_38')
// (7, 12, 'sp4_r_v_b_27')
// (7, 13, 'sp4_r_v_b_14')
// (7, 14, 'sp4_r_v_b_3')
// (7, 19, 'sp4_h_l_36')
// (7, 19, 'sp4_h_r_1')
// (7, 20, 'sp4_h_r_8')
// (8, 0, 'span4_vert_22')
// (8, 1, 'local_g1_6')
// (8, 1, 'lutff_5/in_0')
// (8, 1, 'sp4_v_b_22')
// (8, 2, 'sp4_h_l_39')
// (8, 2, 'sp4_h_l_45')
// (8, 2, 'sp4_h_r_5')
// (8, 2, 'sp4_v_b_11')
// (8, 2, 'sp4_v_t_38')
// (8, 2, 'sp4_v_t_45')
// (8, 3, 'local_g3_6')
// (8, 3, 'lutff_6/in_3')
// (8, 3, 'sp4_h_r_29')
// (8, 3, 'sp4_v_b_38')
// (8, 3, 'sp4_v_b_45')
// (8, 4, 'sp4_v_b_27')
// (8, 4, 'sp4_v_b_32')
// (8, 5, 'sp4_v_b_14')
// (8, 5, 'sp4_v_b_21')
// (8, 6, 'sp4_h_l_46')
// (8, 6, 'sp4_h_r_3')
// (8, 6, 'sp4_v_b_3')
// (8, 6, 'sp4_v_b_8')
// (8, 6, 'sp4_v_t_38')
// (8, 7, 'sp4_h_r_32')
// (8, 7, 'sp4_v_b_38')
// (8, 8, 'local_g0_3')
// (8, 8, 'lutff_5/in_0')
// (8, 8, 'sp4_h_r_19')
// (8, 8, 'sp4_v_b_27')
// (8, 9, 'sp4_v_b_14')
// (8, 10, 'sp4_v_b_3')
// (8, 10, 'sp4_v_t_38')
// (8, 11, 'sp4_v_b_38')
// (8, 12, 'sp4_v_b_27')
// (8, 13, 'local_g0_6')
// (8, 13, 'lutff_3/in_1')
// (8, 13, 'sp4_v_b_14')
// (8, 14, 'sp4_h_r_2')
// (8, 14, 'sp4_v_b_3')
// (8, 19, 'sp4_h_r_12')
// (8, 20, 'local_g1_5')
// (8, 20, 'lutff_2/in_2')
// (8, 20, 'sp4_h_r_21')
// (9, 1, 'sp4_r_v_b_26')
// (9, 2, 'sp4_h_r_16')
// (9, 2, 'sp4_r_v_b_15')
// (9, 3, 'local_g1_2')
// (9, 3, 'lutff_0/in_3')
// (9, 3, 'sp4_h_r_40')
// (9, 3, 'sp4_r_v_b_2')
// (9, 6, 'sp4_h_r_14')
// (9, 7, 'sp4_h_r_45')
// (9, 8, 'sp4_h_r_30')
// (9, 14, 'local_g0_7')
// (9, 14, 'lutff_3/in_2')
// (9, 14, 'sp4_h_r_15')
// (9, 19, 'sp4_h_r_25')
// (9, 20, 'sp4_h_r_32')
// (10, 0, 'span4_vert_26')
// (10, 1, 'local_g3_2')
// (10, 1, 'lutff_3/in_2')
// (10, 1, 'sp4_v_b_26')
// (10, 2, 'sp4_h_r_29')
// (10, 2, 'sp4_v_b_15')
// (10, 3, 'sp4_h_l_40')
// (10, 3, 'sp4_h_r_2')
// (10, 3, 'sp4_v_b_2')
// (10, 6, 'sp4_h_r_27')
// (10, 7, 'sp4_h_l_45')
// (10, 7, 'sp4_h_r_0')
// (10, 8, 'sp4_h_r_43')
// (10, 13, 'sp12_h_r_1')
// (10, 14, 'sp4_h_r_26')
// (10, 14, 'sp4_r_v_b_38')
// (10, 15, 'sp4_r_v_b_27')
// (10, 16, 'sp4_r_v_b_14')
// (10, 16, 'sp4_r_v_b_36')
// (10, 17, 'local_g1_3')
// (10, 17, 'lutff_5/in_1')
// (10, 17, 'sp4_r_v_b_25')
// (10, 17, 'sp4_r_v_b_3')
// (10, 18, 'local_g2_4')
// (10, 18, 'lutff_2/in_2')
// (10, 18, 'sp4_r_v_b_12')
// (10, 18, 'sp4_r_v_b_38')
// (10, 19, 'sp4_h_r_36')
// (10, 19, 'sp4_r_v_b_1')
// (10, 19, 'sp4_r_v_b_27')
// (10, 20, 'local_g2_6')
// (10, 20, 'lutff_1/in_3')
// (10, 20, 'sp4_h_r_45')
// (10, 20, 'sp4_r_v_b_14')
// (10, 21, 'sp4_r_v_b_3')
// (11, 0, 'span12_vert_10')
// (11, 1, 'sp12_v_b_10')
// (11, 2, 'sp12_v_b_9')
// (11, 2, 'sp4_h_r_40')
// (11, 3, 'sp12_v_b_6')
// (11, 3, 'sp4_h_r_15')
// (11, 4, 'local_g3_5')
// (11, 4, 'lutff_4/in_0')
// (11, 4, 'sp12_v_b_5')
// (11, 5, 'sp12_v_b_2')
// (11, 6, 'sp12_h_r_1')
// (11, 6, 'sp12_v_b_1')
// (11, 6, 'sp12_v_t_22')
// (11, 6, 'sp4_h_r_38')
// (11, 7, 'sp12_v_b_22')
// (11, 7, 'sp4_h_r_13')
// (11, 7, 'sp4_r_v_b_43')
// (11, 8, 'sp12_v_b_21')
// (11, 8, 'sp4_h_l_43')
// (11, 8, 'sp4_h_r_3')
// (11, 8, 'sp4_r_v_b_30')
// (11, 9, 'sp12_v_b_18')
// (11, 9, 'sp4_r_v_b_19')
// (11, 10, 'sp12_v_b_17')
// (11, 10, 'sp4_r_v_b_6')
// (11, 11, 'sp12_v_b_14')
// (11, 11, 'sp4_r_v_b_39')
// (11, 12, 'sp12_v_b_13')
// (11, 12, 'sp4_r_v_b_26')
// (11, 13, 'local_g0_2')
// (11, 13, 'lutff_3/in_3')
// (11, 13, 'sp12_h_r_2')
// (11, 13, 'sp12_v_b_10')
// (11, 13, 'sp4_r_v_b_15')
// (11, 13, 'sp4_v_t_38')
// (11, 14, 'sp12_v_b_9')
// (11, 14, 'sp4_h_r_39')
// (11, 14, 'sp4_r_v_b_2')
// (11, 14, 'sp4_v_b_38')
// (11, 15, 'sp12_v_b_6')
// (11, 15, 'sp4_v_b_27')
// (11, 15, 'sp4_v_t_36')
// (11, 16, 'sp12_v_b_5')
// (11, 16, 'sp4_v_b_14')
// (11, 16, 'sp4_v_b_36')
// (11, 17, 'sp12_v_b_2')
// (11, 17, 'sp4_v_b_25')
// (11, 17, 'sp4_v_b_3')
// (11, 17, 'sp4_v_t_38')
// (11, 18, 'sp12_v_b_1')
// (11, 18, 'sp4_v_b_12')
// (11, 18, 'sp4_v_b_38')
// (11, 19, 'sp4_h_l_36')
// (11, 19, 'sp4_v_b_1')
// (11, 19, 'sp4_v_b_27')
// (11, 20, 'sp4_h_l_45')
// (11, 20, 'sp4_h_r_0')
// (11, 20, 'sp4_v_b_14')
// (11, 21, 'sp4_v_b_3')
// (12, 2, 'sp4_h_l_40')
// (12, 2, 'sp4_h_r_5')
// (12, 3, 'sp4_h_r_26')
// (12, 3, 'sp4_r_v_b_44')
// (12, 4, 'sp4_r_v_b_33')
// (12, 5, 'local_g3_4')
// (12, 5, 'lutff_5/in_2')
// (12, 5, 'sp4_r_v_b_20')
// (12, 6, 'sp12_h_r_2')
// (12, 6, 'sp4_h_l_38')
// (12, 6, 'sp4_h_r_0')
// (12, 6, 'sp4_r_v_b_9')
// (12, 6, 'sp4_v_t_43')
// (12, 7, 'sp4_h_r_24')
// (12, 7, 'sp4_v_b_43')
// (12, 8, 'sp4_h_r_14')
// (12, 8, 'sp4_v_b_30')
// (12, 9, 'sp4_v_b_19')
// (12, 10, 'local_g0_6')
// (12, 10, 'lutff_2/in_0')
// (12, 10, 'sp4_v_b_6')
// (12, 10, 'sp4_v_t_39')
// (12, 11, 'sp4_v_b_39')
// (12, 12, 'sp4_v_b_26')
// (12, 13, 'sp12_h_r_5')
// (12, 13, 'sp4_v_b_15')
// (12, 14, 'sp4_h_l_39')
// (12, 14, 'sp4_v_b_2')
// (12, 20, 'local_g1_5')
// (12, 20, 'lutff_7/in_1')
// (12, 20, 'sp4_h_r_13')
// (13, 1, 'sp4_r_v_b_28')
// (13, 2, 'local_g3_1')
// (13, 2, 'lutff_3/in_3')
// (13, 2, 'sp4_h_r_16')
// (13, 2, 'sp4_r_v_b_17')
// (13, 2, 'sp4_v_t_44')
// (13, 3, 'sp4_h_r_39')
// (13, 3, 'sp4_r_v_b_4')
// (13, 3, 'sp4_v_b_44')
// (13, 4, 'sp4_v_b_33')
// (13, 5, 'sp4_v_b_20')
// (13, 6, 'sp12_h_r_5')
// (13, 6, 'sp4_h_r_13')
// (13, 6, 'sp4_h_r_9')
// (13, 6, 'sp4_v_b_9')
// (13, 7, 'sp4_h_r_37')
// (13, 8, 'sp4_h_r_27')
// (13, 13, 'sp12_h_r_6')
// (13, 20, 'sp4_h_r_24')
// (14, 0, 'span4_vert_28')
// (14, 1, 'sp4_v_b_28')
// (14, 2, 'sp4_h_r_29')
// (14, 2, 'sp4_v_b_17')
// (14, 3, 'sp4_h_l_39')
// (14, 3, 'sp4_h_r_11')
// (14, 3, 'sp4_v_b_4')
// (14, 5, 'local_g0_7')
// (14, 5, 'lutff_6/in_1')
// (14, 5, 'sp4_h_r_7')
// (14, 6, 'local_g1_6')
// (14, 6, 'lutff_7/in_0')
// (14, 6, 'sp12_h_r_6')
// (14, 6, 'sp4_h_r_20')
// (14, 6, 'sp4_h_r_24')
// (14, 7, 'sp4_h_l_37')
// (14, 7, 'sp4_h_r_4')
// (14, 8, 'sp4_h_r_38')
// (14, 13, 'sp12_h_r_9')
// (14, 17, 'sp4_r_v_b_42')
// (14, 18, 'sp4_r_v_b_31')
// (14, 19, 'sp4_r_v_b_18')
// (14, 20, 'sp4_h_r_37')
// (14, 20, 'sp4_r_v_b_7')
// (15, 1, 'sp4_r_v_b_16')
// (15, 2, 'local_g1_5')
// (15, 2, 'lutff_2/in_0')
// (15, 2, 'sp4_h_r_40')
// (15, 2, 'sp4_r_v_b_5')
// (15, 3, 'local_g1_6')
// (15, 3, 'lutff_0/in_1')
// (15, 3, 'sp4_h_r_22')
// (15, 3, 'sp4_r_v_b_42')
// (15, 4, 'sp4_r_v_b_31')
// (15, 5, 'local_g3_2')
// (15, 5, 'lutff_6/in_3')
// (15, 5, 'sp4_h_r_18')
// (15, 5, 'sp4_r_v_b_18')
// (15, 6, 'sp12_h_r_9')
// (15, 6, 'sp4_h_r_33')
// (15, 6, 'sp4_h_r_37')
// (15, 6, 'sp4_r_v_b_7')
// (15, 7, 'sp4_h_r_17')
// (15, 8, 'sp4_h_l_38')
// (15, 8, 'sp4_h_r_7')
// (15, 13, 'sp12_h_r_10')
// (15, 16, 'sp4_h_r_1')
// (15, 16, 'sp4_v_t_42')
// (15, 17, 'sp4_v_b_42')
// (15, 18, 'sp4_v_b_31')
// (15, 19, 'sp4_v_b_18')
// (15, 20, 'sp4_h_l_37')
// (15, 20, 'sp4_v_b_7')
// (16, 0, 'span4_vert_16')
// (16, 1, 'sp4_v_b_16')
// (16, 2, 'sp4_h_l_40')
// (16, 2, 'sp4_h_r_5')
// (16, 2, 'sp4_v_b_5')
// (16, 2, 'sp4_v_t_42')
// (16, 3, 'local_g3_3')
// (16, 3, 'lutff_7/in_3')
// (16, 3, 'sp4_h_r_35')
// (16, 3, 'sp4_v_b_42')
// (16, 4, 'sp4_v_b_31')
// (16, 5, 'sp4_h_r_31')
// (16, 5, 'sp4_v_b_18')
// (16, 6, 'sp12_h_r_10')
// (16, 6, 'sp4_h_l_37')
// (16, 6, 'sp4_h_r_2')
// (16, 6, 'sp4_h_r_44')
// (16, 6, 'sp4_h_r_9')
// (16, 6, 'sp4_v_b_7')
// (16, 7, 'sp4_h_r_28')
// (16, 8, 'sp4_h_r_18')
// (16, 13, 'sp12_h_r_13')
// (16, 16, 'sp4_h_r_12')
// (17, 2, 'sp4_h_r_16')
// (17, 3, 'sp4_h_r_46')
// (17, 5, 'sp4_h_r_42')
// (17, 6, 'sp12_h_r_13')
// (17, 6, 'sp4_h_l_44')
// (17, 6, 'sp4_h_r_15')
// (17, 6, 'sp4_h_r_20')
// (17, 6, 'sp4_h_r_6')
// (17, 7, 'sp4_h_r_41')
// (17, 8, 'sp4_h_r_31')
// (17, 13, 'sp12_h_r_14')
// (17, 16, 'sp4_h_r_25')
// (18, 2, 'sp4_h_r_29')
// (18, 3, 'sp4_h_l_46')
// (18, 3, 'sp4_h_r_3')
// (18, 5, 'sp4_h_l_42')
// (18, 5, 'sp4_h_r_11')
// (18, 6, 'sp12_h_r_14')
// (18, 6, 'sp4_h_r_19')
// (18, 6, 'sp4_h_r_26')
// (18, 6, 'sp4_h_r_33')
// (18, 7, 'sp4_h_l_41')
// (18, 7, 'sp4_h_r_8')
// (18, 8, 'sp4_h_r_42')
// (18, 9, 'sp4_r_v_b_36')
// (18, 10, 'sp4_r_v_b_25')
// (18, 11, 'sp4_r_v_b_12')
// (18, 12, 'sp4_r_v_b_1')
// (18, 13, 'sp12_h_r_17')
// (18, 13, 'sp4_r_v_b_36')
// (18, 14, 'sp4_r_v_b_25')
// (18, 15, 'sp4_r_v_b_12')
// (18, 16, 'sp4_h_r_36')
// (18, 16, 'sp4_r_v_b_1')
// (19, 2, 'sp4_h_r_40')
// (19, 3, 'sp4_h_r_14')
// (19, 3, 'sp4_r_v_b_46')
// (19, 4, 'sp4_r_v_b_35')
// (19, 5, 'sp4_h_r_22')
// (19, 5, 'sp4_r_v_b_22')
// (19, 6, 'sp12_h_r_17')
// (19, 6, 'sp4_h_r_30')
// (19, 6, 'sp4_h_r_39')
// (19, 6, 'sp4_h_r_44')
// (19, 6, 'sp4_r_v_b_11')
// (19, 7, 'sp4_h_r_21')
// (19, 8, 'sp4_h_l_42')
// (19, 8, 'sp4_h_r_7')
// (19, 8, 'sp4_v_t_36')
// (19, 9, 'sp4_v_b_36')
// (19, 10, 'sp4_v_b_25')
// (19, 11, 'sp4_v_b_12')
// (19, 12, 'sp4_v_b_1')
// (19, 12, 'sp4_v_t_36')
// (19, 13, 'sp12_h_r_18')
// (19, 13, 'sp4_v_b_36')
// (19, 14, 'sp4_v_b_25')
// (19, 15, 'sp4_v_b_12')
// (19, 16, 'sp4_h_l_36')
// (19, 16, 'sp4_v_b_1')
// (20, 2, 'sp4_h_l_40')
// (20, 2, 'sp4_v_t_46')
// (20, 3, 'sp4_h_r_27')
// (20, 3, 'sp4_v_b_46')
// (20, 4, 'sp4_v_b_35')
// (20, 5, 'sp4_h_r_35')
// (20, 5, 'sp4_v_b_22')
// (20, 6, 'sp12_h_r_18')
// (20, 6, 'sp4_h_l_39')
// (20, 6, 'sp4_h_l_44')
// (20, 6, 'sp4_h_r_43')
// (20, 6, 'sp4_h_r_6')
// (20, 6, 'sp4_v_b_11')
// (20, 7, 'sp4_h_r_32')
// (20, 8, 'sp4_h_r_18')
// (20, 13, 'sp12_h_r_21')
// (21, 3, 'sp4_h_r_38')
// (21, 4, 'sp4_r_v_b_38')
// (21, 5, 'neigh_op_tnr_7')
// (21, 5, 'sp4_h_r_46')
// (21, 5, 'sp4_r_v_b_27')
// (21, 6, 'neigh_op_rgt_7')
// (21, 6, 'sp12_h_r_21')
// (21, 6, 'sp4_h_l_43')
// (21, 6, 'sp4_h_r_19')
// (21, 6, 'sp4_h_r_3')
// (21, 6, 'sp4_r_v_b_14')
// (21, 6, 'sp4_r_v_b_46')
// (21, 7, 'neigh_op_bnr_7')
// (21, 7, 'sp4_h_r_45')
// (21, 7, 'sp4_r_v_b_3')
// (21, 7, 'sp4_r_v_b_35')
// (21, 8, 'sp4_h_r_31')
// (21, 8, 'sp4_r_v_b_22')
// (21, 9, 'sp4_r_v_b_11')
// (21, 13, 'sp12_h_r_22')
// (22, 1, 'sp12_v_t_22')
// (22, 2, 'sp12_v_b_22')
// (22, 3, 'sp12_v_b_21')
// (22, 3, 'sp4_h_l_38')
// (22, 3, 'sp4_v_t_38')
// (22, 4, 'sp12_v_b_18')
// (22, 4, 'sp4_v_b_38')
// (22, 5, 'neigh_op_top_7')
// (22, 5, 'sp12_v_b_17')
// (22, 5, 'sp4_h_l_46')
// (22, 5, 'sp4_r_v_b_42')
// (22, 5, 'sp4_v_b_27')
// (22, 5, 'sp4_v_t_46')
// (22, 6, 'lutff_7/out')
// (22, 6, 'sp12_h_r_22')
// (22, 6, 'sp12_v_b_14')
// (22, 6, 'sp4_h_r_14')
// (22, 6, 'sp4_h_r_30')
// (22, 6, 'sp4_r_v_b_31')
// (22, 6, 'sp4_v_b_14')
// (22, 6, 'sp4_v_b_46')
// (22, 7, 'neigh_op_bot_7')
// (22, 7, 'sp12_v_b_13')
// (22, 7, 'sp4_h_l_45')
// (22, 7, 'sp4_r_v_b_18')
// (22, 7, 'sp4_v_b_3')
// (22, 7, 'sp4_v_b_35')
// (22, 8, 'sp12_v_b_10')
// (22, 8, 'sp4_h_r_42')
// (22, 8, 'sp4_r_v_b_7')
// (22, 8, 'sp4_v_b_22')
// (22, 9, 'sp12_v_b_9')
// (22, 9, 'sp4_v_b_11')
// (22, 10, 'sp12_v_b_6')
// (22, 11, 'sp12_v_b_5')
// (22, 12, 'sp12_v_b_2')
// (22, 13, 'sp12_h_l_22')
// (22, 13, 'sp12_v_b_1')
// (23, 4, 'sp4_v_t_42')
// (23, 5, 'neigh_op_tnl_7')
// (23, 5, 'sp4_v_b_42')
// (23, 6, 'neigh_op_lft_7')
// (23, 6, 'sp12_h_l_22')
// (23, 6, 'sp4_h_r_27')
// (23, 6, 'sp4_h_r_43')
// (23, 6, 'sp4_v_b_31')
// (23, 7, 'neigh_op_bnl_7')
// (23, 7, 'sp4_v_b_18')
// (23, 8, 'sp4_h_l_42')
// (23, 8, 'sp4_v_b_7')
// (24, 6, 'sp4_h_l_43')
// (24, 6, 'sp4_h_r_38')
// (25, 6, 'sp4_h_l_38')

reg n180 = 0;
// (1, 2, 'neigh_op_tnr_0')
// (1, 3, 'neigh_op_rgt_0')
// (1, 4, 'neigh_op_bnr_0')
// (2, 2, 'neigh_op_top_0')
// (2, 3, 'local_g0_0')
// (2, 3, 'lutff_0/out')
// (2, 3, 'lutff_1/in_1')
// (2, 3, 'lutff_5/in_1')
// (2, 4, 'neigh_op_bot_0')
// (3, 2, 'neigh_op_tnl_0')
// (3, 3, 'neigh_op_lft_0')
// (3, 4, 'neigh_op_bnl_0')

reg n181 = 0;
// (1, 2, 'neigh_op_tnr_1')
// (1, 3, 'neigh_op_rgt_1')
// (1, 4, 'neigh_op_bnr_1')
// (2, 2, 'neigh_op_top_1')
// (2, 3, 'local_g2_1')
// (2, 3, 'lutff_1/out')
// (2, 3, 'lutff_6/in_3')
// (2, 4, 'local_g1_1')
// (2, 4, 'lutff_2/in_2')
// (2, 4, 'neigh_op_bot_1')
// (3, 2, 'neigh_op_tnl_1')
// (3, 3, 'neigh_op_lft_1')
// (3, 4, 'neigh_op_bnl_1')

wire n182;
// (1, 2, 'neigh_op_tnr_2')
// (1, 3, 'neigh_op_rgt_2')
// (1, 4, 'neigh_op_bnr_2')
// (2, 2, 'neigh_op_top_2')
// (2, 3, 'local_g3_2')
// (2, 3, 'lutff_2/out')
// (2, 3, 'lutff_5/in_0')
// (2, 4, 'neigh_op_bot_2')
// (3, 2, 'neigh_op_tnl_2')
// (3, 3, 'neigh_op_lft_2')
// (3, 4, 'neigh_op_bnl_2')

wire n183;
// (1, 2, 'neigh_op_tnr_3')
// (1, 3, 'neigh_op_rgt_3')
// (1, 4, 'neigh_op_bnr_3')
// (2, 2, 'neigh_op_top_3')
// (2, 2, 'sp12_v_t_22')
// (2, 3, 'lutff_3/out')
// (2, 3, 'sp12_v_b_22')
// (2, 4, 'neigh_op_bot_3')
// (2, 4, 'sp12_v_b_21')
// (2, 5, 'sp12_v_b_18')
// (2, 6, 'sp12_v_b_17')
// (2, 7, 'sp12_v_b_14')
// (2, 8, 'sp12_v_b_13')
// (2, 9, 'sp12_v_b_10')
// (2, 10, 'sp12_v_b_9')
// (2, 11, 'sp12_v_b_6')
// (2, 12, 'sp12_v_b_5')
// (2, 13, 'sp12_v_b_2')
// (2, 14, 'local_g2_1')
// (2, 14, 'lutff_1/in_2')
// (2, 14, 'sp12_v_b_1')
// (3, 2, 'neigh_op_tnl_3')
// (3, 3, 'neigh_op_lft_3')
// (3, 4, 'neigh_op_bnl_3')

reg n184 = 0;
// (1, 2, 'neigh_op_tnr_4')
// (1, 3, 'neigh_op_rgt_4')
// (1, 4, 'neigh_op_bnr_4')
// (2, 2, 'neigh_op_top_4')
// (2, 3, 'local_g0_4')
// (2, 3, 'lutff_2/in_2')
// (2, 3, 'lutff_4/out')
// (2, 3, 'lutff_7/in_3')
// (2, 4, 'neigh_op_bot_4')
// (3, 2, 'neigh_op_tnl_4')
// (3, 3, 'neigh_op_lft_4')
// (3, 4, 'neigh_op_bnl_4')

wire n185;
// (1, 2, 'neigh_op_tnr_5')
// (1, 3, 'neigh_op_rgt_5')
// (1, 4, 'neigh_op_bnr_5')
// (2, 2, 'neigh_op_top_5')
// (2, 3, 'local_g1_5')
// (2, 3, 'lutff_3/in_1')
// (2, 3, 'lutff_5/out')
// (2, 4, 'neigh_op_bot_5')
// (3, 2, 'neigh_op_tnl_5')
// (3, 3, 'neigh_op_lft_5')
// (3, 4, 'neigh_op_bnl_5')

reg n186 = 0;
// (1, 2, 'neigh_op_tnr_6')
// (1, 3, 'local_g3_6')
// (1, 3, 'lutff_0/in_1')
// (1, 3, 'lutff_2/in_1')
// (1, 3, 'neigh_op_rgt_6')
// (1, 4, 'neigh_op_bnr_6')
// (2, 2, 'neigh_op_top_6')
// (2, 3, 'lutff_6/out')
// (2, 4, 'neigh_op_bot_6')
// (3, 2, 'neigh_op_tnl_6')
// (3, 3, 'neigh_op_lft_6')
// (3, 4, 'neigh_op_bnl_6')

reg n187 = 0;
// (1, 2, 'neigh_op_tnr_7')
// (1, 3, 'neigh_op_rgt_7')
// (1, 4, 'neigh_op_bnr_7')
// (2, 2, 'neigh_op_top_7')
// (2, 3, 'local_g1_7')
// (2, 3, 'lutff_0/in_0')
// (2, 3, 'lutff_2/in_0')
// (2, 3, 'lutff_7/out')
// (2, 4, 'neigh_op_bot_7')
// (3, 2, 'neigh_op_tnl_7')
// (3, 3, 'neigh_op_lft_7')
// (3, 4, 'neigh_op_bnl_7')

reg n188 = 0;
// (1, 2, 'sp4_h_r_7')
// (2, 2, 'local_g1_2')
// (2, 2, 'lutff_3/in_0')
// (2, 2, 'sp4_h_r_18')
// (2, 2, 'sp4_r_v_b_41')
// (2, 3, 'sp4_r_v_b_28')
// (2, 4, 'sp4_r_v_b_17')
// (2, 5, 'sp4_r_v_b_4')
// (2, 6, 'sp4_r_v_b_36')
// (2, 7, 'sp4_r_v_b_25')
// (2, 8, 'sp4_r_v_b_12')
// (2, 9, 'sp4_r_v_b_1')
// (3, 1, 'local_g1_0')
// (3, 1, 'lutff_1/in_0')
// (3, 1, 'sp4_h_r_0')
// (3, 1, 'sp4_v_t_41')
// (3, 2, 'sp4_h_r_31')
// (3, 2, 'sp4_v_b_41')
// (3, 3, 'sp4_v_b_28')
// (3, 4, 'local_g1_1')
// (3, 4, 'lutff_2/in_0')
// (3, 4, 'sp4_v_b_17')
// (3, 5, 'local_g1_4')
// (3, 5, 'lutff_7/in_0')
// (3, 5, 'sp4_h_r_4')
// (3, 5, 'sp4_v_b_4')
// (3, 5, 'sp4_v_t_36')
// (3, 6, 'sp4_v_b_36')
// (3, 7, 'local_g2_1')
// (3, 7, 'lutff_2/in_3')
// (3, 7, 'sp4_v_b_25')
// (3, 8, 'sp4_v_b_12')
// (3, 9, 'sp4_h_r_8')
// (3, 9, 'sp4_v_b_1')
// (4, 1, 'sp4_h_r_13')
// (4, 2, 'sp4_h_r_42')
// (4, 3, 'sp4_r_v_b_41')
// (4, 4, 'sp4_r_v_b_28')
// (4, 5, 'sp4_h_r_17')
// (4, 5, 'sp4_r_v_b_17')
// (4, 6, 'sp4_r_v_b_4')
// (4, 7, 'sp4_r_v_b_47')
// (4, 8, 'sp4_r_v_b_34')
// (4, 9, 'sp4_h_r_21')
// (4, 9, 'sp4_r_v_b_23')
// (4, 10, 'local_g2_2')
// (4, 10, 'lutff_0/in_0')
// (4, 10, 'sp4_r_v_b_10')
// (4, 11, 'sp4_r_v_b_45')
// (4, 12, 'sp4_r_v_b_32')
// (4, 13, 'sp4_r_v_b_21')
// (4, 14, 'sp4_r_v_b_8')
// (4, 15, 'sp4_r_v_b_46')
// (4, 16, 'sp4_r_v_b_35')
// (4, 17, 'sp4_r_v_b_22')
// (4, 18, 'sp4_r_v_b_11')
// (5, 1, 'sp4_h_r_24')
// (5, 2, 'sp4_h_l_42')
// (5, 2, 'sp4_h_r_4')
// (5, 2, 'sp4_h_r_7')
// (5, 2, 'sp4_v_t_41')
// (5, 3, 'local_g2_1')
// (5, 3, 'lutff_0/in_1')
// (5, 3, 'sp4_v_b_41')
// (5, 4, 'sp4_v_b_28')
// (5, 5, 'sp4_h_r_28')
// (5, 5, 'sp4_v_b_17')
// (5, 6, 'sp4_h_r_4')
// (5, 6, 'sp4_v_b_4')
// (5, 6, 'sp4_v_t_47')
// (5, 7, 'sp4_v_b_47')
// (5, 8, 'sp4_v_b_34')
// (5, 9, 'sp4_h_r_32')
// (5, 9, 'sp4_v_b_23')
// (5, 10, 'sp4_h_r_10')
// (5, 10, 'sp4_h_r_2')
// (5, 10, 'sp4_v_b_10')
// (5, 10, 'sp4_v_t_45')
// (5, 11, 'sp4_v_b_45')
// (5, 12, 'sp4_v_b_32')
// (5, 13, 'sp4_v_b_21')
// (5, 14, 'sp4_v_b_8')
// (5, 14, 'sp4_v_t_46')
// (5, 15, 'sp4_v_b_46')
// (5, 16, 'sp4_v_b_35')
// (5, 17, 'sp4_v_b_22')
// (5, 18, 'local_g1_3')
// (5, 18, 'lutff_0/in_2')
// (5, 18, 'sp4_v_b_11')
// (6, 1, 'sp4_h_r_37')
// (6, 2, 'sp4_h_r_17')
// (6, 2, 'sp4_h_r_18')
// (6, 2, 'sp4_r_v_b_39')
// (6, 3, 'sp4_r_v_b_26')
// (6, 4, 'sp4_r_v_b_15')
// (6, 5, 'sp4_h_r_41')
// (6, 5, 'sp4_r_v_b_2')
// (6, 6, 'sp4_h_r_17')
// (6, 9, 'sp4_h_r_45')
// (6, 10, 'sp4_h_r_15')
// (6, 10, 'sp4_h_r_23')
// (7, 1, 'sp4_h_l_37')
// (7, 1, 'sp4_h_r_9')
// (7, 1, 'sp4_v_t_39')
// (7, 2, 'local_g2_4')
// (7, 2, 'lutff_7/in_3')
// (7, 2, 'sp4_h_r_28')
// (7, 2, 'sp4_h_r_31')
// (7, 2, 'sp4_v_b_39')
// (7, 3, 'local_g2_2')
// (7, 3, 'lutff_5/in_3')
// (7, 3, 'sp4_v_b_26')
// (7, 4, 'sp4_v_b_15')
// (7, 5, 'sp4_h_l_41')
// (7, 5, 'sp4_h_r_8')
// (7, 5, 'sp4_h_r_9')
// (7, 5, 'sp4_v_b_2')
// (7, 6, 'sp4_h_r_28')
// (7, 6, 'sp4_r_v_b_45')
// (7, 7, 'sp4_r_v_b_32')
// (7, 8, 'sp4_r_v_b_21')
// (7, 9, 'sp4_h_l_45')
// (7, 9, 'sp4_h_r_0')
// (7, 9, 'sp4_r_v_b_8')
// (7, 10, 'sp4_h_r_26')
// (7, 10, 'sp4_h_r_34')
// (7, 13, 'sp4_h_r_9')
// (8, 1, 'local_g3_4')
// (8, 1, 'lutff_2/in_3')
// (8, 1, 'sp4_h_r_20')
// (8, 1, 'sp4_r_v_b_20')
// (8, 2, 'sp4_h_r_41')
// (8, 2, 'sp4_h_r_42')
// (8, 2, 'sp4_r_v_b_9')
// (8, 3, 'local_g3_3')
// (8, 3, 'lutff_5/in_1')
// (8, 3, 'sp4_r_v_b_43')
// (8, 4, 'sp4_r_v_b_30')
// (8, 5, 'sp4_h_r_20')
// (8, 5, 'sp4_h_r_21')
// (8, 5, 'sp4_r_v_b_19')
// (8, 5, 'sp4_v_t_45')
// (8, 6, 'sp4_h_r_41')
// (8, 6, 'sp4_r_v_b_6')
// (8, 6, 'sp4_v_b_45')
// (8, 7, 'sp4_v_b_32')
// (8, 8, 'local_g0_5')
// (8, 8, 'lutff_2/in_1')
// (8, 8, 'sp4_v_b_21')
// (8, 9, 'sp4_h_r_13')
// (8, 9, 'sp4_h_r_3')
// (8, 9, 'sp4_v_b_8')
// (8, 10, 'sp4_h_r_39')
// (8, 10, 'sp4_h_r_47')
// (8, 13, 'local_g0_4')
// (8, 13, 'lutff_5/in_3')
// (8, 13, 'sp4_h_r_20')
// (9, 0, 'span4_vert_20')
// (9, 1, 'local_g3_4')
// (9, 1, 'lutff_5/in_0')
// (9, 1, 'sp4_h_r_33')
// (9, 1, 'sp4_r_v_b_20')
// (9, 1, 'sp4_v_b_20')
// (9, 2, 'sp4_h_l_41')
// (9, 2, 'sp4_h_l_42')
// (9, 2, 'sp4_h_r_11')
// (9, 2, 'sp4_h_r_4')
// (9, 2, 'sp4_r_v_b_9')
// (9, 2, 'sp4_v_b_9')
// (9, 2, 'sp4_v_t_43')
// (9, 3, 'sp4_v_b_43')
// (9, 4, 'sp4_v_b_30')
// (9, 5, 'sp4_h_r_32')
// (9, 5, 'sp4_h_r_33')
// (9, 5, 'sp4_v_b_19')
// (9, 6, 'sp4_h_l_41')
// (9, 6, 'sp4_h_r_1')
// (9, 6, 'sp4_v_b_6')
// (9, 9, 'sp4_h_r_14')
// (9, 9, 'sp4_h_r_24')
// (9, 10, 'sp4_h_l_39')
// (9, 10, 'sp4_h_l_47')
// (9, 10, 'sp4_h_r_2')
// (9, 13, 'sp4_h_r_33')
// (9, 27, 'sp4_r_v_b_40')
// (9, 28, 'sp4_r_v_b_29')
// (9, 29, 'sp4_r_v_b_16')
// (9, 30, 'sp4_r_v_b_5')
// (10, 0, 'span12_vert_17')
// (10, 0, 'span4_vert_20')
// (10, 1, 'sp12_v_b_17')
// (10, 1, 'sp4_h_r_44')
// (10, 1, 'sp4_v_b_20')
// (10, 2, 'sp12_v_b_14')
// (10, 2, 'sp4_h_r_17')
// (10, 2, 'sp4_h_r_22')
// (10, 2, 'sp4_r_v_b_44')
// (10, 2, 'sp4_v_b_9')
// (10, 3, 'sp12_v_b_13')
// (10, 3, 'sp4_r_v_b_33')
// (10, 4, 'sp12_v_b_10')
// (10, 4, 'sp4_r_v_b_20')
// (10, 5, 'sp12_v_b_9')
// (10, 5, 'sp4_h_r_44')
// (10, 5, 'sp4_h_r_45')
// (10, 5, 'sp4_r_v_b_9')
// (10, 6, 'sp12_v_b_6')
// (10, 6, 'sp4_h_r_12')
// (10, 6, 'sp4_r_v_b_44')
// (10, 7, 'sp12_v_b_5')
// (10, 7, 'sp4_r_v_b_33')
// (10, 8, 'sp12_v_b_2')
// (10, 8, 'sp4_r_v_b_20')
// (10, 9, 'sp12_h_r_1')
// (10, 9, 'sp12_v_b_1')
// (10, 9, 'sp12_v_t_22')
// (10, 9, 'sp4_h_r_27')
// (10, 9, 'sp4_h_r_37')
// (10, 9, 'sp4_r_v_b_9')
// (10, 10, 'sp12_v_b_22')
// (10, 10, 'sp4_h_r_15')
// (10, 10, 'sp4_r_v_b_44')
// (10, 11, 'sp12_v_b_21')
// (10, 11, 'sp4_r_v_b_33')
// (10, 12, 'sp12_v_b_18')
// (10, 12, 'sp4_r_v_b_20')
// (10, 13, 'sp12_v_b_17')
// (10, 13, 'sp4_h_r_44')
// (10, 13, 'sp4_r_v_b_9')
// (10, 14, 'sp12_v_b_14')
// (10, 14, 'sp4_r_v_b_44')
// (10, 15, 'sp12_v_b_13')
// (10, 15, 'sp4_r_v_b_33')
// (10, 16, 'sp12_v_b_10')
// (10, 16, 'sp4_r_v_b_20')
// (10, 17, 'sp12_v_b_9')
// (10, 17, 'sp4_r_v_b_9')
// (10, 18, 'local_g2_6')
// (10, 18, 'lutff_0/in_2')
// (10, 18, 'sp12_v_b_6')
// (10, 18, 'sp4_r_v_b_44')
// (10, 19, 'local_g3_5')
// (10, 19, 'lutff_2/in_2')
// (10, 19, 'sp12_v_b_5')
// (10, 19, 'sp4_r_v_b_33')
// (10, 20, 'sp12_v_b_2')
// (10, 20, 'sp4_r_v_b_20')
// (10, 21, 'sp12_v_b_1')
// (10, 21, 'sp12_v_t_22')
// (10, 21, 'sp4_r_v_b_9')
// (10, 22, 'sp12_v_b_22')
// (10, 23, 'sp12_v_b_21')
// (10, 24, 'sp12_v_b_18')
// (10, 25, 'sp12_v_b_17')
// (10, 26, 'sp12_v_b_14')
// (10, 26, 'sp4_v_t_40')
// (10, 27, 'sp12_v_b_13')
// (10, 27, 'sp4_v_b_40')
// (10, 28, 'sp12_v_b_10')
// (10, 28, 'sp4_v_b_29')
// (10, 29, 'sp12_v_b_9')
// (10, 29, 'sp4_v_b_16')
// (10, 30, 'sp12_v_b_6')
// (10, 30, 'sp4_h_r_5')
// (10, 30, 'sp4_v_b_5')
// (10, 31, 'span12_vert_5')
// (11, 1, 'sp4_h_l_44')
// (11, 1, 'sp4_h_r_9')
// (11, 1, 'sp4_v_t_44')
// (11, 2, 'local_g2_4')
// (11, 2, 'lutff_4/in_0')
// (11, 2, 'sp4_h_r_28')
// (11, 2, 'sp4_h_r_35')
// (11, 2, 'sp4_v_b_44')
// (11, 3, 'local_g2_1')
// (11, 3, 'lutff_1/in_0')
// (11, 3, 'sp4_v_b_33')
// (11, 4, 'sp4_v_b_20')
// (11, 5, 'sp4_h_l_44')
// (11, 5, 'sp4_h_l_45')
// (11, 5, 'sp4_h_r_8')
// (11, 5, 'sp4_v_b_9')
// (11, 5, 'sp4_v_t_44')
// (11, 6, 'local_g3_4')
// (11, 6, 'lutff_6/in_1')
// (11, 6, 'sp4_h_r_25')
// (11, 6, 'sp4_r_v_b_37')
// (11, 6, 'sp4_r_v_b_39')
// (11, 6, 'sp4_v_b_44')
// (11, 7, 'sp4_r_v_b_24')
// (11, 7, 'sp4_r_v_b_26')
// (11, 7, 'sp4_v_b_33')
// (11, 8, 'sp4_r_v_b_13')
// (11, 8, 'sp4_r_v_b_15')
// (11, 8, 'sp4_v_b_20')
// (11, 9, 'sp12_h_r_2')
// (11, 9, 'sp4_h_l_37')
// (11, 9, 'sp4_h_r_38')
// (11, 9, 'sp4_h_r_9')
// (11, 9, 'sp4_r_v_b_0')
// (11, 9, 'sp4_r_v_b_2')
// (11, 9, 'sp4_v_b_9')
// (11, 9, 'sp4_v_t_44')
// (11, 10, 'sp4_h_r_26')
// (11, 10, 'sp4_v_b_44')
// (11, 11, 'sp4_v_b_33')
// (11, 12, 'sp4_v_b_20')
// (11, 13, 'sp4_h_l_44')
// (11, 13, 'sp4_v_b_9')
// (11, 13, 'sp4_v_t_44')
// (11, 14, 'sp4_v_b_44')
// (11, 15, 'sp4_v_b_33')
// (11, 16, 'sp4_v_b_20')
// (11, 17, 'local_g1_1')
// (11, 17, 'lutff_5/in_1')
// (11, 17, 'sp4_v_b_9')
// (11, 17, 'sp4_v_t_44')
// (11, 18, 'sp4_v_b_44')
// (11, 19, 'sp4_v_b_33')
// (11, 20, 'local_g1_4')
// (11, 20, 'lutff_3/in_2')
// (11, 20, 'sp4_v_b_20')
// (11, 21, 'sp4_v_b_9')
// (11, 30, 'local_g1_0')
// (11, 30, 'lutff_0/in_1')
// (11, 30, 'sp4_h_r_16')
// (12, 1, 'sp4_h_r_20')
// (12, 2, 'sp4_h_r_41')
// (12, 2, 'sp4_h_r_46')
// (12, 3, 'sp4_r_v_b_47')
// (12, 4, 'sp4_r_v_b_34')
// (12, 5, 'sp4_h_r_21')
// (12, 5, 'sp4_r_v_b_23')
// (12, 5, 'sp4_v_t_37')
// (12, 5, 'sp4_v_t_39')
// (12, 6, 'sp4_h_r_36')
// (12, 6, 'sp4_r_v_b_10')
// (12, 6, 'sp4_v_b_37')
// (12, 6, 'sp4_v_b_39')
// (12, 7, 'local_g2_0')
// (12, 7, 'lutff_6/in_2')
// (12, 7, 'sp4_v_b_24')
// (12, 7, 'sp4_v_b_26')
// (12, 8, 'local_g0_7')
// (12, 8, 'lutff_4/in_3')
// (12, 8, 'sp4_v_b_13')
// (12, 8, 'sp4_v_b_15')
// (12, 9, 'sp12_h_r_5')
// (12, 9, 'sp4_h_l_38')
// (12, 9, 'sp4_h_r_20')
// (12, 9, 'sp4_h_r_7')
// (12, 9, 'sp4_h_r_9')
// (12, 9, 'sp4_v_b_0')
// (12, 9, 'sp4_v_b_2')
// (12, 10, 'sp4_h_r_39')
// (12, 30, 'sp4_h_r_29')
// (13, 1, 'sp4_h_r_33')
// (13, 2, 'local_g0_2')
// (13, 2, 'lutff_2/in_2')
// (13, 2, 'sp4_h_l_41')
// (13, 2, 'sp4_h_l_46')
// (13, 2, 'sp4_h_r_10')
// (13, 2, 'sp4_h_r_8')
// (13, 2, 'sp4_v_t_47')
// (13, 3, 'sp4_v_b_47')
// (13, 4, 'sp4_v_b_34')
// (13, 5, 'sp4_h_r_32')
// (13, 5, 'sp4_v_b_23')
// (13, 6, 'sp4_h_l_36')
// (13, 6, 'sp4_h_r_5')
// (13, 6, 'sp4_v_b_10')
// (13, 9, 'sp12_h_r_6')
// (13, 9, 'sp4_h_r_18')
// (13, 9, 'sp4_h_r_20')
// (13, 9, 'sp4_h_r_33')
// (13, 10, 'sp4_h_l_39')
// (13, 10, 'sp4_h_r_11')
// (13, 30, 'sp4_h_r_40')
// (14, 1, 'sp4_h_r_44')
// (14, 2, 'sp4_h_r_21')
// (14, 2, 'sp4_h_r_23')
// (14, 2, 'sp4_r_v_b_37')
// (14, 3, 'sp4_r_v_b_24')
// (14, 4, 'sp4_r_v_b_13')
// (14, 5, 'sp4_h_r_45')
// (14, 5, 'sp4_r_v_b_0')
// (14, 6, 'sp4_h_r_16')
// (14, 9, 'sp12_h_r_9')
// (14, 9, 'sp4_h_r_31')
// (14, 9, 'sp4_h_r_33')
// (14, 9, 'sp4_h_r_44')
// (14, 10, 'sp4_h_r_22')
// (14, 30, 'sp4_h_l_40')
// (15, 1, 'sp4_h_l_44')
// (15, 1, 'sp4_h_r_6')
// (15, 1, 'sp4_v_t_37')
// (15, 2, 'sp4_h_r_32')
// (15, 2, 'sp4_h_r_34')
// (15, 2, 'sp4_v_b_37')
// (15, 3, 'local_g2_0')
// (15, 3, 'lutff_2/in_0')
// (15, 3, 'sp4_v_b_24')
// (15, 4, 'sp4_v_b_13')
// (15, 5, 'sp4_h_l_45')
// (15, 5, 'sp4_h_r_0')
// (15, 5, 'sp4_v_b_0')
// (15, 6, 'sp4_h_r_29')
// (15, 9, 'sp12_h_r_10')
// (15, 9, 'sp4_h_l_44')
// (15, 9, 'sp4_h_r_42')
// (15, 9, 'sp4_h_r_44')
// (15, 9, 'sp4_h_r_6')
// (15, 10, 'sp4_h_r_35')
// (16, 1, 'sp4_h_r_19')
// (16, 1, 'sp4_r_v_b_16')
// (16, 2, 'local_g1_5')
// (16, 2, 'lutff_3/in_1')
// (16, 2, 'sp4_h_r_45')
// (16, 2, 'sp4_h_r_47')
// (16, 2, 'sp4_r_v_b_5')
// (16, 3, 'local_g3_4')
// (16, 3, 'lutff_2/in_1')
// (16, 3, 'sp4_r_v_b_44')
// (16, 4, 'sp4_r_v_b_33')
// (16, 5, 'local_g3_4')
// (16, 5, 'lutff_0/in_3')
// (16, 5, 'sp4_h_r_13')
// (16, 5, 'sp4_r_v_b_20')
// (16, 6, 'local_g2_1')
// (16, 6, 'lutff_3/in_0')
// (16, 6, 'sp4_h_r_40')
// (16, 6, 'sp4_r_v_b_9')
// (16, 9, 'sp12_h_r_13')
// (16, 9, 'sp4_h_l_42')
// (16, 9, 'sp4_h_l_44')
// (16, 9, 'sp4_h_r_11')
// (16, 9, 'sp4_h_r_19')
// (16, 9, 'sp4_h_r_6')
// (16, 10, 'sp4_h_r_46')
// (17, 0, 'span4_vert_16')
// (17, 1, 'sp4_h_r_30')
// (17, 1, 'sp4_v_b_16')
// (17, 2, 'sp4_h_l_45')
// (17, 2, 'sp4_h_l_47')
// (17, 2, 'sp4_h_r_0')
// (17, 2, 'sp4_v_b_5')
// (17, 2, 'sp4_v_t_44')
// (17, 3, 'sp4_v_b_44')
// (17, 4, 'sp4_v_b_33')
// (17, 5, 'sp4_h_r_24')
// (17, 5, 'sp4_v_b_20')
// (17, 6, 'sp4_h_l_40')
// (17, 6, 'sp4_h_r_9')
// (17, 6, 'sp4_v_b_9')
// (17, 9, 'sp12_h_r_14')
// (17, 9, 'sp4_h_r_19')
// (17, 9, 'sp4_h_r_22')
// (17, 9, 'sp4_h_r_30')
// (17, 10, 'sp4_h_l_46')
// (17, 10, 'sp4_h_r_3')
// (18, 1, 'sp4_h_r_43')
// (18, 2, 'sp4_h_r_13')
// (18, 2, 'sp4_r_v_b_43')
// (18, 3, 'sp4_r_v_b_30')
// (18, 4, 'sp4_r_v_b_19')
// (18, 5, 'sp4_h_r_37')
// (18, 5, 'sp4_r_v_b_6')
// (18, 6, 'sp4_h_r_20')
// (18, 6, 'sp4_r_v_b_43')
// (18, 7, 'sp4_r_v_b_30')
// (18, 8, 'sp4_r_v_b_19')
// (18, 9, 'sp12_h_r_17')
// (18, 9, 'sp4_h_r_30')
// (18, 9, 'sp4_h_r_35')
// (18, 9, 'sp4_h_r_43')
// (18, 9, 'sp4_r_v_b_6')
// (18, 10, 'sp4_h_r_14')
// (19, 1, 'sp4_h_l_43')
// (19, 1, 'sp4_v_t_43')
// (19, 2, 'sp4_h_r_24')
// (19, 2, 'sp4_v_b_43')
// (19, 3, 'sp4_v_b_30')
// (19, 4, 'sp4_v_b_19')
// (19, 5, 'sp4_h_l_37')
// (19, 5, 'sp4_v_b_6')
// (19, 5, 'sp4_v_t_43')
// (19, 6, 'sp4_h_r_33')
// (19, 6, 'sp4_v_b_43')
// (19, 7, 'sp4_v_b_30')
// (19, 8, 'sp4_v_b_19')
// (19, 9, 'sp12_h_r_18')
// (19, 9, 'sp4_h_l_43')
// (19, 9, 'sp4_h_r_43')
// (19, 9, 'sp4_h_r_46')
// (19, 9, 'sp4_h_r_6')
// (19, 9, 'sp4_v_b_6')
// (19, 10, 'sp4_h_r_27')
// (20, 2, 'sp4_h_r_37')
// (20, 3, 'sp4_r_v_b_43')
// (20, 4, 'sp4_r_v_b_30')
// (20, 5, 'sp4_r_v_b_19')
// (20, 6, 'sp4_h_r_44')
// (20, 6, 'sp4_r_v_b_6')
// (20, 7, 'sp4_r_v_b_38')
// (20, 8, 'neigh_op_tnr_7')
// (20, 8, 'sp4_r_v_b_27')
// (20, 9, 'neigh_op_rgt_7')
// (20, 9, 'sp12_h_r_21')
// (20, 9, 'sp4_h_l_43')
// (20, 9, 'sp4_h_l_46')
// (20, 9, 'sp4_h_r_19')
// (20, 9, 'sp4_h_r_3')
// (20, 9, 'sp4_r_v_b_14')
// (20, 10, 'neigh_op_bnr_7')
// (20, 10, 'sp4_h_r_38')
// (20, 10, 'sp4_r_v_b_3')
// (21, 2, 'sp4_h_l_37')
// (21, 2, 'sp4_v_t_43')
// (21, 3, 'sp4_v_b_43')
// (21, 4, 'sp4_v_b_30')
// (21, 5, 'sp4_v_b_19')
// (21, 6, 'sp4_h_l_44')
// (21, 6, 'sp4_v_b_6')
// (21, 6, 'sp4_v_t_38')
// (21, 7, 'sp4_v_b_38')
// (21, 8, 'neigh_op_top_7')
// (21, 8, 'sp4_v_b_27')
// (21, 9, 'lutff_7/out')
// (21, 9, 'sp12_h_r_22')
// (21, 9, 'sp4_h_r_14')
// (21, 9, 'sp4_h_r_30')
// (21, 9, 'sp4_v_b_14')
// (21, 10, 'neigh_op_bot_7')
// (21, 10, 'sp4_h_l_38')
// (21, 10, 'sp4_v_b_3')
// (22, 8, 'neigh_op_tnl_7')
// (22, 9, 'neigh_op_lft_7')
// (22, 9, 'sp12_h_l_22')
// (22, 9, 'sp4_h_r_27')
// (22, 9, 'sp4_h_r_43')
// (22, 10, 'neigh_op_bnl_7')
// (23, 9, 'sp4_h_l_43')
// (23, 9, 'sp4_h_r_38')
// (24, 9, 'sp4_h_l_38')

reg n189 = 0;
// (1, 2, 'sp4_r_v_b_38')
// (1, 3, 'sp4_r_v_b_27')
// (1, 4, 'sp4_r_v_b_14')
// (1, 5, 'sp4_r_v_b_3')
// (2, 1, 'sp4_h_r_9')
// (2, 1, 'sp4_v_t_38')
// (2, 2, 'local_g3_6')
// (2, 2, 'lutff_7/in_0')
// (2, 2, 'sp4_v_b_38')
// (2, 3, 'sp4_v_b_27')
// (2, 4, 'sp4_v_b_14')
// (2, 5, 'sp4_v_b_3')
// (2, 7, 'sp4_h_r_8')
// (3, 1, 'local_g1_4')
// (3, 1, 'lutff_4/in_3')
// (3, 1, 'sp4_h_r_20')
// (3, 7, 'local_g0_5')
// (3, 7, 'lutff_7/in_0')
// (3, 7, 'sp4_h_r_21')
// (4, 1, 'sp4_h_r_33')
// (4, 1, 'sp4_r_v_b_26')
// (4, 2, 'sp4_r_v_b_15')
// (4, 2, 'sp4_r_v_b_47')
// (4, 3, 'local_g1_2')
// (4, 3, 'lutff_5/in_2')
// (4, 3, 'sp4_r_v_b_2')
// (4, 3, 'sp4_r_v_b_34')
// (4, 4, 'local_g3_7')
// (4, 4, 'lutff_6/in_2')
// (4, 4, 'sp4_r_v_b_23')
// (4, 4, 'sp4_r_v_b_37')
// (4, 4, 'sp4_r_v_b_46')
// (4, 5, 'sp4_r_v_b_10')
// (4, 5, 'sp4_r_v_b_24')
// (4, 5, 'sp4_r_v_b_35')
// (4, 6, 'sp4_r_v_b_13')
// (4, 6, 'sp4_r_v_b_22')
// (4, 7, 'sp4_h_r_32')
// (4, 7, 'sp4_r_v_b_0')
// (4, 7, 'sp4_r_v_b_11')
// (4, 8, 'sp4_r_v_b_38')
// (4, 9, 'sp4_r_v_b_27')
// (4, 10, 'local_g2_6')
// (4, 10, 'lutff_3/in_3')
// (4, 10, 'sp4_r_v_b_14')
// (4, 11, 'sp4_r_v_b_3')
// (5, 0, 'span4_vert_26')
// (5, 1, 'sp4_h_r_4')
// (5, 1, 'sp4_h_r_44')
// (5, 1, 'sp4_v_b_26')
// (5, 1, 'sp4_v_t_47')
// (5, 2, 'sp4_r_v_b_43')
// (5, 2, 'sp4_v_b_15')
// (5, 2, 'sp4_v_b_47')
// (5, 3, 'sp4_h_r_2')
// (5, 3, 'sp4_h_r_5')
// (5, 3, 'sp4_h_r_6')
// (5, 3, 'sp4_r_v_b_30')
// (5, 3, 'sp4_v_b_2')
// (5, 3, 'sp4_v_b_34')
// (5, 3, 'sp4_v_t_37')
// (5, 3, 'sp4_v_t_46')
// (5, 4, 'sp4_r_v_b_19')
// (5, 4, 'sp4_v_b_23')
// (5, 4, 'sp4_v_b_37')
// (5, 4, 'sp4_v_b_46')
// (5, 5, 'local_g1_6')
// (5, 5, 'lutff_6/in_1')
// (5, 5, 'sp4_r_v_b_6')
// (5, 5, 'sp4_v_b_10')
// (5, 5, 'sp4_v_b_24')
// (5, 5, 'sp4_v_b_35')
// (5, 6, 'sp12_h_r_1')
// (5, 6, 'sp12_v_t_22')
// (5, 6, 'sp4_v_b_13')
// (5, 6, 'sp4_v_b_22')
// (5, 7, 'local_g1_3')
// (5, 7, 'lutff_3/in_1')
// (5, 7, 'sp12_v_b_22')
// (5, 7, 'sp4_h_r_45')
// (5, 7, 'sp4_v_b_0')
// (5, 7, 'sp4_v_b_11')
// (5, 7, 'sp4_v_t_38')
// (5, 8, 'sp12_v_b_21')
// (5, 8, 'sp4_v_b_38')
// (5, 9, 'sp12_v_b_18')
// (5, 9, 'sp4_v_b_27')
// (5, 10, 'sp12_v_b_17')
// (5, 10, 'sp4_v_b_14')
// (5, 11, 'sp12_v_b_14')
// (5, 11, 'sp4_v_b_3')
// (5, 12, 'sp12_v_b_13')
// (5, 13, 'sp12_v_b_10')
// (5, 14, 'sp12_v_b_9')
// (5, 15, 'sp12_v_b_6')
// (5, 16, 'sp12_v_b_5')
// (5, 17, 'sp12_v_b_2')
// (5, 18, 'local_g3_1')
// (5, 18, 'lutff_6/in_0')
// (5, 18, 'sp12_h_r_1')
// (5, 18, 'sp12_v_b_1')
// (6, 1, 'sp4_h_l_44')
// (6, 1, 'sp4_h_r_17')
// (6, 1, 'sp4_h_r_6')
// (6, 1, 'sp4_v_t_43')
// (6, 2, 'sp4_v_b_43')
// (6, 3, 'sp4_h_r_15')
// (6, 3, 'sp4_h_r_16')
// (6, 3, 'sp4_h_r_19')
// (6, 3, 'sp4_v_b_30')
// (6, 4, 'sp4_v_b_19')
// (6, 5, 'sp4_v_b_6')
// (6, 6, 'sp12_h_r_2')
// (6, 7, 'sp4_h_l_45')
// (6, 7, 'sp4_h_r_5')
// (6, 18, 'sp12_h_r_2')
// (7, 1, 'local_g0_3')
// (7, 1, 'lutff_3/in_0')
// (7, 1, 'sp4_h_r_19')
// (7, 1, 'sp4_h_r_28')
// (7, 3, 'sp4_h_r_26')
// (7, 3, 'sp4_h_r_29')
// (7, 3, 'sp4_h_r_30')
// (7, 6, 'sp12_h_r_5')
// (7, 7, 'sp4_h_r_16')
// (7, 18, 'sp12_h_r_5')
// (8, 1, 'local_g1_1')
// (8, 1, 'lutff_4/in_0')
// (8, 1, 'sp12_h_r_1')
// (8, 1, 'sp12_v_t_22')
// (8, 1, 'sp4_h_r_30')
// (8, 1, 'sp4_h_r_41')
// (8, 1, 'sp4_r_v_b_26')
// (8, 2, 'sp12_v_b_22')
// (8, 2, 'sp4_r_v_b_15')
// (8, 3, 'local_g1_2')
// (8, 3, 'lutff_3/in_2')
// (8, 3, 'sp12_v_b_21')
// (8, 3, 'sp4_h_r_39')
// (8, 3, 'sp4_h_r_40')
// (8, 3, 'sp4_h_r_43')
// (8, 3, 'sp4_r_v_b_2')
// (8, 4, 'sp12_v_b_18')
// (8, 4, 'sp4_r_v_b_39')
// (8, 5, 'sp12_v_b_17')
// (8, 5, 'sp4_r_v_b_26')
// (8, 6, 'sp12_h_r_6')
// (8, 6, 'sp12_v_b_14')
// (8, 6, 'sp4_r_v_b_15')
// (8, 7, 'sp12_v_b_13')
// (8, 7, 'sp4_h_r_29')
// (8, 7, 'sp4_r_v_b_2')
// (8, 8, 'sp12_v_b_10')
// (8, 8, 'sp4_r_v_b_40')
// (8, 9, 'local_g2_1')
// (8, 9, 'lutff_7/in_2')
// (8, 9, 'sp12_v_b_9')
// (8, 9, 'sp4_r_v_b_29')
// (8, 10, 'sp12_v_b_6')
// (8, 10, 'sp4_r_v_b_16')
// (8, 11, 'sp12_v_b_5')
// (8, 11, 'sp4_r_v_b_5')
// (8, 12, 'sp12_v_b_2')
// (8, 12, 'sp4_r_v_b_40')
// (8, 13, 'local_g3_1')
// (8, 13, 'lutff_1/in_3')
// (8, 13, 'sp12_v_b_1')
// (8, 13, 'sp12_v_t_22')
// (8, 13, 'sp4_r_v_b_29')
// (8, 14, 'sp12_v_b_22')
// (8, 14, 'sp4_r_v_b_16')
// (8, 15, 'sp12_v_b_21')
// (8, 15, 'sp4_r_v_b_5')
// (8, 16, 'sp12_v_b_18')
// (8, 17, 'sp12_v_b_17')
// (8, 18, 'sp12_h_r_6')
// (8, 18, 'sp12_v_b_14')
// (8, 19, 'sp12_v_b_13')
// (8, 20, 'local_g2_2')
// (8, 20, 'lutff_5/in_1')
// (8, 20, 'sp12_v_b_10')
// (8, 21, 'sp12_v_b_9')
// (8, 22, 'sp12_v_b_6')
// (8, 23, 'sp12_v_b_5')
// (8, 24, 'sp12_v_b_2')
// (8, 25, 'sp12_v_b_1')
// (9, 0, 'span4_vert_26')
// (9, 1, 'sp12_h_r_2')
// (9, 1, 'sp4_h_l_41')
// (9, 1, 'sp4_h_r_1')
// (9, 1, 'sp4_h_r_43')
// (9, 1, 'sp4_v_b_26')
// (9, 2, 'sp4_r_v_b_38')
// (9, 2, 'sp4_r_v_b_41')
// (9, 2, 'sp4_v_b_15')
// (9, 3, 'local_g0_3')
// (9, 3, 'lutff_4/in_3')
// (9, 3, 'sp4_h_l_39')
// (9, 3, 'sp4_h_l_40')
// (9, 3, 'sp4_h_l_43')
// (9, 3, 'sp4_h_r_10')
// (9, 3, 'sp4_h_r_2')
// (9, 3, 'sp4_r_v_b_27')
// (9, 3, 'sp4_r_v_b_28')
// (9, 3, 'sp4_v_b_2')
// (9, 3, 'sp4_v_t_39')
// (9, 4, 'sp4_r_v_b_14')
// (9, 4, 'sp4_r_v_b_17')
// (9, 4, 'sp4_v_b_39')
// (9, 5, 'sp4_r_v_b_3')
// (9, 5, 'sp4_r_v_b_4')
// (9, 5, 'sp4_v_b_26')
// (9, 6, 'sp12_h_r_9')
// (9, 6, 'sp4_r_v_b_41')
// (9, 6, 'sp4_v_b_15')
// (9, 7, 'sp4_h_r_40')
// (9, 7, 'sp4_r_v_b_28')
// (9, 7, 'sp4_v_b_2')
// (9, 7, 'sp4_v_t_40')
// (9, 8, 'sp4_r_v_b_17')
// (9, 8, 'sp4_v_b_40')
// (9, 9, 'sp4_r_v_b_4')
// (9, 9, 'sp4_v_b_29')
// (9, 10, 'sp4_r_v_b_41')
// (9, 10, 'sp4_v_b_16')
// (9, 11, 'sp4_r_v_b_28')
// (9, 11, 'sp4_v_b_5')
// (9, 11, 'sp4_v_t_40')
// (9, 12, 'sp4_r_v_b_17')
// (9, 12, 'sp4_v_b_40')
// (9, 13, 'sp4_r_v_b_4')
// (9, 13, 'sp4_v_b_29')
// (9, 14, 'local_g1_0')
// (9, 14, 'lutff_7/in_2')
// (9, 14, 'sp4_r_v_b_37')
// (9, 14, 'sp4_v_b_16')
// (9, 15, 'sp4_r_v_b_24')
// (9, 15, 'sp4_v_b_5')
// (9, 16, 'sp4_r_v_b_13')
// (9, 17, 'sp4_r_v_b_0')
// (9, 18, 'sp12_h_r_9')
// (9, 18, 'sp4_r_v_b_37')
// (9, 19, 'sp4_r_v_b_24')
// (9, 20, 'sp4_r_v_b_13')
// (9, 21, 'sp4_r_v_b_0')
// (10, 1, 'local_g0_2')
// (10, 1, 'lutff_5/in_1')
// (10, 1, 'sp12_h_r_5')
// (10, 1, 'sp4_h_l_43')
// (10, 1, 'sp4_h_r_10')
// (10, 1, 'sp4_h_r_12')
// (10, 1, 'sp4_h_r_3')
// (10, 1, 'sp4_v_t_38')
// (10, 1, 'sp4_v_t_41')
// (10, 2, 'sp4_v_b_38')
// (10, 2, 'sp4_v_b_41')
// (10, 3, 'sp4_h_r_15')
// (10, 3, 'sp4_h_r_23')
// (10, 3, 'sp4_v_b_27')
// (10, 3, 'sp4_v_b_28')
// (10, 4, 'sp4_v_b_14')
// (10, 4, 'sp4_v_b_17')
// (10, 5, 'local_g0_3')
// (10, 5, 'lutff_4/in_3')
// (10, 5, 'sp4_v_b_3')
// (10, 5, 'sp4_v_b_4')
// (10, 5, 'sp4_v_t_41')
// (10, 6, 'sp12_h_r_10')
// (10, 6, 'sp4_r_v_b_42')
// (10, 6, 'sp4_v_b_41')
// (10, 7, 'sp4_h_l_40')
// (10, 7, 'sp4_h_r_2')
// (10, 7, 'sp4_r_v_b_31')
// (10, 7, 'sp4_v_b_28')
// (10, 8, 'sp4_r_v_b_18')
// (10, 8, 'sp4_v_b_17')
// (10, 9, 'sp4_r_v_b_7')
// (10, 9, 'sp4_v_b_4')
// (10, 9, 'sp4_v_t_41')
// (10, 10, 'sp4_r_v_b_42')
// (10, 10, 'sp4_v_b_41')
// (10, 11, 'sp4_r_v_b_31')
// (10, 11, 'sp4_v_b_28')
// (10, 12, 'sp4_r_v_b_18')
// (10, 12, 'sp4_v_b_17')
// (10, 13, 'sp4_r_v_b_7')
// (10, 13, 'sp4_v_b_4')
// (10, 13, 'sp4_v_t_37')
// (10, 14, 'sp4_v_b_37')
// (10, 15, 'sp4_v_b_24')
// (10, 16, 'sp4_v_b_13')
// (10, 17, 'local_g0_0')
// (10, 17, 'lutff_1/in_1')
// (10, 17, 'sp4_v_b_0')
// (10, 17, 'sp4_v_t_37')
// (10, 18, 'local_g1_2')
// (10, 18, 'lutff_1/in_2')
// (10, 18, 'sp12_h_r_10')
// (10, 18, 'sp4_v_b_37')
// (10, 19, 'sp4_v_b_24')
// (10, 20, 'local_g1_5')
// (10, 20, 'lutff_6/in_0')
// (10, 20, 'sp4_v_b_13')
// (10, 21, 'sp4_v_b_0')
// (11, 1, 'sp12_h_r_6')
// (11, 1, 'sp4_h_r_14')
// (11, 1, 'sp4_h_r_23')
// (11, 1, 'sp4_h_r_25')
// (11, 3, 'sp4_h_r_26')
// (11, 3, 'sp4_h_r_34')
// (11, 5, 'sp4_h_r_7')
// (11, 5, 'sp4_v_t_42')
// (11, 6, 'sp12_h_r_13')
// (11, 6, 'sp4_v_b_42')
// (11, 7, 'sp4_h_r_15')
// (11, 7, 'sp4_v_b_31')
// (11, 8, 'sp4_v_b_18')
// (11, 9, 'sp4_v_b_7')
// (11, 9, 'sp4_v_t_42')
// (11, 10, 'sp4_v_b_42')
// (11, 11, 'sp4_v_b_31')
// (11, 12, 'sp4_v_b_18')
// (11, 13, 'local_g1_7')
// (11, 13, 'lutff_4/in_2')
// (11, 13, 'sp4_v_b_7')
// (11, 18, 'sp12_h_r_13')
// (12, 1, 'sp12_h_r_9')
// (12, 1, 'sp4_h_r_27')
// (12, 1, 'sp4_h_r_34')
// (12, 1, 'sp4_h_r_36')
// (12, 3, 'sp4_h_r_39')
// (12, 3, 'sp4_h_r_47')
// (12, 5, 'local_g1_2')
// (12, 5, 'lutff_3/in_0')
// (12, 5, 'sp4_h_r_18')
// (12, 5, 'sp4_r_v_b_42')
// (12, 6, 'sp12_h_r_14')
// (12, 6, 'sp4_r_v_b_31')
// (12, 7, 'sp4_h_r_26')
// (12, 7, 'sp4_r_v_b_18')
// (12, 8, 'local_g1_7')
// (12, 8, 'lutff_2/in_2')
// (12, 8, 'sp4_r_v_b_7')
// (12, 14, 'sp4_r_v_b_41')
// (12, 15, 'sp4_r_v_b_28')
// (12, 16, 'sp4_r_v_b_17')
// (12, 17, 'sp4_r_v_b_4')
// (12, 18, 'sp12_h_r_14')
// (12, 18, 'sp4_r_v_b_37')
// (12, 19, 'sp4_r_v_b_24')
// (12, 20, 'sp4_r_v_b_13')
// (12, 21, 'local_g1_0')
// (12, 21, 'lutff_5/in_2')
// (12, 21, 'sp4_r_v_b_0')
// (13, 1, 'sp12_h_r_10')
// (13, 1, 'sp4_h_l_36')
// (13, 1, 'sp4_h_r_10')
// (13, 1, 'sp4_h_r_38')
// (13, 1, 'sp4_h_r_47')
// (13, 3, 'sp4_h_l_39')
// (13, 3, 'sp4_h_l_47')
// (13, 3, 'sp4_h_r_2')
// (13, 4, 'sp4_h_r_7')
// (13, 4, 'sp4_v_t_42')
// (13, 5, 'sp4_h_r_31')
// (13, 5, 'sp4_r_v_b_37')
// (13, 5, 'sp4_v_b_42')
// (13, 6, 'sp12_h_r_17')
// (13, 6, 'sp4_r_v_b_24')
// (13, 6, 'sp4_v_b_31')
// (13, 7, 'sp4_h_r_39')
// (13, 7, 'sp4_r_v_b_13')
// (13, 7, 'sp4_v_b_18')
// (13, 8, 'sp4_r_v_b_0')
// (13, 8, 'sp4_v_b_7')
// (13, 13, 'sp4_h_r_10')
// (13, 13, 'sp4_v_t_41')
// (13, 14, 'sp4_v_b_41')
// (13, 15, 'sp4_v_b_28')
// (13, 16, 'sp4_v_b_17')
// (13, 17, 'sp4_v_b_4')
// (13, 17, 'sp4_v_t_37')
// (13, 18, 'sp12_h_r_17')
// (13, 18, 'sp4_v_b_37')
// (13, 19, 'sp4_v_b_24')
// (13, 20, 'sp4_v_b_13')
// (13, 21, 'sp4_v_b_0')
// (14, 1, 'sp12_h_r_13')
// (14, 1, 'sp4_h_l_38')
// (14, 1, 'sp4_h_l_47')
// (14, 1, 'sp4_h_r_23')
// (14, 1, 'sp4_h_r_7')
// (14, 2, 'local_g2_7')
// (14, 2, 'lutff_3/in_2')
// (14, 2, 'sp4_r_v_b_39')
// (14, 3, 'sp4_h_r_15')
// (14, 3, 'sp4_r_v_b_26')
// (14, 4, 'sp4_h_r_18')
// (14, 4, 'sp4_h_r_6')
// (14, 4, 'sp4_r_v_b_15')
// (14, 4, 'sp4_v_t_37')
// (14, 5, 'local_g1_2')
// (14, 5, 'lutff_7/in_2')
// (14, 5, 'sp4_h_r_42')
// (14, 5, 'sp4_r_v_b_2')
// (14, 5, 'sp4_v_b_37')
// (14, 6, 'sp12_h_r_18')
// (14, 6, 'sp4_v_b_24')
// (14, 7, 'local_g1_5')
// (14, 7, 'lutff_4/in_2')
// (14, 7, 'sp4_h_l_39')
// (14, 7, 'sp4_h_r_11')
// (14, 7, 'sp4_v_b_13')
// (14, 8, 'sp4_v_b_0')
// (14, 13, 'sp4_h_r_23')
// (14, 18, 'sp12_h_r_18')
// (15, 1, 'sp12_h_r_14')
// (15, 1, 'sp4_h_r_18')
// (15, 1, 'sp4_h_r_2')
// (15, 1, 'sp4_h_r_34')
// (15, 1, 'sp4_v_t_39')
// (15, 2, 'sp4_v_b_39')
// (15, 3, 'sp4_h_r_26')
// (15, 3, 'sp4_v_b_26')
// (15, 4, 'local_g2_7')
// (15, 4, 'lutff_3/in_2')
// (15, 4, 'sp4_h_r_19')
// (15, 4, 'sp4_h_r_31')
// (15, 4, 'sp4_v_b_15')
// (15, 5, 'sp4_h_l_42')
// (15, 5, 'sp4_v_b_2')
// (15, 6, 'sp12_h_r_21')
// (15, 7, 'sp4_h_r_22')
// (15, 13, 'sp4_h_r_34')
// (15, 18, 'sp12_h_r_21')
// (16, 0, 'logic_op_tnr_5')
// (16, 1, 'neigh_op_rgt_5')
// (16, 1, 'sp12_h_r_17')
// (16, 1, 'sp4_h_r_15')
// (16, 1, 'sp4_h_r_31')
// (16, 1, 'sp4_h_r_47')
// (16, 1, 'sp4_r_v_b_10')
// (16, 1, 'sp4_r_v_b_26')
// (16, 1, 'sp4_r_v_b_42')
// (16, 2, 'local_g0_5')
// (16, 2, 'lutff_7/in_0')
// (16, 2, 'neigh_op_bnr_5')
// (16, 2, 'sp4_r_v_b_15')
// (16, 2, 'sp4_r_v_b_31')
// (16, 2, 'sp4_r_v_b_47')
// (16, 3, 'local_g1_2')
// (16, 3, 'lutff_6/in_3')
// (16, 3, 'sp4_h_r_39')
// (16, 3, 'sp4_r_v_b_18')
// (16, 3, 'sp4_r_v_b_2')
// (16, 3, 'sp4_r_v_b_34')
// (16, 4, 'sp4_h_r_30')
// (16, 4, 'sp4_h_r_42')
// (16, 4, 'sp4_r_v_b_23')
// (16, 4, 'sp4_r_v_b_7')
// (16, 5, 'local_g2_2')
// (16, 5, 'lutff_2/in_0')
// (16, 5, 'sp4_r_v_b_10')
// (16, 6, 'sp12_h_r_22')
// (16, 6, 'sp4_r_v_b_47')
// (16, 7, 'sp4_h_r_35')
// (16, 7, 'sp4_r_v_b_34')
// (16, 8, 'sp4_r_v_b_23')
// (16, 9, 'sp4_r_v_b_10')
// (16, 10, 'sp4_r_v_b_47')
// (16, 11, 'sp4_r_v_b_34')
// (16, 12, 'sp4_r_v_b_23')
// (16, 13, 'sp4_h_r_47')
// (16, 13, 'sp4_r_v_b_10')
// (16, 18, 'sp12_h_r_22')
// (17, 0, 'logic_op_top_5')
// (17, 0, 'span12_vert_10')
// (17, 0, 'span4_vert_10')
// (17, 0, 'span4_vert_26')
// (17, 0, 'span4_vert_42')
// (17, 1, 'lutff_5/out')
// (17, 1, 'sp12_h_r_18')
// (17, 1, 'sp12_v_b_10')
// (17, 1, 'sp4_h_l_47')
// (17, 1, 'sp4_h_r_26')
// (17, 1, 'sp4_h_r_42')
// (17, 1, 'sp4_r_v_b_27')
// (17, 1, 'sp4_r_v_b_43')
// (17, 1, 'sp4_v_b_10')
// (17, 1, 'sp4_v_b_26')
// (17, 1, 'sp4_v_b_42')
// (17, 1, 'sp4_v_t_47')
// (17, 2, 'neigh_op_bot_5')
// (17, 2, 'sp12_v_b_9')
// (17, 2, 'sp4_r_v_b_14')
// (17, 2, 'sp4_r_v_b_30')
// (17, 2, 'sp4_v_b_15')
// (17, 2, 'sp4_v_b_31')
// (17, 2, 'sp4_v_b_47')
// (17, 3, 'sp12_v_b_6')
// (17, 3, 'sp4_h_l_39')
// (17, 3, 'sp4_r_v_b_19')
// (17, 3, 'sp4_r_v_b_3')
// (17, 3, 'sp4_v_b_18')
// (17, 3, 'sp4_v_b_2')
// (17, 3, 'sp4_v_b_34')
// (17, 4, 'sp12_v_b_5')
// (17, 4, 'sp4_h_l_42')
// (17, 4, 'sp4_h_r_43')
// (17, 4, 'sp4_r_v_b_46')
// (17, 4, 'sp4_r_v_b_6')
// (17, 4, 'sp4_v_b_23')
// (17, 4, 'sp4_v_b_7')
// (17, 5, 'sp12_v_b_2')
// (17, 5, 'sp4_r_v_b_35')
// (17, 5, 'sp4_v_b_10')
// (17, 5, 'sp4_v_t_47')
// (17, 6, 'sp12_h_l_22')
// (17, 6, 'sp12_v_b_1')
// (17, 6, 'sp12_v_t_22')
// (17, 6, 'sp4_r_v_b_22')
// (17, 6, 'sp4_v_b_47')
// (17, 7, 'sp12_v_b_22')
// (17, 7, 'sp4_h_r_46')
// (17, 7, 'sp4_r_v_b_11')
// (17, 7, 'sp4_v_b_34')
// (17, 8, 'sp12_v_b_21')
// (17, 8, 'sp4_v_b_23')
// (17, 9, 'sp12_v_b_18')
// (17, 9, 'sp4_v_b_10')
// (17, 9, 'sp4_v_t_47')
// (17, 10, 'sp12_v_b_17')
// (17, 10, 'sp4_v_b_47')
// (17, 11, 'sp12_v_b_14')
// (17, 11, 'sp4_v_b_34')
// (17, 12, 'sp12_v_b_13')
// (17, 12, 'sp4_v_b_23')
// (17, 13, 'sp12_v_b_10')
// (17, 13, 'sp4_h_l_47')
// (17, 13, 'sp4_v_b_10')
// (17, 14, 'sp12_v_b_9')
// (17, 15, 'sp12_v_b_6')
// (17, 16, 'sp12_v_b_5')
// (17, 17, 'sp12_v_b_2')
// (17, 18, 'sp12_h_l_22')
// (17, 18, 'sp12_v_b_1')
// (18, 0, 'logic_op_tnl_5')
// (18, 0, 'span4_vert_27')
// (18, 0, 'span4_vert_43')
// (18, 1, 'neigh_op_lft_5')
// (18, 1, 'sp12_h_r_21')
// (18, 1, 'sp4_h_l_42')
// (18, 1, 'sp4_h_r_39')
// (18, 1, 'sp4_v_b_27')
// (18, 1, 'sp4_v_b_43')
// (18, 2, 'neigh_op_bnl_5')
// (18, 2, 'sp4_v_b_14')
// (18, 2, 'sp4_v_b_30')
// (18, 3, 'sp4_v_b_19')
// (18, 3, 'sp4_v_b_3')
// (18, 3, 'sp4_v_t_46')
// (18, 4, 'sp4_h_l_43')
// (18, 4, 'sp4_v_b_46')
// (18, 4, 'sp4_v_b_6')
// (18, 5, 'sp4_v_b_35')
// (18, 6, 'sp4_v_b_22')
// (18, 7, 'sp4_h_l_46')
// (18, 7, 'sp4_v_b_11')
// (19, 1, 'sp12_h_r_22')
// (19, 1, 'sp4_h_l_39')
// (20, 1, 'sp12_h_l_22')

wire n190;
// (1, 3, 'local_g2_2')
// (1, 3, 'lutff_1/in_1')
// (1, 3, 'neigh_op_tnr_2')
// (1, 4, 'neigh_op_rgt_2')
// (1, 5, 'neigh_op_bnr_2')
// (2, 3, 'neigh_op_top_2')
// (2, 4, 'lutff_2/out')
// (2, 5, 'neigh_op_bot_2')
// (3, 3, 'neigh_op_tnl_2')
// (3, 4, 'neigh_op_lft_2')
// (3, 5, 'neigh_op_bnl_2')

reg n191 = 0;
// (1, 3, 'local_g2_6')
// (1, 3, 'lutff_2/in_0')
// (1, 3, 'neigh_op_tnr_6')
// (1, 4, 'neigh_op_rgt_6')
// (1, 5, 'neigh_op_bnr_6')
// (2, 3, 'neigh_op_top_6')
// (2, 4, 'lutff_6/out')
// (2, 5, 'local_g0_6')
// (2, 5, 'lutff_5/in_3')
// (2, 5, 'lutff_6/in_2')
// (2, 5, 'neigh_op_bot_6')
// (3, 3, 'neigh_op_tnl_6')
// (3, 4, 'neigh_op_lft_6')
// (3, 5, 'neigh_op_bnl_6')

reg n192 = 0;
// (1, 3, 'neigh_op_tnr_0')
// (1, 4, 'neigh_op_rgt_0')
// (1, 5, 'neigh_op_bnr_0')
// (2, 3, 'local_g1_0')
// (2, 3, 'lutff_2/in_1')
// (2, 3, 'neigh_op_top_0')
// (2, 4, 'local_g2_0')
// (2, 4, 'lutff_0/out')
// (2, 4, 'lutff_1/in_3')
// (2, 5, 'neigh_op_bot_0')
// (3, 3, 'neigh_op_tnl_0')
// (3, 4, 'local_g1_0')
// (3, 4, 'lutff_5/in_0')
// (3, 4, 'neigh_op_lft_0')
// (3, 5, 'neigh_op_bnl_0')

reg n193 = 0;
// (1, 3, 'neigh_op_tnr_1')
// (1, 4, 'neigh_op_rgt_1')
// (1, 5, 'neigh_op_bnr_1')
// (2, 3, 'local_g1_1')
// (2, 3, 'lutff_5/in_3')
// (2, 3, 'neigh_op_top_1')
// (2, 4, 'local_g0_1')
// (2, 4, 'lutff_1/out')
// (2, 4, 'lutff_3/in_0')
// (2, 4, 'lutff_7/in_2')
// (2, 5, 'neigh_op_bot_1')
// (3, 3, 'neigh_op_tnl_1')
// (3, 4, 'neigh_op_lft_1')
// (3, 5, 'neigh_op_bnl_1')

reg n194 = 0;
// (1, 3, 'neigh_op_tnr_3')
// (1, 4, 'neigh_op_rgt_3')
// (1, 5, 'neigh_op_bnr_3')
// (2, 3, 'neigh_op_top_3')
// (2, 4, 'local_g3_3')
// (2, 4, 'lutff_2/in_0')
// (2, 4, 'lutff_3/out')
// (2, 4, 'lutff_6/in_2')
// (2, 5, 'local_g1_3')
// (2, 5, 'lutff_3/in_1')
// (2, 5, 'neigh_op_bot_3')
// (3, 3, 'neigh_op_tnl_3')
// (3, 4, 'neigh_op_lft_3')
// (3, 5, 'neigh_op_bnl_3')

reg n195 = 0;
// (1, 3, 'neigh_op_tnr_4')
// (1, 4, 'neigh_op_rgt_4')
// (1, 5, 'neigh_op_bnr_4')
// (2, 3, 'local_g1_4')
// (2, 3, 'lutff_2/in_3')
// (2, 3, 'neigh_op_top_4')
// (2, 4, 'local_g0_4')
// (2, 4, 'lutff_0/in_2')
// (2, 4, 'lutff_4/out')
// (2, 5, 'neigh_op_bot_4')
// (3, 3, 'neigh_op_tnl_4')
// (3, 4, 'local_g1_4')
// (3, 4, 'lutff_5/in_2')
// (3, 4, 'neigh_op_lft_4')
// (3, 5, 'neigh_op_bnl_4')

wire n196;
// (1, 3, 'neigh_op_tnr_5')
// (1, 4, 'neigh_op_rgt_5')
// (1, 5, 'neigh_op_bnr_5')
// (2, 3, 'neigh_op_top_5')
// (2, 4, 'lutff_5/out')
// (2, 5, 'local_g1_5')
// (2, 5, 'lutff_0/in_2')
// (2, 5, 'neigh_op_bot_5')
// (3, 3, 'neigh_op_tnl_5')
// (3, 4, 'neigh_op_lft_5')
// (3, 5, 'neigh_op_bnl_5')

wire n197;
// (1, 3, 'neigh_op_tnr_7')
// (1, 4, 'neigh_op_rgt_7')
// (1, 5, 'neigh_op_bnr_7')
// (2, 3, 'neigh_op_top_7')
// (2, 4, 'lutff_7/out')
// (2, 5, 'neigh_op_bot_7')
// (3, 3, 'neigh_op_tnl_7')
// (3, 4, 'local_g0_7')
// (3, 4, 'lutff_4/in_1')
// (3, 4, 'neigh_op_lft_7')
// (3, 5, 'neigh_op_bnl_7')

wire n198;
// (1, 3, 'sp4_h_r_3')
// (2, 3, 'sp4_h_r_14')
// (3, 2, 'sp4_r_v_b_43')
// (3, 3, 'local_g3_3')
// (3, 3, 'lutff_global/cen')
// (3, 3, 'sp4_h_r_27')
// (3, 3, 'sp4_r_v_b_30')
// (3, 4, 'sp4_r_v_b_19')
// (3, 5, 'sp4_r_v_b_6')
// (4, 1, 'sp4_v_t_43')
// (4, 2, 'sp4_v_b_43')
// (4, 3, 'sp4_h_r_38')
// (4, 3, 'sp4_v_b_30')
// (4, 4, 'local_g1_3')
// (4, 4, 'lutff_global/cen')
// (4, 4, 'sp4_v_b_19')
// (4, 5, 'sp4_h_r_6')
// (4, 5, 'sp4_v_b_6')
// (5, 2, 'sp4_r_v_b_39')
// (5, 3, 'local_g0_2')
// (5, 3, 'lutff_global/cen')
// (5, 3, 'sp4_h_l_38')
// (5, 3, 'sp4_h_r_3')
// (5, 3, 'sp4_r_v_b_26')
// (5, 4, 'sp4_r_v_b_15')
// (5, 5, 'sp4_h_r_19')
// (5, 5, 'sp4_r_v_b_2')
// (6, 1, 'sp4_v_t_39')
// (6, 2, 'sp4_v_b_39')
// (6, 3, 'sp4_h_r_14')
// (6, 3, 'sp4_v_b_26')
// (6, 4, 'sp4_v_b_15')
// (6, 5, 'sp4_h_r_2')
// (6, 5, 'sp4_h_r_30')
// (6, 5, 'sp4_v_b_2')
// (7, 3, 'sp4_h_r_27')
// (7, 4, 'neigh_op_tnr_5')
// (7, 5, 'neigh_op_rgt_5')
// (7, 5, 'sp4_h_r_15')
// (7, 5, 'sp4_h_r_43')
// (7, 6, 'neigh_op_bnr_5')
// (8, 3, 'sp4_h_r_38')
// (8, 4, 'neigh_op_top_5')
// (8, 4, 'sp4_r_v_b_38')
// (8, 5, 'lutff_5/out')
// (8, 5, 'sp4_h_l_43')
// (8, 5, 'sp4_h_r_10')
// (8, 5, 'sp4_h_r_26')
// (8, 5, 'sp4_r_v_b_27')
// (8, 6, 'neigh_op_bot_5')
// (8, 6, 'sp4_r_v_b_14')
// (8, 7, 'sp4_r_v_b_3')
// (9, 3, 'sp4_h_l_38')
// (9, 3, 'sp4_v_t_38')
// (9, 4, 'neigh_op_tnl_5')
// (9, 4, 'sp4_v_b_38')
// (9, 5, 'neigh_op_lft_5')
// (9, 5, 'sp4_h_r_23')
// (9, 5, 'sp4_h_r_39')
// (9, 5, 'sp4_v_b_27')
// (9, 6, 'neigh_op_bnl_5')
// (9, 6, 'sp4_v_b_14')
// (9, 7, 'sp4_v_b_3')
// (10, 5, 'sp4_h_l_39')
// (10, 5, 'sp4_h_r_34')
// (11, 5, 'sp4_h_r_47')
// (12, 5, 'sp4_h_l_47')

reg n199 = 0;
// (1, 3, 'sp4_r_v_b_36')
// (1, 4, 'sp4_r_v_b_25')
// (1, 5, 'sp4_r_v_b_12')
// (1, 6, 'sp4_r_v_b_1')
// (1, 7, 'sp4_r_v_b_47')
// (1, 8, 'sp4_r_v_b_34')
// (1, 9, 'neigh_op_tnr_5')
// (1, 9, 'sp4_r_v_b_23')
// (1, 10, 'neigh_op_rgt_5')
// (1, 10, 'sp4_r_v_b_10')
// (1, 10, 'sp4_r_v_b_42')
// (1, 11, 'neigh_op_bnr_5')
// (1, 11, 'sp4_r_v_b_31')
// (1, 12, 'sp4_r_v_b_18')
// (1, 13, 'sp4_r_v_b_7')
// (1, 14, 'sp4_r_v_b_42')
// (1, 15, 'sp4_r_v_b_31')
// (1, 16, 'sp4_r_v_b_18')
// (1, 17, 'sp4_r_v_b_7')
// (2, 2, 'sp4_v_t_36')
// (2, 3, 'sp4_r_v_b_39')
// (2, 3, 'sp4_v_b_36')
// (2, 4, 'sp4_r_v_b_26')
// (2, 4, 'sp4_v_b_25')
// (2, 5, 'local_g1_4')
// (2, 5, 'lutff_0/in_3')
// (2, 5, 'sp4_r_v_b_15')
// (2, 5, 'sp4_v_b_12')
// (2, 6, 'sp4_r_v_b_2')
// (2, 6, 'sp4_v_b_1')
// (2, 6, 'sp4_v_t_47')
// (2, 7, 'sp4_r_v_b_46')
// (2, 7, 'sp4_v_b_47')
// (2, 8, 'sp4_r_v_b_35')
// (2, 8, 'sp4_v_b_34')
// (2, 9, 'neigh_op_top_5')
// (2, 9, 'sp4_r_v_b_22')
// (2, 9, 'sp4_v_b_23')
// (2, 9, 'sp4_v_t_42')
// (2, 10, 'local_g0_5')
// (2, 10, 'lutff_5/in_0')
// (2, 10, 'lutff_5/out')
// (2, 10, 'sp4_r_v_b_11')
// (2, 10, 'sp4_v_b_10')
// (2, 10, 'sp4_v_b_42')
// (2, 11, 'neigh_op_bot_5')
// (2, 11, 'sp4_v_b_31')
// (2, 12, 'sp4_v_b_18')
// (2, 13, 'sp4_v_b_7')
// (2, 13, 'sp4_v_t_42')
// (2, 14, 'sp4_v_b_42')
// (2, 15, 'local_g2_7')
// (2, 15, 'lutff_2/in_1')
// (2, 15, 'sp4_v_b_31')
// (2, 16, 'sp4_v_b_18')
// (2, 17, 'sp4_v_b_7')
// (3, 2, 'sp4_v_t_39')
// (3, 3, 'sp4_v_b_39')
// (3, 4, 'local_g2_2')
// (3, 4, 'lutff_3/in_1')
// (3, 4, 'sp4_v_b_26')
// (3, 5, 'sp4_v_b_15')
// (3, 6, 'sp4_v_b_2')
// (3, 6, 'sp4_v_t_46')
// (3, 7, 'sp4_v_b_46')
// (3, 8, 'sp4_v_b_35')
// (3, 9, 'neigh_op_tnl_5')
// (3, 9, 'sp4_v_b_22')
// (3, 10, 'neigh_op_lft_5')
// (3, 10, 'sp4_v_b_11')
// (3, 11, 'local_g3_5')
// (3, 11, 'lutff_0/in_2')
// (3, 11, 'neigh_op_bnl_5')

reg n200 = 0;
// (1, 3, 'sp4_r_v_b_43')
// (1, 4, 'sp4_r_v_b_30')
// (1, 4, 'sp4_r_v_b_46')
// (1, 5, 'neigh_op_tnr_3')
// (1, 5, 'sp4_r_v_b_19')
// (1, 5, 'sp4_r_v_b_35')
// (1, 6, 'neigh_op_rgt_3')
// (1, 6, 'sp4_h_r_11')
// (1, 6, 'sp4_r_v_b_22')
// (1, 6, 'sp4_r_v_b_6')
// (1, 7, 'neigh_op_bnr_3')
// (1, 7, 'sp4_r_v_b_11')
// (2, 2, 'local_g0_3')
// (2, 2, 'lutff_1/in_0')
// (2, 2, 'sp4_h_r_11')
// (2, 2, 'sp4_v_t_43')
// (2, 3, 'sp4_h_r_4')
// (2, 3, 'sp4_r_v_b_42')
// (2, 3, 'sp4_v_b_43')
// (2, 3, 'sp4_v_t_46')
// (2, 4, 'sp4_r_v_b_31')
// (2, 4, 'sp4_r_v_b_47')
// (2, 4, 'sp4_v_b_30')
// (2, 4, 'sp4_v_b_46')
// (2, 5, 'neigh_op_top_3')
// (2, 5, 'sp4_r_v_b_18')
// (2, 5, 'sp4_r_v_b_34')
// (2, 5, 'sp4_v_b_19')
// (2, 5, 'sp4_v_b_35')
// (2, 6, 'local_g1_3')
// (2, 6, 'lutff_3/in_1')
// (2, 6, 'lutff_3/out')
// (2, 6, 'lutff_6/in_2')
// (2, 6, 'lutff_7/in_3')
// (2, 6, 'sp4_h_r_22')
// (2, 6, 'sp4_r_v_b_23')
// (2, 6, 'sp4_r_v_b_7')
// (2, 6, 'sp4_v_b_22')
// (2, 6, 'sp4_v_b_6')
// (2, 7, 'neigh_op_bot_3')
// (2, 7, 'sp4_r_v_b_10')
// (2, 7, 'sp4_v_b_11')
// (3, 2, 'sp4_h_r_0')
// (3, 2, 'sp4_h_r_22')
// (3, 2, 'sp4_h_r_7')
// (3, 2, 'sp4_v_t_42')
// (3, 3, 'sp4_h_r_17')
// (3, 3, 'sp4_h_r_3')
// (3, 3, 'sp4_v_b_42')
// (3, 3, 'sp4_v_t_47')
// (3, 4, 'local_g3_7')
// (3, 4, 'lutff_4/in_2')
// (3, 4, 'sp4_v_b_31')
// (3, 4, 'sp4_v_b_47')
// (3, 5, 'local_g2_3')
// (3, 5, 'lutff_2/in_1')
// (3, 5, 'lutff_4/in_3')
// (3, 5, 'neigh_op_tnl_3')
// (3, 5, 'sp4_v_b_18')
// (3, 5, 'sp4_v_b_34')
// (3, 6, 'local_g1_3')
// (3, 6, 'lutff_0/in_0')
// (3, 6, 'neigh_op_lft_3')
// (3, 6, 'sp4_h_r_35')
// (3, 6, 'sp4_v_b_23')
// (3, 6, 'sp4_v_b_7')
// (3, 7, 'neigh_op_bnl_3')
// (3, 7, 'sp4_h_r_4')
// (3, 7, 'sp4_v_b_10')
// (4, 1, 'local_g3_5')
// (4, 1, 'lutff_1/in_1')
// (4, 1, 'sp4_r_v_b_21')
// (4, 2, 'sp4_h_r_13')
// (4, 2, 'sp4_h_r_18')
// (4, 2, 'sp4_h_r_35')
// (4, 2, 'sp4_r_v_b_8')
// (4, 3, 'local_g2_4')
// (4, 3, 'lutff_2/in_0')
// (4, 3, 'sp4_h_r_14')
// (4, 3, 'sp4_h_r_28')
// (4, 3, 'sp4_r_v_b_40')
// (4, 3, 'sp4_r_v_b_46')
// (4, 4, 'local_g2_3')
// (4, 4, 'lutff_2/in_3')
// (4, 4, 'sp4_r_v_b_29')
// (4, 4, 'sp4_r_v_b_35')
// (4, 5, 'sp4_r_v_b_16')
// (4, 5, 'sp4_r_v_b_22')
// (4, 6, 'sp4_h_r_46')
// (4, 6, 'sp4_r_v_b_11')
// (4, 6, 'sp4_r_v_b_5')
// (4, 7, 'local_g1_1')
// (4, 7, 'lutff_4/in_2')
// (4, 7, 'lutff_5/in_1')
// (4, 7, 'sp4_h_r_17')
// (4, 7, 'sp4_r_v_b_46')
// (4, 8, 'local_g2_3')
// (4, 8, 'lutff_5/in_2')
// (4, 8, 'sp4_r_v_b_35')
// (4, 9, 'sp4_r_v_b_22')
// (4, 10, 'sp4_r_v_b_11')
// (5, 0, 'span4_vert_21')
// (5, 1, 'local_g3_0')
// (5, 1, 'lutff_5/in_0')
// (5, 1, 'sp4_r_v_b_16')
// (5, 1, 'sp4_v_b_21')
// (5, 2, 'sp4_h_r_10')
// (5, 2, 'sp4_h_r_24')
// (5, 2, 'sp4_h_r_31')
// (5, 2, 'sp4_h_r_46')
// (5, 2, 'sp4_r_v_b_5')
// (5, 2, 'sp4_v_b_8')
// (5, 2, 'sp4_v_t_40')
// (5, 2, 'sp4_v_t_46')
// (5, 3, 'local_g2_3')
// (5, 3, 'lutff_6/in_1')
// (5, 3, 'sp4_h_r_27')
// (5, 3, 'sp4_h_r_41')
// (5, 3, 'sp4_v_b_40')
// (5, 3, 'sp4_v_b_46')
// (5, 4, 'sp4_v_b_29')
// (5, 4, 'sp4_v_b_35')
// (5, 5, 'sp4_v_b_16')
// (5, 5, 'sp4_v_b_22')
// (5, 6, 'sp4_h_l_46')
// (5, 6, 'sp4_v_b_11')
// (5, 6, 'sp4_v_b_5')
// (5, 6, 'sp4_v_t_46')
// (5, 7, 'local_g3_4')
// (5, 7, 'lutff_2/in_1')
// (5, 7, 'sp4_h_r_28')
// (5, 7, 'sp4_v_b_46')
// (5, 8, 'sp4_v_b_35')
// (5, 9, 'sp4_v_b_22')
// (5, 10, 'sp4_v_b_11')
// (6, 0, 'span4_vert_16')
// (6, 1, 'sp4_v_b_16')
// (6, 2, 'sp4_h_l_46')
// (6, 2, 'sp4_h_r_23')
// (6, 2, 'sp4_h_r_37')
// (6, 2, 'sp4_h_r_42')
// (6, 2, 'sp4_h_r_7')
// (6, 2, 'sp4_v_b_5')
// (6, 3, 'sp4_h_l_41')
// (6, 3, 'sp4_h_r_38')
// (6, 7, 'sp4_h_r_41')
// (7, 2, 'local_g0_0')
// (7, 2, 'lutff_1/in_1')
// (7, 2, 'lutff_4/in_2')
// (7, 2, 'lutff_5/in_1')
// (7, 2, 'sp4_h_l_37')
// (7, 2, 'sp4_h_l_42')
// (7, 2, 'sp4_h_r_18')
// (7, 2, 'sp4_h_r_34')
// (7, 2, 'sp4_h_r_7')
// (7, 2, 'sp4_h_r_8')
// (7, 3, 'sp4_h_l_38')
// (7, 3, 'sp4_h_r_11')
// (7, 7, 'sp4_h_l_41')
// (8, 1, 'local_g3_7')
// (8, 1, 'lutff_3/in_3')
// (8, 1, 'sp4_r_v_b_23')
// (8, 2, 'local_g1_2')
// (8, 2, 'local_g3_7')
// (8, 2, 'lutff_0/in_3')
// (8, 2, 'lutff_1/in_1')
// (8, 2, 'sp4_h_r_18')
// (8, 2, 'sp4_h_r_21')
// (8, 2, 'sp4_h_r_31')
// (8, 2, 'sp4_h_r_47')
// (8, 2, 'sp4_r_v_b_10')
// (8, 3, 'sp4_h_r_22')
// (9, 0, 'span4_vert_23')
// (9, 1, 'sp4_v_b_23')
// (9, 2, 'sp4_h_l_47')
// (9, 2, 'sp4_h_r_31')
// (9, 2, 'sp4_h_r_32')
// (9, 2, 'sp4_h_r_42')
// (9, 2, 'sp4_v_b_10')
// (9, 3, 'local_g2_3')
// (9, 3, 'lutff_3/in_2')
// (9, 3, 'lutff_6/in_1')
// (9, 3, 'sp4_h_r_35')
// (10, 2, 'sp4_h_l_42')
// (10, 2, 'sp4_h_r_42')
// (10, 2, 'sp4_h_r_45')
// (10, 3, 'sp4_h_r_46')
// (11, 2, 'sp4_h_l_42')
// (11, 2, 'sp4_h_l_45')
// (11, 3, 'sp4_h_l_46')

wire n201;
// (1, 3, 'sp4_r_v_b_47')
// (1, 4, 'local_g2_2')
// (1, 4, 'lutff_global/cen')
// (1, 4, 'sp4_r_v_b_34')
// (1, 4, 'sp4_r_v_b_38')
// (1, 5, 'local_g1_3')
// (1, 5, 'lutff_global/cen')
// (1, 5, 'sp4_r_v_b_23')
// (1, 5, 'sp4_r_v_b_27')
// (1, 6, 'sp4_r_v_b_10')
// (1, 6, 'sp4_r_v_b_14')
// (1, 7, 'sp4_r_v_b_3')
// (1, 7, 'sp4_r_v_b_39')
// (1, 8, 'sp4_r_v_b_26')
// (1, 8, 'sp4_r_v_b_42')
// (1, 9, 'neigh_op_tnr_1')
// (1, 9, 'sp4_r_v_b_15')
// (1, 9, 'sp4_r_v_b_31')
// (1, 10, 'neigh_op_rgt_1')
// (1, 10, 'sp4_r_v_b_18')
// (1, 10, 'sp4_r_v_b_2')
// (1, 11, 'neigh_op_bnr_1')
// (1, 11, 'sp4_r_v_b_7')
// (2, 2, 'sp4_v_t_47')
// (2, 3, 'sp4_r_v_b_43')
// (2, 3, 'sp4_v_b_47')
// (2, 3, 'sp4_v_t_38')
// (2, 4, 'local_g2_2')
// (2, 4, 'lutff_global/cen')
// (2, 4, 'sp4_r_v_b_30')
// (2, 4, 'sp4_v_b_34')
// (2, 4, 'sp4_v_b_38')
// (2, 5, 'local_g3_3')
// (2, 5, 'lutff_global/cen')
// (2, 5, 'sp4_r_v_b_19')
// (2, 5, 'sp4_v_b_23')
// (2, 5, 'sp4_v_b_27')
// (2, 6, 'sp4_r_v_b_6')
// (2, 6, 'sp4_v_b_10')
// (2, 6, 'sp4_v_b_14')
// (2, 6, 'sp4_v_t_39')
// (2, 7, 'sp4_r_v_b_38')
// (2, 7, 'sp4_v_b_3')
// (2, 7, 'sp4_v_b_39')
// (2, 7, 'sp4_v_t_42')
// (2, 8, 'sp4_r_v_b_27')
// (2, 8, 'sp4_v_b_26')
// (2, 8, 'sp4_v_b_42')
// (2, 9, 'neigh_op_top_1')
// (2, 9, 'sp4_r_v_b_14')
// (2, 9, 'sp4_v_b_15')
// (2, 9, 'sp4_v_b_31')
// (2, 10, 'lutff_1/out')
// (2, 10, 'sp4_r_v_b_3')
// (2, 10, 'sp4_v_b_18')
// (2, 10, 'sp4_v_b_2')
// (2, 11, 'neigh_op_bot_1')
// (2, 11, 'sp4_v_b_7')
// (3, 2, 'sp4_v_t_43')
// (3, 3, 'sp4_v_b_43')
// (3, 4, 'sp4_v_b_30')
// (3, 5, 'sp4_v_b_19')
// (3, 6, 'sp4_v_b_6')
// (3, 6, 'sp4_v_t_38')
// (3, 7, 'sp4_v_b_38')
// (3, 8, 'sp4_v_b_27')
// (3, 9, 'neigh_op_tnl_1')
// (3, 9, 'sp4_v_b_14')
// (3, 10, 'neigh_op_lft_1')
// (3, 10, 'sp4_v_b_3')
// (3, 11, 'neigh_op_bnl_1')

wire n202;
// (1, 4, 'neigh_op_tnr_0')
// (1, 5, 'neigh_op_rgt_0')
// (1, 6, 'neigh_op_bnr_0')
// (2, 4, 'neigh_op_top_0')
// (2, 5, 'local_g3_0')
// (2, 5, 'lutff_0/out')
// (2, 5, 'lutff_4/in_3')
// (2, 6, 'neigh_op_bot_0')
// (3, 4, 'neigh_op_tnl_0')
// (3, 5, 'neigh_op_lft_0')
// (3, 6, 'neigh_op_bnl_0')

wire n203;
// (1, 4, 'neigh_op_tnr_2')
// (1, 5, 'neigh_op_rgt_2')
// (1, 6, 'neigh_op_bnr_2')
// (2, 4, 'neigh_op_top_2')
// (2, 5, 'lutff_2/out')
// (2, 6, 'neigh_op_bot_2')
// (3, 4, 'neigh_op_tnl_2')
// (3, 5, 'local_g1_2')
// (3, 5, 'lutff_3/in_2')
// (3, 5, 'neigh_op_lft_2')
// (3, 6, 'neigh_op_bnl_2')

wire n204;
// (1, 4, 'neigh_op_tnr_3')
// (1, 5, 'neigh_op_rgt_3')
// (1, 6, 'neigh_op_bnr_3')
// (2, 4, 'neigh_op_top_3')
// (2, 5, 'lutff_3/out')
// (2, 6, 'neigh_op_bot_3')
// (3, 4, 'neigh_op_tnl_3')
// (3, 5, 'local_g1_3')
// (3, 5, 'lutff_2/in_2')
// (3, 5, 'neigh_op_lft_3')
// (3, 6, 'neigh_op_bnl_3')

wire n205;
// (1, 4, 'neigh_op_tnr_4')
// (1, 5, 'neigh_op_rgt_4')
// (1, 6, 'neigh_op_bnr_4')
// (2, 4, 'neigh_op_top_4')
// (2, 5, 'lutff_4/out')
// (2, 6, 'neigh_op_bot_4')
// (3, 4, 'local_g3_4')
// (3, 4, 'lutff_3/in_0')
// (3, 4, 'neigh_op_tnl_4')
// (3, 5, 'neigh_op_lft_4')
// (3, 6, 'neigh_op_bnl_4')

wire n206;
// (1, 4, 'neigh_op_tnr_5')
// (1, 5, 'neigh_op_rgt_5')
// (1, 6, 'neigh_op_bnr_5')
// (2, 4, 'neigh_op_top_5')
// (2, 5, 'lutff_5/out')
// (2, 6, 'neigh_op_bot_5')
// (3, 4, 'neigh_op_tnl_5')
// (3, 5, 'local_g1_5')
// (3, 5, 'lutff_2/in_0')
// (3, 5, 'neigh_op_lft_5')
// (3, 6, 'neigh_op_bnl_5')

wire n207;
// (1, 4, 'neigh_op_tnr_7')
// (1, 5, 'neigh_op_rgt_7')
// (1, 6, 'neigh_op_bnr_7')
// (2, 4, 'neigh_op_top_7')
// (2, 5, 'lutff_7/out')
// (2, 6, 'local_g0_7')
// (2, 6, 'lutff_7/in_2')
// (2, 6, 'neigh_op_bot_7')
// (3, 4, 'neigh_op_tnl_7')
// (3, 5, 'neigh_op_lft_7')
// (3, 6, 'local_g3_7')
// (3, 6, 'lutff_5/in_1')
// (3, 6, 'neigh_op_bnl_7')

reg n208 = 0;
// (1, 4, 'sp4_r_v_b_42')
// (1, 5, 'sp4_r_v_b_31')
// (1, 6, 'local_g3_2')
// (1, 6, 'lutff_1/in_2')
// (1, 6, 'sp4_r_v_b_18')
// (1, 7, 'sp4_r_v_b_7')
// (1, 9, 'sp4_h_r_5')
// (2, 3, 'sp4_v_t_42')
// (2, 4, 'sp4_v_b_42')
// (2, 5, 'sp4_v_b_31')
// (2, 6, 'sp4_v_b_18')
// (2, 7, 'sp4_h_r_7')
// (2, 7, 'sp4_v_b_7')
// (2, 9, 'local_g0_0')
// (2, 9, 'lutff_1/in_1')
// (2, 9, 'sp4_h_r_16')
// (3, 7, 'sp4_h_r_18')
// (3, 9, 'sp4_h_r_29')
// (4, 7, 'sp4_h_r_31')
// (4, 9, 'sp4_h_r_40')
// (5, 7, 'sp4_h_r_42')
// (5, 9, 'sp4_h_l_40')
// (5, 9, 'sp4_h_r_2')
// (6, 7, 'sp4_h_l_42')
// (6, 7, 'sp4_h_r_7')
// (6, 9, 'sp4_h_r_15')
// (7, 7, 'sp4_h_r_18')
// (7, 9, 'sp4_h_r_26')
// (8, 6, 'neigh_op_tnr_5')
// (8, 6, 'sp4_r_v_b_39')
// (8, 7, 'neigh_op_rgt_5')
// (8, 7, 'sp4_h_r_31')
// (8, 7, 'sp4_r_v_b_26')
// (8, 8, 'neigh_op_bnr_5')
// (8, 8, 'sp4_r_v_b_15')
// (8, 9, 'sp4_h_r_39')
// (8, 9, 'sp4_r_v_b_2')
// (9, 5, 'sp4_v_t_39')
// (9, 6, 'neigh_op_top_5')
// (9, 6, 'sp4_v_b_39')
// (9, 7, 'local_g3_5')
// (9, 7, 'lutff_0/in_2')
// (9, 7, 'lutff_5/out')
// (9, 7, 'sp4_h_r_42')
// (9, 7, 'sp4_v_b_26')
// (9, 8, 'neigh_op_bot_5')
// (9, 8, 'sp4_v_b_15')
// (9, 9, 'sp4_h_l_39')
// (9, 9, 'sp4_v_b_2')
// (10, 6, 'neigh_op_tnl_5')
// (10, 7, 'neigh_op_lft_5')
// (10, 7, 'sp4_h_l_42')
// (10, 8, 'neigh_op_bnl_5')

reg n209 = 0;
// (1, 4, 'sp4_r_v_b_47')
// (1, 5, 'sp4_r_v_b_34')
// (1, 6, 'local_g3_7')
// (1, 6, 'lutff_0/in_2')
// (1, 6, 'sp4_r_v_b_23')
// (1, 7, 'sp4_r_v_b_10')
// (1, 8, 'local_g1_6')
// (1, 8, 'lutff_0/in_1')
// (1, 8, 'sp4_h_r_6')
// (1, 9, 'sp4_h_r_0')
// (2, 3, 'sp4_v_t_47')
// (2, 4, 'sp4_v_b_47')
// (2, 5, 'sp4_v_b_34')
// (2, 6, 'sp4_v_b_23')
// (2, 7, 'sp4_h_r_5')
// (2, 7, 'sp4_v_b_10')
// (2, 8, 'sp4_h_r_19')
// (2, 8, 'sp4_h_r_5')
// (2, 9, 'local_g1_5')
// (2, 9, 'lutff_0/in_2')
// (2, 9, 'lutff_1/in_3')
// (2, 9, 'sp4_h_r_13')
// (3, 7, 'sp4_h_r_16')
// (3, 8, 'local_g0_0')
// (3, 8, 'lutff_4/in_0')
// (3, 8, 'sp4_h_r_16')
// (3, 8, 'sp4_h_r_30')
// (3, 9, 'sp4_h_r_24')
// (4, 7, 'sp4_h_r_29')
// (4, 8, 'sp4_h_r_29')
// (4, 8, 'sp4_h_r_43')
// (4, 9, 'sp4_h_r_37')
// (5, 7, 'sp4_h_r_40')
// (5, 8, 'sp4_h_l_43')
// (5, 8, 'sp4_h_r_40')
// (5, 8, 'sp4_h_r_6')
// (5, 9, 'sp4_h_l_37')
// (5, 9, 'sp4_h_r_9')
// (6, 7, 'sp4_h_l_40')
// (6, 7, 'sp4_h_r_9')
// (6, 8, 'sp4_h_l_40')
// (6, 8, 'sp4_h_r_19')
// (6, 8, 'sp4_h_r_5')
// (6, 9, 'sp4_h_r_20')
// (7, 7, 'sp4_h_r_20')
// (7, 8, 'sp4_h_r_16')
// (7, 8, 'sp4_h_r_30')
// (7, 9, 'sp4_h_r_33')
// (8, 5, 'sp4_r_v_b_36')
// (8, 6, 'neigh_op_tnr_6')
// (8, 6, 'sp4_r_v_b_25')
// (8, 6, 'sp4_r_v_b_41')
// (8, 7, 'neigh_op_rgt_6')
// (8, 7, 'sp4_h_r_33')
// (8, 7, 'sp4_r_v_b_12')
// (8, 7, 'sp4_r_v_b_28')
// (8, 8, 'neigh_op_bnr_6')
// (8, 8, 'sp4_h_r_29')
// (8, 8, 'sp4_h_r_43')
// (8, 8, 'sp4_r_v_b_1')
// (8, 8, 'sp4_r_v_b_17')
// (8, 9, 'sp4_h_r_44')
// (8, 9, 'sp4_r_v_b_4')
// (9, 4, 'sp4_v_t_36')
// (9, 5, 'sp4_r_v_b_37')
// (9, 5, 'sp4_v_b_36')
// (9, 5, 'sp4_v_t_41')
// (9, 6, 'neigh_op_top_6')
// (9, 6, 'sp4_r_v_b_24')
// (9, 6, 'sp4_v_b_25')
// (9, 6, 'sp4_v_b_41')
// (9, 7, 'lutff_6/out')
// (9, 7, 'sp4_h_r_44')
// (9, 7, 'sp4_r_v_b_13')
// (9, 7, 'sp4_v_b_12')
// (9, 7, 'sp4_v_b_28')
// (9, 8, 'local_g0_6')
// (9, 8, 'lutff_0/in_0')
// (9, 8, 'neigh_op_bot_6')
// (9, 8, 'sp4_h_l_43')
// (9, 8, 'sp4_h_r_40')
// (9, 8, 'sp4_r_v_b_0')
// (9, 8, 'sp4_v_b_1')
// (9, 8, 'sp4_v_b_17')
// (9, 9, 'sp4_h_l_44')
// (9, 9, 'sp4_v_b_4')
// (10, 4, 'sp4_v_t_37')
// (10, 5, 'sp4_v_b_37')
// (10, 6, 'neigh_op_tnl_6')
// (10, 6, 'sp4_v_b_24')
// (10, 7, 'neigh_op_lft_6')
// (10, 7, 'sp4_h_l_44')
// (10, 7, 'sp4_v_b_13')
// (10, 8, 'neigh_op_bnl_6')
// (10, 8, 'sp4_h_l_40')
// (10, 8, 'sp4_v_b_0')

wire n210;
// (1, 5, 'neigh_op_tnr_6')
// (1, 6, 'neigh_op_rgt_6')
// (1, 7, 'neigh_op_bnr_6')
// (2, 5, 'neigh_op_top_6')
// (2, 6, 'lutff_6/out')
// (2, 7, 'neigh_op_bot_6')
// (3, 5, 'local_g3_6')
// (3, 5, 'lutff_2/in_3')
// (3, 5, 'neigh_op_tnl_6')
// (3, 6, 'neigh_op_lft_6')
// (3, 7, 'neigh_op_bnl_6')

wire n211;
// (1, 5, 'neigh_op_tnr_7')
// (1, 6, 'neigh_op_rgt_7')
// (1, 7, 'neigh_op_bnr_7')
// (2, 5, 'local_g1_7')
// (2, 5, 'lutff_2/in_2')
// (2, 5, 'neigh_op_top_7')
// (2, 6, 'lutff_7/out')
// (2, 7, 'neigh_op_bot_7')
// (3, 5, 'neigh_op_tnl_7')
// (3, 6, 'neigh_op_lft_7')
// (3, 7, 'neigh_op_bnl_7')

reg n212 = 0;
// (1, 5, 'sp4_h_r_11')
// (1, 16, 'sp12_h_r_0')
// (2, 5, 'local_g1_6')
// (2, 5, 'lutff_2/in_3')
// (2, 5, 'sp4_h_r_22')
// (2, 9, 'sp4_r_v_b_39')
// (2, 9, 'sp4_r_v_b_41')
// (2, 10, 'sp4_r_v_b_26')
// (2, 10, 'sp4_r_v_b_28')
// (2, 11, 'sp4_r_v_b_15')
// (2, 11, 'sp4_r_v_b_17')
// (2, 12, 'local_g1_2')
// (2, 12, 'lutff_7/in_2')
// (2, 12, 'sp4_r_v_b_2')
// (2, 12, 'sp4_r_v_b_4')
// (2, 13, 'sp4_r_v_b_41')
// (2, 14, 'sp4_r_v_b_28')
// (2, 15, 'local_g3_1')
// (2, 15, 'lutff_7/in_1')
// (2, 15, 'sp4_r_v_b_17')
// (2, 16, 'sp12_h_r_3')
// (2, 16, 'sp4_r_v_b_4')
// (3, 5, 'sp4_h_r_35')
// (3, 8, 'sp4_h_r_4')
// (3, 8, 'sp4_h_r_8')
// (3, 8, 'sp4_v_t_39')
// (3, 8, 'sp4_v_t_41')
// (3, 9, 'sp4_v_b_39')
// (3, 9, 'sp4_v_b_41')
// (3, 10, 'sp4_v_b_26')
// (3, 10, 'sp4_v_b_28')
// (3, 11, 'sp4_v_b_15')
// (3, 11, 'sp4_v_b_17')
// (3, 12, 'sp4_v_b_2')
// (3, 12, 'sp4_v_b_4')
// (3, 12, 'sp4_v_t_41')
// (3, 13, 'sp4_v_b_41')
// (3, 14, 'sp4_v_b_28')
// (3, 15, 'sp4_v_b_17')
// (3, 16, 'sp12_h_r_4')
// (3, 16, 'sp4_v_b_4')
// (4, 1, 'sp4_r_v_b_39')
// (4, 2, 'local_g3_1')
// (4, 2, 'lutff_7/in_1')
// (4, 2, 'sp4_r_v_b_26')
// (4, 2, 'sp4_r_v_b_41')
// (4, 2, 'sp4_r_v_b_46')
// (4, 3, 'sp4_r_v_b_15')
// (4, 3, 'sp4_r_v_b_28')
// (4, 3, 'sp4_r_v_b_35')
// (4, 4, 'sp4_r_v_b_17')
// (4, 4, 'sp4_r_v_b_2')
// (4, 4, 'sp4_r_v_b_22')
// (4, 5, 'local_g2_3')
// (4, 5, 'lutff_4/in_3')
// (4, 5, 'sp4_h_r_46')
// (4, 5, 'sp4_r_v_b_11')
// (4, 5, 'sp4_r_v_b_4')
// (4, 5, 'sp4_r_v_b_41')
// (4, 6, 'sp4_r_v_b_28')
// (4, 7, 'sp4_r_v_b_17')
// (4, 8, 'local_g1_1')
// (4, 8, 'lutff_6/in_2')
// (4, 8, 'sp4_h_r_17')
// (4, 8, 'sp4_h_r_21')
// (4, 8, 'sp4_r_v_b_4')
// (4, 9, 'sp4_r_v_b_40')
// (4, 10, 'sp4_r_v_b_29')
// (4, 11, 'sp4_r_v_b_16')
// (4, 12, 'sp4_r_v_b_5')
// (4, 13, 'sp4_r_v_b_36')
// (4, 14, 'sp4_r_v_b_25')
// (4, 15, 'sp4_r_v_b_12')
// (4, 16, 'sp12_h_r_7')
// (4, 16, 'sp4_r_v_b_1')
// (5, 0, 'span4_vert_39')
// (5, 1, 'sp4_v_b_39')
// (5, 1, 'sp4_v_t_41')
// (5, 1, 'sp4_v_t_46')
// (5, 2, 'sp4_v_b_26')
// (5, 2, 'sp4_v_b_41')
// (5, 2, 'sp4_v_b_46')
// (5, 3, 'local_g1_7')
// (5, 3, 'lutff_2/in_2')
// (5, 3, 'sp4_v_b_15')
// (5, 3, 'sp4_v_b_28')
// (5, 3, 'sp4_v_b_35')
// (5, 4, 'sp4_h_r_2')
// (5, 4, 'sp4_v_b_17')
// (5, 4, 'sp4_v_b_2')
// (5, 4, 'sp4_v_b_22')
// (5, 4, 'sp4_v_t_41')
// (5, 5, 'sp4_h_l_46')
// (5, 5, 'sp4_h_r_11')
// (5, 5, 'sp4_v_b_11')
// (5, 5, 'sp4_v_b_4')
// (5, 5, 'sp4_v_b_41')
// (5, 6, 'sp4_v_b_28')
// (5, 7, 'local_g0_1')
// (5, 7, 'lutff_6/in_1')
// (5, 7, 'sp4_v_b_17')
// (5, 8, 'sp4_h_r_11')
// (5, 8, 'sp4_h_r_28')
// (5, 8, 'sp4_h_r_32')
// (5, 8, 'sp4_h_r_4')
// (5, 8, 'sp4_v_b_4')
// (5, 8, 'sp4_v_t_40')
// (5, 9, 'sp4_v_b_40')
// (5, 10, 'sp4_v_b_29')
// (5, 11, 'sp4_v_b_16')
// (5, 12, 'local_g1_5')
// (5, 12, 'lutff_2/in_2')
// (5, 12, 'sp4_v_b_5')
// (5, 12, 'sp4_v_t_36')
// (5, 13, 'sp4_v_b_36')
// (5, 14, 'sp4_v_b_25')
// (5, 15, 'local_g1_4')
// (5, 15, 'lutff_3/in_2')
// (5, 15, 'sp4_v_b_12')
// (5, 16, 'local_g1_0')
// (5, 16, 'lutff_4/in_3')
// (5, 16, 'sp12_h_r_8')
// (5, 16, 'sp4_v_b_1')
// (6, 4, 'sp4_h_r_15')
// (6, 5, 'sp4_h_r_22')
// (6, 8, 'sp4_h_r_17')
// (6, 8, 'sp4_h_r_22')
// (6, 8, 'sp4_h_r_41')
// (6, 8, 'sp4_h_r_45')
// (6, 9, 'sp4_r_v_b_47')
// (6, 10, 'sp4_r_v_b_34')
// (6, 11, 'sp4_r_v_b_23')
// (6, 12, 'sp4_r_v_b_10')
// (6, 16, 'sp12_h_r_11')
// (7, 4, 'sp4_h_r_26')
// (7, 5, 'sp4_h_r_35')
// (7, 8, 'sp4_h_l_41')
// (7, 8, 'sp4_h_l_45')
// (7, 8, 'sp4_h_r_28')
// (7, 8, 'sp4_h_r_35')
// (7, 8, 'sp4_h_r_4')
// (7, 8, 'sp4_h_r_8')
// (7, 8, 'sp4_v_t_47')
// (7, 9, 'sp4_v_b_47')
// (7, 10, 'sp4_v_b_34')
// (7, 11, 'local_g0_7')
// (7, 11, 'lutff_6/in_1')
// (7, 11, 'sp4_v_b_23')
// (7, 12, 'sp4_v_b_10')
// (7, 16, 'sp12_h_r_12')
// (7, 16, 'sp4_h_r_8')
// (8, 4, 'sp4_h_r_39')
// (8, 5, 'sp4_h_r_46')
// (8, 8, 'sp4_h_r_17')
// (8, 8, 'sp4_h_r_21')
// (8, 8, 'sp4_h_r_41')
// (8, 8, 'sp4_h_r_46')
// (8, 15, 'sp4_r_v_b_44')
// (8, 16, 'local_g0_5')
// (8, 16, 'lutff_1/in_0')
// (8, 16, 'sp12_h_r_15')
// (8, 16, 'sp4_h_r_21')
// (8, 16, 'sp4_r_v_b_33')
// (8, 17, 'sp4_r_v_b_20')
// (8, 18, 'local_g2_1')
// (8, 18, 'lutff_1/in_2')
// (8, 18, 'sp4_r_v_b_9')
// (9, 4, 'sp4_h_l_39')
// (9, 4, 'sp4_h_r_6')
// (9, 5, 'sp4_h_l_46')
// (9, 5, 'sp4_h_r_11')
// (9, 8, 'sp4_h_l_41')
// (9, 8, 'sp4_h_l_46')
// (9, 8, 'sp4_h_r_28')
// (9, 8, 'sp4_h_r_32')
// (9, 8, 'sp4_h_r_8')
// (9, 9, 'sp4_h_r_5')
// (9, 13, 'sp4_h_r_6')
// (9, 14, 'sp4_h_r_9')
// (9, 14, 'sp4_v_t_44')
// (9, 15, 'sp4_v_b_44')
// (9, 16, 'sp12_h_r_16')
// (9, 16, 'sp4_h_r_32')
// (9, 16, 'sp4_v_b_33')
// (9, 17, 'sp4_v_b_20')
// (9, 18, 'sp4_v_b_9')
// (10, 4, 'sp4_h_r_19')
// (10, 5, 'local_g0_6')
// (10, 5, 'lutff_1/in_3')
// (10, 5, 'sp4_h_r_22')
// (10, 5, 'sp4_r_v_b_45')
// (10, 6, 'sp4_r_v_b_32')
// (10, 7, 'sp4_r_v_b_21')
// (10, 8, 'sp4_h_r_21')
// (10, 8, 'sp4_h_r_41')
// (10, 8, 'sp4_h_r_45')
// (10, 8, 'sp4_r_v_b_8')
// (10, 9, 'sp4_h_r_16')
// (10, 9, 'sp4_r_v_b_39')
// (10, 9, 'sp4_r_v_b_45')
// (10, 10, 'sp4_r_v_b_26')
// (10, 10, 'sp4_r_v_b_32')
// (10, 11, 'local_g2_7')
// (10, 11, 'lutff_5/in_2')
// (10, 11, 'sp4_r_v_b_15')
// (10, 11, 'sp4_r_v_b_21')
// (10, 12, 'local_g2_0')
// (10, 12, 'lutff_0/in_2')
// (10, 12, 'sp4_r_v_b_2')
// (10, 12, 'sp4_r_v_b_8')
// (10, 13, 'local_g1_3')
// (10, 13, 'lutff_2/in_2')
// (10, 13, 'lutff_6/in_0')
// (10, 13, 'sp4_h_r_19')
// (10, 13, 'sp4_r_v_b_41')
// (10, 13, 'sp4_r_v_b_45')
// (10, 14, 'local_g1_4')
// (10, 14, 'lutff_0/in_3')
// (10, 14, 'sp4_h_r_20')
// (10, 14, 'sp4_r_v_b_28')
// (10, 14, 'sp4_r_v_b_32')
// (10, 15, 'local_g3_1')
// (10, 15, 'lutff_0/in_0')
// (10, 15, 'lutff_4/in_2')
// (10, 15, 'sp4_r_v_b_17')
// (10, 15, 'sp4_r_v_b_21')
// (10, 16, 'local_g2_0')
// (10, 16, 'lutff_6/in_0')
// (10, 16, 'sp12_h_r_19')
// (10, 16, 'sp4_h_r_45')
// (10, 16, 'sp4_r_v_b_4')
// (10, 16, 'sp4_r_v_b_8')
// (10, 17, 'sp4_r_v_b_46')
// (10, 18, 'sp4_r_v_b_35')
// (10, 19, 'sp4_r_v_b_22')
// (10, 20, 'sp4_r_v_b_11')
// (11, 4, 'local_g3_6')
// (11, 4, 'lutff_1/in_2')
// (11, 4, 'lutff_7/in_2')
// (11, 4, 'sp4_h_r_30')
// (11, 4, 'sp4_v_t_45')
// (11, 5, 'local_g2_3')
// (11, 5, 'lutff_5/in_0')
// (11, 5, 'lutff_7/in_2')
// (11, 5, 'sp4_h_r_35')
// (11, 5, 'sp4_v_b_45')
// (11, 6, 'local_g3_0')
// (11, 6, 'lutff_4/in_3')
// (11, 6, 'sp4_v_b_32')
// (11, 7, 'sp4_v_b_21')
// (11, 8, 'local_g1_0')
// (11, 8, 'lutff_0/in_1')
// (11, 8, 'lutff_4/in_1')
// (11, 8, 'sp4_h_l_41')
// (11, 8, 'sp4_h_l_45')
// (11, 8, 'sp4_h_r_32')
// (11, 8, 'sp4_h_r_8')
// (11, 8, 'sp4_v_b_8')
// (11, 8, 'sp4_v_t_39')
// (11, 8, 'sp4_v_t_45')
// (11, 9, 'local_g2_5')
// (11, 9, 'lutff_0/in_1')
// (11, 9, 'sp4_h_r_29')
// (11, 9, 'sp4_r_v_b_40')
// (11, 9, 'sp4_v_b_39')
// (11, 9, 'sp4_v_b_45')
// (11, 10, 'local_g3_0')
// (11, 10, 'lutff_3/in_0')
// (11, 10, 'sp4_r_v_b_29')
// (11, 10, 'sp4_v_b_26')
// (11, 10, 'sp4_v_b_32')
// (11, 11, 'sp4_r_v_b_16')
// (11, 11, 'sp4_v_b_15')
// (11, 11, 'sp4_v_b_21')
// (11, 12, 'local_g1_0')
// (11, 12, 'lutff_4/in_1')
// (11, 12, 'sp4_r_v_b_5')
// (11, 12, 'sp4_v_b_2')
// (11, 12, 'sp4_v_b_8')
// (11, 12, 'sp4_v_t_41')
// (11, 12, 'sp4_v_t_45')
// (11, 13, 'sp4_h_r_30')
// (11, 13, 'sp4_v_b_41')
// (11, 13, 'sp4_v_b_45')
// (11, 14, 'local_g3_0')
// (11, 14, 'lutff_2/in_1')
// (11, 14, 'sp4_h_r_33')
// (11, 14, 'sp4_v_b_28')
// (11, 14, 'sp4_v_b_32')
// (11, 15, 'sp4_v_b_17')
// (11, 15, 'sp4_v_b_21')
// (11, 16, 'local_g1_4')
// (11, 16, 'lutff_4/in_3')
// (11, 16, 'sp12_h_r_20')
// (11, 16, 'sp4_h_l_45')
// (11, 16, 'sp4_v_b_4')
// (11, 16, 'sp4_v_b_8')
// (11, 16, 'sp4_v_t_46')
// (11, 17, 'local_g2_6')
// (11, 17, 'lutff_6/in_0')
// (11, 17, 'lutff_7/in_3')
// (11, 17, 'sp4_v_b_46')
// (11, 18, 'sp4_v_b_35')
// (11, 19, 'sp4_v_b_22')
// (11, 20, 'sp4_v_b_11')
// (12, 4, 'local_g2_3')
// (12, 4, 'lutff_6/in_3')
// (12, 4, 'sp4_h_r_43')
// (12, 5, 'sp4_h_r_46')
// (12, 5, 'sp4_r_v_b_37')
// (12, 6, 'sp4_r_v_b_24')
// (12, 6, 'sp4_r_v_b_40')
// (12, 7, 'neigh_op_tnr_0')
// (12, 7, 'sp4_r_v_b_13')
// (12, 7, 'sp4_r_v_b_29')
// (12, 7, 'sp4_r_v_b_45')
// (12, 8, 'neigh_op_rgt_0')
// (12, 8, 'sp4_h_r_21')
// (12, 8, 'sp4_h_r_45')
// (12, 8, 'sp4_h_r_5')
// (12, 8, 'sp4_r_v_b_0')
// (12, 8, 'sp4_r_v_b_16')
// (12, 8, 'sp4_r_v_b_32')
// (12, 8, 'sp4_v_t_40')
// (12, 9, 'local_g0_0')
// (12, 9, 'lutff_6/in_2')
// (12, 9, 'neigh_op_bnr_0')
// (12, 9, 'sp4_h_r_40')
// (12, 9, 'sp4_r_v_b_21')
// (12, 9, 'sp4_r_v_b_5')
// (12, 9, 'sp4_v_b_40')
// (12, 10, 'local_g2_0')
// (12, 10, 'lutff_1/in_3')
// (12, 10, 'sp4_r_v_b_36')
// (12, 10, 'sp4_r_v_b_8')
// (12, 10, 'sp4_v_b_29')
// (12, 11, 'sp4_r_v_b_25')
// (12, 11, 'sp4_r_v_b_41')
// (12, 11, 'sp4_v_b_16')
// (12, 12, 'local_g1_5')
// (12, 12, 'lutff_0/in_2')
// (12, 12, 'sp4_r_v_b_12')
// (12, 12, 'sp4_r_v_b_28')
// (12, 12, 'sp4_v_b_5')
// (12, 13, 'local_g3_1')
// (12, 13, 'lutff_2/in_2')
// (12, 13, 'sp4_h_r_43')
// (12, 13, 'sp4_r_v_b_1')
// (12, 13, 'sp4_r_v_b_17')
// (12, 14, 'sp4_h_r_44')
// (12, 14, 'sp4_r_v_b_4')
// (12, 16, 'sp12_h_r_23')
// (13, 1, 'sp4_r_v_b_36')
// (13, 2, 'sp4_r_v_b_25')
// (13, 3, 'sp4_r_v_b_12')
// (13, 4, 'sp12_v_t_23')
// (13, 4, 'sp4_h_l_43')
// (13, 4, 'sp4_r_v_b_1')
// (13, 4, 'sp4_v_t_37')
// (13, 5, 'sp12_v_b_23')
// (13, 5, 'sp4_h_l_46')
// (13, 5, 'sp4_r_v_b_36')
// (13, 5, 'sp4_v_b_37')
// (13, 5, 'sp4_v_t_40')
// (13, 6, 'sp12_v_b_20')
// (13, 6, 'sp4_r_v_b_25')
// (13, 6, 'sp4_v_b_24')
// (13, 6, 'sp4_v_b_40')
// (13, 6, 'sp4_v_t_45')
// (13, 7, 'neigh_op_top_0')
// (13, 7, 'sp12_v_b_19')
// (13, 7, 'sp4_r_v_b_12')
// (13, 7, 'sp4_v_b_13')
// (13, 7, 'sp4_v_b_29')
// (13, 7, 'sp4_v_b_45')
// (13, 8, 'lutff_0/out')
// (13, 8, 'sp12_v_b_16')
// (13, 8, 'sp4_h_l_45')
// (13, 8, 'sp4_h_r_0')
// (13, 8, 'sp4_h_r_16')
// (13, 8, 'sp4_h_r_32')
// (13, 8, 'sp4_r_v_b_1')
// (13, 8, 'sp4_v_b_0')
// (13, 8, 'sp4_v_b_16')
// (13, 8, 'sp4_v_b_32')
// (13, 9, 'local_g0_0')
// (13, 9, 'lutff_0/in_0')
// (13, 9, 'neigh_op_bot_0')
// (13, 9, 'sp12_v_b_15')
// (13, 9, 'sp4_h_l_40')
// (13, 9, 'sp4_v_b_21')
// (13, 9, 'sp4_v_b_5')
// (13, 9, 'sp4_v_t_36')
// (13, 10, 'sp12_v_b_12')
// (13, 10, 'sp4_v_b_36')
// (13, 10, 'sp4_v_b_8')
// (13, 10, 'sp4_v_t_41')
// (13, 11, 'sp12_v_b_11')
// (13, 11, 'sp4_v_b_25')
// (13, 11, 'sp4_v_b_41')
// (13, 12, 'sp12_v_b_8')
// (13, 12, 'sp4_v_b_12')
// (13, 12, 'sp4_v_b_28')
// (13, 13, 'sp12_v_b_7')
// (13, 13, 'sp4_h_l_43')
// (13, 13, 'sp4_v_b_1')
// (13, 13, 'sp4_v_b_17')
// (13, 14, 'sp12_v_b_4')
// (13, 14, 'sp4_h_l_44')
// (13, 14, 'sp4_v_b_4')
// (13, 15, 'sp12_v_b_3')
// (13, 16, 'local_g3_0')
// (13, 16, 'lutff_6/in_3')
// (13, 16, 'lutff_7/in_2')
// (13, 16, 'sp12_h_l_23')
// (13, 16, 'sp12_v_b_0')
// (14, 0, 'span4_vert_36')
// (14, 1, 'sp4_v_b_36')
// (14, 2, 'local_g2_1')
// (14, 2, 'lutff_5/in_0')
// (14, 2, 'sp4_v_b_25')
// (14, 3, 'sp4_v_b_12')
// (14, 4, 'sp4_v_b_1')
// (14, 4, 'sp4_v_t_36')
// (14, 5, 'sp4_v_b_36')
// (14, 6, 'sp4_v_b_25')
// (14, 7, 'neigh_op_tnl_0')
// (14, 7, 'sp4_v_b_12')
// (14, 8, 'neigh_op_lft_0')
// (14, 8, 'sp4_h_r_13')
// (14, 8, 'sp4_h_r_29')
// (14, 8, 'sp4_h_r_45')
// (14, 8, 'sp4_v_b_1')
// (14, 9, 'neigh_op_bnl_0')
// (15, 8, 'sp4_h_l_45')
// (15, 8, 'sp4_h_r_24')
// (15, 8, 'sp4_h_r_4')
// (15, 8, 'sp4_h_r_40')
// (15, 9, 'sp4_r_v_b_40')
// (15, 9, 'sp4_r_v_b_47')
// (15, 10, 'sp4_r_v_b_29')
// (15, 10, 'sp4_r_v_b_34')
// (15, 11, 'sp4_r_v_b_16')
// (15, 11, 'sp4_r_v_b_23')
// (15, 12, 'sp4_r_v_b_10')
// (15, 12, 'sp4_r_v_b_5')
// (15, 13, 'sp4_r_v_b_40')
// (15, 13, 'sp4_r_v_b_43')
// (15, 14, 'sp4_r_v_b_29')
// (15, 14, 'sp4_r_v_b_30')
// (15, 15, 'local_g3_0')
// (15, 15, 'local_g3_3')
// (15, 15, 'lutff_0/in_1')
// (15, 15, 'lutff_4/in_2')
// (15, 15, 'lutff_5/in_1')
// (15, 15, 'sp4_r_v_b_16')
// (15, 15, 'sp4_r_v_b_19')
// (15, 16, 'sp4_r_v_b_5')
// (15, 16, 'sp4_r_v_b_6')
// (16, 8, 'sp4_h_l_40')
// (16, 8, 'sp4_h_r_17')
// (16, 8, 'sp4_h_r_37')
// (16, 8, 'sp4_v_t_40')
// (16, 8, 'sp4_v_t_47')
// (16, 9, 'sp4_v_b_40')
// (16, 9, 'sp4_v_b_47')
// (16, 10, 'sp4_v_b_29')
// (16, 10, 'sp4_v_b_34')
// (16, 11, 'sp4_v_b_16')
// (16, 11, 'sp4_v_b_23')
// (16, 12, 'sp4_v_b_10')
// (16, 12, 'sp4_v_b_5')
// (16, 12, 'sp4_v_t_40')
// (16, 12, 'sp4_v_t_43')
// (16, 13, 'sp4_v_b_40')
// (16, 13, 'sp4_v_b_43')
// (16, 14, 'local_g3_5')
// (16, 14, 'local_g3_6')
// (16, 14, 'lutff_4/in_3')
// (16, 14, 'lutff_6/in_2')
// (16, 14, 'lutff_7/in_3')
// (16, 14, 'sp4_v_b_29')
// (16, 14, 'sp4_v_b_30')
// (16, 15, 'sp4_v_b_16')
// (16, 15, 'sp4_v_b_19')
// (16, 16, 'sp4_v_b_5')
// (16, 16, 'sp4_v_b_6')
// (17, 8, 'sp4_h_l_37')
// (17, 8, 'sp4_h_r_28')
// (18, 8, 'sp4_h_r_41')
// (18, 9, 'sp4_r_v_b_44')
// (18, 10, 'local_g2_1')
// (18, 10, 'lutff_6/in_3')
// (18, 10, 'sp4_r_v_b_33')
// (18, 11, 'sp4_r_v_b_20')
// (18, 12, 'sp4_r_v_b_9')
// (19, 8, 'sp4_h_l_41')
// (19, 8, 'sp4_v_t_44')
// (19, 9, 'sp4_v_b_44')
// (19, 10, 'sp4_v_b_33')
// (19, 11, 'sp4_v_b_20')
// (19, 12, 'sp4_v_b_9')

reg n213 = 0;
// (1, 5, 'sp4_h_r_6')
// (2, 4, 'neigh_op_tnr_7')
// (2, 5, 'neigh_op_rgt_7')
// (2, 5, 'sp4_h_r_19')
// (2, 6, 'neigh_op_bnr_7')
// (3, 3, 'sp4_r_v_b_39')
// (3, 4, 'neigh_op_top_7')
// (3, 4, 'sp4_r_v_b_26')
// (3, 4, 'sp4_r_v_b_42')
// (3, 5, 'lutff_7/out')
// (3, 5, 'sp4_h_r_30')
// (3, 5, 'sp4_r_v_b_15')
// (3, 5, 'sp4_r_v_b_31')
// (3, 6, 'neigh_op_bot_7')
// (3, 6, 'sp4_r_v_b_18')
// (3, 6, 'sp4_r_v_b_2')
// (3, 7, 'sp4_r_v_b_7')
// (4, 2, 'sp4_r_v_b_37')
// (4, 2, 'sp4_v_t_39')
// (4, 3, 'sp4_r_v_b_24')
// (4, 3, 'sp4_v_b_39')
// (4, 3, 'sp4_v_t_42')
// (4, 4, 'neigh_op_tnl_7')
// (4, 4, 'sp4_r_v_b_13')
// (4, 4, 'sp4_v_b_26')
// (4, 4, 'sp4_v_b_42')
// (4, 5, 'neigh_op_lft_7')
// (4, 5, 'sp4_h_r_43')
// (4, 5, 'sp4_r_v_b_0')
// (4, 5, 'sp4_v_b_15')
// (4, 5, 'sp4_v_b_31')
// (4, 6, 'local_g3_7')
// (4, 6, 'lutff_3/in_1')
// (4, 6, 'neigh_op_bnl_7')
// (4, 6, 'sp4_h_r_2')
// (4, 6, 'sp4_r_v_b_43')
// (4, 6, 'sp4_v_b_18')
// (4, 6, 'sp4_v_b_2')
// (4, 7, 'local_g1_7')
// (4, 7, 'lutff_5/in_3')
// (4, 7, 'sp4_r_v_b_30')
// (4, 7, 'sp4_v_b_7')
// (4, 8, 'sp4_r_v_b_19')
// (4, 9, 'sp4_r_v_b_6')
// (5, 1, 'sp4_v_t_37')
// (5, 2, 'sp4_v_b_37')
// (5, 3, 'sp4_v_b_24')
// (5, 4, 'local_g1_5')
// (5, 4, 'lutff_1/in_1')
// (5, 4, 'sp4_v_b_13')
// (5, 5, 'sp4_h_l_43')
// (5, 5, 'sp4_v_b_0')
// (5, 5, 'sp4_v_t_43')
// (5, 6, 'local_g1_7')
// (5, 6, 'lutff_0/in_2')
// (5, 6, 'lutff_1/in_3')
// (5, 6, 'sp4_h_r_15')
// (5, 6, 'sp4_v_b_43')
// (5, 7, 'sp4_v_b_30')
// (5, 8, 'local_g1_3')
// (5, 8, 'lutff_4/in_2')
// (5, 8, 'sp4_v_b_19')
// (5, 9, 'sp4_v_b_6')
// (6, 6, 'sp4_h_r_26')
// (7, 6, 'sp4_h_r_39')
// (8, 6, 'sp4_h_l_39')

wire n214;
// (1, 5, 'sp4_r_v_b_47')
// (1, 6, 'local_g0_1')
// (1, 6, 'lutff_0/in_1')
// (1, 6, 'sp4_r_v_b_34')
// (1, 7, 'local_g2_5')
// (1, 7, 'lutff_0/in_1')
// (1, 7, 'neigh_op_tnr_5')
// (1, 7, 'sp4_r_v_b_23')
// (1, 8, 'local_g2_5')
// (1, 8, 'lutff_6/in_3')
// (1, 8, 'neigh_op_rgt_5')
// (1, 8, 'sp4_r_v_b_10')
// (1, 9, 'neigh_op_bnr_5')
// (2, 4, 'sp4_v_t_47')
// (2, 5, 'sp4_v_b_47')
// (2, 6, 'sp4_v_b_34')
// (2, 7, 'neigh_op_top_5')
// (2, 7, 'sp4_v_b_23')
// (2, 8, 'lutff_5/out')
// (2, 8, 'sp4_v_b_10')
// (2, 9, 'neigh_op_bot_5')
// (3, 7, 'neigh_op_tnl_5')
// (3, 8, 'neigh_op_lft_5')
// (3, 9, 'neigh_op_bnl_5')

wire n215;
// (1, 6, 'local_g2_4')
// (1, 6, 'lutff_4/in_2')
// (1, 6, 'neigh_op_tnr_4')
// (1, 7, 'neigh_op_rgt_4')
// (1, 8, 'neigh_op_bnr_4')
// (2, 6, 'neigh_op_top_4')
// (2, 7, 'lutff_4/out')
// (2, 8, 'neigh_op_bot_4')
// (3, 6, 'neigh_op_tnl_4')
// (3, 7, 'neigh_op_lft_4')
// (3, 8, 'neigh_op_bnl_4')

wire n216;
// (1, 6, 'lutff_4/cout')
// (1, 6, 'lutff_5/in_3')

wire n217;
// (1, 6, 'neigh_op_tnr_0')
// (1, 7, 'neigh_op_rgt_0')
// (1, 8, 'neigh_op_bnr_0')
// (2, 0, 'span12_vert_12')
// (2, 1, 'sp12_v_b_12')
// (2, 2, 'sp12_v_b_11')
// (2, 3, 'sp12_v_b_8')
// (2, 4, 'sp12_v_b_7')
// (2, 5, 'sp12_v_b_4')
// (2, 6, 'local_g3_3')
// (2, 6, 'lutff_global/cen')
// (2, 6, 'neigh_op_top_0')
// (2, 6, 'sp12_v_b_3')
// (2, 7, 'lutff_0/out')
// (2, 7, 'sp12_v_b_0')
// (2, 7, 'sp4_h_r_0')
// (2, 8, 'neigh_op_bot_0')
// (3, 6, 'neigh_op_tnl_0')
// (3, 7, 'neigh_op_lft_0')
// (3, 7, 'sp4_h_r_13')
// (3, 8, 'neigh_op_bnl_0')
// (4, 7, 'sp4_h_r_24')
// (5, 4, 'local_g3_3')
// (5, 4, 'lutff_global/cen')
// (5, 4, 'sp4_r_v_b_43')
// (5, 5, 'sp4_r_v_b_30')
// (5, 6, 'sp4_r_v_b_19')
// (5, 7, 'sp4_h_r_37')
// (5, 7, 'sp4_r_v_b_6')
// (6, 3, 'sp4_v_t_43')
// (6, 4, 'sp4_v_b_43')
// (6, 5, 'sp4_v_b_30')
// (6, 6, 'sp4_v_b_19')
// (6, 7, 'sp4_h_l_37')
// (6, 7, 'sp4_v_b_6')

wire n218;
// (1, 6, 'neigh_op_tnr_1')
// (1, 7, 'neigh_op_rgt_1')
// (1, 8, 'neigh_op_bnr_1')
// (2, 6, 'neigh_op_top_1')
// (2, 7, 'local_g2_1')
// (2, 7, 'lutff_1/out')
// (2, 7, 'lutff_2/in_3')
// (2, 8, 'neigh_op_bot_1')
// (3, 6, 'neigh_op_tnl_1')
// (3, 7, 'neigh_op_lft_1')
// (3, 8, 'neigh_op_bnl_1')

wire n219;
// (1, 6, 'neigh_op_tnr_2')
// (1, 7, 'neigh_op_rgt_2')
// (1, 8, 'neigh_op_bnr_2')
// (2, 6, 'neigh_op_top_2')
// (2, 7, 'local_g3_2')
// (2, 7, 'lutff_2/out')
// (2, 7, 'lutff_6/in_3')
// (2, 8, 'neigh_op_bot_2')
// (3, 6, 'neigh_op_tnl_2')
// (3, 7, 'neigh_op_lft_2')
// (3, 8, 'neigh_op_bnl_2')

wire n220;
// (1, 6, 'neigh_op_tnr_3')
// (1, 7, 'neigh_op_rgt_3')
// (1, 8, 'neigh_op_bnr_3')
// (2, 6, 'neigh_op_top_3')
// (2, 7, 'local_g1_3')
// (2, 7, 'lutff_2/in_2')
// (2, 7, 'lutff_3/out')
// (2, 8, 'neigh_op_bot_3')
// (3, 6, 'neigh_op_tnl_3')
// (3, 7, 'neigh_op_lft_3')
// (3, 8, 'neigh_op_bnl_3')

reg n221 = 0;
// (1, 6, 'neigh_op_tnr_5')
// (1, 7, 'neigh_op_rgt_5')
// (1, 8, 'neigh_op_bnr_5')
// (2, 6, 'neigh_op_top_5')
// (2, 6, 'sp4_r_v_b_38')
// (2, 7, 'lutff_5/out')
// (2, 7, 'sp4_r_v_b_27')
// (2, 8, 'neigh_op_bot_5')
// (2, 8, 'sp4_r_v_b_14')
// (2, 9, 'sp4_r_v_b_3')
// (3, 5, 'sp4_h_r_3')
// (3, 5, 'sp4_v_t_38')
// (3, 6, 'neigh_op_tnl_5')
// (3, 6, 'sp4_v_b_38')
// (3, 7, 'neigh_op_lft_5')
// (3, 7, 'sp4_v_b_27')
// (3, 8, 'neigh_op_bnl_5')
// (3, 8, 'sp4_v_b_14')
// (3, 9, 'sp4_h_r_9')
// (3, 9, 'sp4_v_b_3')
// (4, 5, 'sp4_h_r_14')
// (4, 9, 'local_g1_4')
// (4, 9, 'lutff_6/in_3')
// (4, 9, 'sp4_h_r_20')
// (5, 5, 'local_g2_3')
// (5, 5, 'lutff_5/in_0')
// (5, 5, 'sp4_h_r_27')
// (5, 9, 'sp4_h_r_33')
// (6, 5, 'sp4_h_r_38')
// (6, 9, 'sp4_h_r_44')
// (7, 5, 'sp4_h_l_38')
// (7, 9, 'sp4_h_l_44')

wire n222;
// (1, 6, 'neigh_op_tnr_6')
// (1, 7, 'neigh_op_rgt_6')
// (1, 8, 'neigh_op_bnr_6')
// (2, 5, 'sp4_r_v_b_37')
// (2, 6, 'local_g0_6')
// (2, 6, 'local_g1_6')
// (2, 6, 'lutff_2/in_0')
// (2, 6, 'lutff_3/in_0')
// (2, 6, 'lutff_4/in_0')
// (2, 6, 'lutff_5/in_0')
// (2, 6, 'neigh_op_top_6')
// (2, 6, 'sp4_r_v_b_24')
// (2, 7, 'local_g0_6')
// (2, 7, 'lutff_0/in_0')
// (2, 7, 'lutff_6/out')
// (2, 7, 'sp4_r_v_b_13')
// (2, 8, 'neigh_op_bot_6')
// (2, 8, 'sp4_r_v_b_0')
// (3, 4, 'sp4_h_r_5')
// (3, 4, 'sp4_v_t_37')
// (3, 5, 'sp4_v_b_37')
// (3, 6, 'neigh_op_tnl_6')
// (3, 6, 'sp4_v_b_24')
// (3, 7, 'neigh_op_lft_6')
// (3, 7, 'sp4_v_b_13')
// (3, 8, 'neigh_op_bnl_6')
// (3, 8, 'sp4_v_b_0')
// (4, 4, 'sp4_h_r_16')
// (5, 4, 'local_g2_5')
// (5, 4, 'lutff_3/in_0')
// (5, 4, 'lutff_5/in_2')
// (5, 4, 'sp4_h_r_29')
// (6, 4, 'sp4_h_r_40')
// (7, 4, 'sp4_h_l_40')

wire n223;
// (1, 6, 'neigh_op_tnr_7')
// (1, 7, 'neigh_op_rgt_7')
// (1, 8, 'neigh_op_bnr_7')
// (2, 1, 'sp4_r_v_b_39')
// (2, 2, 'sp4_r_v_b_26')
// (2, 3, 'sp4_r_v_b_15')
// (2, 4, 'sp4_r_v_b_2')
// (2, 5, 'sp4_r_v_b_39')
// (2, 6, 'neigh_op_top_7')
// (2, 6, 'sp4_r_v_b_26')
// (2, 7, 'lutff_7/out')
// (2, 7, 'sp4_r_v_b_15')
// (2, 8, 'neigh_op_bot_7')
// (2, 8, 'sp4_r_v_b_2')
// (3, 0, 'span4_vert_39')
// (3, 1, 'sp4_v_b_39')
// (3, 2, 'sp4_v_b_26')
// (3, 3, 'local_g0_7')
// (3, 3, 'lutff_5/in_2')
// (3, 3, 'sp4_v_b_15')
// (3, 4, 'sp4_v_b_2')
// (3, 4, 'sp4_v_t_39')
// (3, 5, 'sp4_v_b_39')
// (3, 6, 'neigh_op_tnl_7')
// (3, 6, 'sp4_v_b_26')
// (3, 7, 'neigh_op_lft_7')
// (3, 7, 'sp4_v_b_15')
// (3, 8, 'neigh_op_bnl_7')
// (3, 8, 'sp4_v_b_2')

wire n224;
// (1, 6, 'sp4_h_r_2')
// (1, 7, 'sp4_r_v_b_43')
// (1, 8, 'sp4_r_v_b_30')
// (1, 9, 'sp4_r_v_b_19')
// (1, 10, 'sp4_r_v_b_6')
// (2, 6, 'sp4_h_r_15')
// (2, 6, 'sp4_h_r_6')
// (2, 6, 'sp4_v_t_43')
// (2, 7, 'local_g3_3')
// (2, 7, 'lutff_global/cen')
// (2, 7, 'sp4_v_b_43')
// (2, 8, 'sp4_v_b_30')
// (2, 9, 'sp4_v_b_19')
// (2, 10, 'sp4_v_b_6')
// (3, 4, 'sp4_r_v_b_38')
// (3, 5, 'sp4_r_v_b_27')
// (3, 6, 'local_g2_2')
// (3, 6, 'lutff_global/cen')
// (3, 6, 'sp4_h_r_19')
// (3, 6, 'sp4_h_r_26')
// (3, 6, 'sp4_r_v_b_14')
// (3, 7, 'local_g1_3')
// (3, 7, 'lutff_global/cen')
// (3, 7, 'sp4_r_v_b_3')
// (4, 3, 'sp4_v_t_38')
// (4, 4, 'sp4_v_b_38')
// (4, 5, 'sp4_v_b_27')
// (4, 6, 'sp4_h_r_30')
// (4, 6, 'sp4_h_r_39')
// (4, 6, 'sp4_v_b_14')
// (4, 7, 'sp4_h_r_3')
// (4, 7, 'sp4_v_b_3')
// (5, 6, 'sp4_h_l_39')
// (5, 6, 'sp4_h_r_11')
// (5, 6, 'sp4_h_r_43')
// (5, 7, 'sp4_h_r_14')
// (6, 3, 'sp4_r_v_b_38')
// (6, 4, 'sp4_r_v_b_27')
// (6, 5, 'sp4_r_v_b_14')
// (6, 6, 'sp4_h_l_43')
// (6, 6, 'sp4_h_r_22')
// (6, 6, 'sp4_h_r_6')
// (6, 6, 'sp4_r_v_b_3')
// (6, 7, 'sp4_h_r_27')
// (7, 2, 'sp4_v_t_38')
// (7, 3, 'sp4_v_b_38')
// (7, 4, 'local_g3_3')
// (7, 4, 'lutff_global/cen')
// (7, 4, 'sp4_r_v_b_38')
// (7, 4, 'sp4_v_b_27')
// (7, 5, 'neigh_op_tnr_7')
// (7, 5, 'sp4_r_v_b_27')
// (7, 5, 'sp4_v_b_14')
// (7, 6, 'neigh_op_rgt_7')
// (7, 6, 'sp4_h_r_19')
// (7, 6, 'sp4_h_r_3')
// (7, 6, 'sp4_h_r_35')
// (7, 6, 'sp4_r_v_b_14')
// (7, 6, 'sp4_v_b_3')
// (7, 7, 'neigh_op_bnr_7')
// (7, 7, 'sp4_h_r_38')
// (7, 7, 'sp4_r_v_b_3')
// (8, 3, 'sp4_v_t_38')
// (8, 4, 'sp4_v_b_38')
// (8, 5, 'neigh_op_top_7')
// (8, 5, 'sp4_v_b_27')
// (8, 6, 'lutff_7/out')
// (8, 6, 'sp4_h_r_14')
// (8, 6, 'sp4_h_r_30')
// (8, 6, 'sp4_h_r_46')
// (8, 6, 'sp4_v_b_14')
// (8, 7, 'neigh_op_bot_7')
// (8, 7, 'sp4_h_l_38')
// (8, 7, 'sp4_v_b_3')
// (9, 5, 'neigh_op_tnl_7')
// (9, 6, 'neigh_op_lft_7')
// (9, 6, 'sp4_h_l_46')
// (9, 6, 'sp4_h_r_27')
// (9, 6, 'sp4_h_r_43')
// (9, 7, 'neigh_op_bnl_7')
// (10, 6, 'sp4_h_l_43')
// (10, 6, 'sp4_h_r_38')
// (11, 6, 'sp4_h_l_38')

wire n225;
// (1, 6, 'sp4_r_v_b_38')
// (1, 7, 'sp4_r_v_b_27')
// (1, 8, 'sp4_r_v_b_14')
// (1, 9, 'sp4_r_v_b_3')
// (1, 10, 'sp4_r_v_b_37')
// (1, 11, 'sp4_r_v_b_24')
// (1, 12, 'neigh_op_tnr_0')
// (1, 12, 'sp4_r_v_b_13')
// (1, 13, 'neigh_op_rgt_0')
// (1, 13, 'sp4_r_v_b_0')
// (1, 14, 'local_g1_0')
// (1, 14, 'lutff_4/in_3')
// (1, 14, 'neigh_op_bnr_0')
// (2, 5, 'sp4_v_t_38')
// (2, 6, 'sp4_v_b_38')
// (2, 7, 'local_g2_3')
// (2, 7, 'lutff_0/in_1')
// (2, 7, 'sp4_v_b_27')
// (2, 8, 'sp4_v_b_14')
// (2, 9, 'sp4_v_b_3')
// (2, 9, 'sp4_v_t_37')
// (2, 10, 'sp4_v_b_37')
// (2, 11, 'sp4_v_b_24')
// (2, 12, 'local_g1_0')
// (2, 12, 'lutff_2/in_3')
// (2, 12, 'neigh_op_top_0')
// (2, 12, 'sp4_v_b_13')
// (2, 13, 'lutff_0/out')
// (2, 13, 'sp4_v_b_0')
// (2, 14, 'neigh_op_bot_0')
// (3, 12, 'neigh_op_tnl_0')
// (3, 13, 'neigh_op_lft_0')
// (3, 14, 'neigh_op_bnl_0')

reg n226 = 0;
// (1, 7, 'local_g2_2')
// (1, 7, 'lutff_4/in_0')
// (1, 7, 'neigh_op_tnr_2')
// (1, 8, 'neigh_op_rgt_2')
// (1, 9, 'neigh_op_bnr_2')
// (2, 7, 'neigh_op_top_2')
// (2, 8, 'local_g0_2')
// (2, 8, 'lutff_2/in_2')
// (2, 8, 'lutff_2/out')
// (2, 9, 'local_g0_2')
// (2, 9, 'lutff_6/in_2')
// (2, 9, 'neigh_op_bot_2')
// (3, 7, 'neigh_op_tnl_2')
// (3, 8, 'local_g1_2')
// (3, 8, 'lutff_2/in_1')
// (3, 8, 'neigh_op_lft_2')
// (3, 9, 'local_g2_2')
// (3, 9, 'lutff_5/in_3')
// (3, 9, 'neigh_op_bnl_2')

reg n227 = 0;
// (1, 7, 'local_g3_3')
// (1, 7, 'lutff_6/in_2')
// (1, 7, 'neigh_op_tnr_3')
// (1, 8, 'neigh_op_rgt_3')
// (1, 9, 'neigh_op_bnr_3')
// (2, 7, 'neigh_op_top_3')
// (2, 8, 'local_g1_3')
// (2, 8, 'lutff_3/in_1')
// (2, 8, 'lutff_3/out')
// (2, 9, 'neigh_op_bot_3')
// (3, 7, 'neigh_op_tnl_3')
// (3, 8, 'local_g1_3')
// (3, 8, 'lutff_3/in_1')
// (3, 8, 'lutff_6/in_0')
// (3, 8, 'neigh_op_lft_3')
// (3, 9, 'neigh_op_bnl_3')

wire n228;
// (1, 7, 'lutff_0/cout')
// (1, 7, 'lutff_1/in_3')

wire n229;
// (1, 7, 'lutff_1/cout')
// (1, 7, 'lutff_2/in_3')

reg n230 = 0;
// (1, 7, 'neigh_op_tnr_4')
// (1, 8, 'neigh_op_rgt_4')
// (1, 9, 'neigh_op_bnr_4')
// (2, 7, 'local_g1_4')
// (2, 7, 'lutff_4/in_1')
// (2, 7, 'neigh_op_top_4')
// (2, 8, 'local_g2_4')
// (2, 8, 'lutff_4/in_0')
// (2, 8, 'lutff_4/out')
// (2, 9, 'neigh_op_bot_4')
// (3, 7, 'neigh_op_tnl_4')
// (3, 8, 'local_g0_4')
// (3, 8, 'lutff_6/in_2')
// (3, 8, 'neigh_op_lft_4')
// (3, 9, 'neigh_op_bnl_4')

wire n231;
// (1, 7, 'neigh_op_tnr_7')
// (1, 8, 'local_g3_7')
// (1, 8, 'lutff_1/in_1')
// (1, 8, 'neigh_op_rgt_7')
// (1, 9, 'neigh_op_bnr_7')
// (2, 7, 'neigh_op_top_7')
// (2, 8, 'lutff_7/out')
// (2, 9, 'neigh_op_bot_7')
// (3, 7, 'neigh_op_tnl_7')
// (3, 8, 'neigh_op_lft_7')
// (3, 9, 'neigh_op_bnl_7')

wire n232;
// (1, 7, 'sp4_h_r_5')
// (2, 7, 'local_g0_0')
// (2, 7, 'lutff_3/in_1')
// (2, 7, 'sp4_h_r_16')
// (3, 1, 'local_g0_0')
// (3, 1, 'lutff_3/in_1')
// (3, 1, 'sp4_r_v_b_35')
// (3, 2, 'sp4_r_v_b_22')
// (3, 3, 'sp4_r_v_b_11')
// (3, 4, 'sp4_r_v_b_45')
// (3, 5, 'sp4_r_v_b_32')
// (3, 6, 'local_g2_4')
// (3, 6, 'lutff_2/in_2')
// (3, 6, 'neigh_op_tnr_4')
// (3, 6, 'sp4_r_v_b_21')
// (3, 7, 'neigh_op_rgt_4')
// (3, 7, 'sp4_h_r_29')
// (3, 7, 'sp4_r_v_b_8')
// (3, 8, 'neigh_op_bnr_4')
// (4, 0, 'span4_vert_35')
// (4, 1, 'sp4_v_b_35')
// (4, 2, 'sp4_v_b_22')
// (4, 3, 'sp4_v_b_11')
// (4, 3, 'sp4_v_t_45')
// (4, 4, 'local_g2_5')
// (4, 4, 'lutff_0/in_1')
// (4, 4, 'lutff_7/in_2')
// (4, 4, 'sp4_v_b_45')
// (4, 5, 'sp4_v_b_32')
// (4, 6, 'local_g1_4')
// (4, 6, 'lutff_5/in_0')
// (4, 6, 'neigh_op_top_4')
// (4, 6, 'sp4_v_b_21')
// (4, 7, 'lutff_4/out')
// (4, 7, 'sp4_h_r_40')
// (4, 7, 'sp4_v_b_8')
// (4, 8, 'neigh_op_bot_4')
// (5, 6, 'neigh_op_tnl_4')
// (5, 7, 'neigh_op_lft_4')
// (5, 7, 'sp4_h_l_40')
// (5, 8, 'neigh_op_bnl_4')

reg n233 = 0;
// (1, 7, 'sp4_h_r_6')
// (2, 0, 'span12_vert_4')
// (2, 1, 'local_g3_4')
// (2, 1, 'lutff_5/in_0')
// (2, 1, 'sp12_v_b_4')
// (2, 1, 'sp4_r_v_b_26')
// (2, 2, 'sp12_v_b_3')
// (2, 2, 'sp4_r_v_b_15')
// (2, 3, 'sp12_h_r_0')
// (2, 3, 'sp12_v_b_0')
// (2, 3, 'sp4_r_v_b_2')
// (2, 7, 'local_g0_3')
// (2, 7, 'lutff_5/in_0')
// (2, 7, 'sp4_h_r_19')
// (2, 18, 'sp4_r_v_b_36')
// (2, 19, 'sp4_r_v_b_25')
// (2, 20, 'sp4_r_v_b_12')
// (2, 21, 'sp4_r_v_b_1')
// (3, 0, 'span4_vert_26')
// (3, 1, 'sp4_v_b_26')
// (3, 2, 'local_g0_7')
// (3, 2, 'lutff_1/in_2')
// (3, 2, 'sp4_v_b_15')
// (3, 3, 'local_g0_3')
// (3, 3, 'lutff_4/in_3')
// (3, 3, 'sp12_h_r_3')
// (3, 3, 'sp4_h_r_9')
// (3, 3, 'sp4_v_b_2')
// (3, 7, 'sp4_h_r_30')
// (3, 7, 'sp4_r_v_b_41')
// (3, 8, 'sp4_r_v_b_28')
// (3, 9, 'sp4_r_v_b_17')
// (3, 10, 'local_g1_4')
// (3, 10, 'lutff_7/in_0')
// (3, 10, 'sp4_r_v_b_4')
// (3, 17, 'sp4_h_r_7')
// (3, 17, 'sp4_v_t_36')
// (3, 18, 'sp4_v_b_36')
// (3, 19, 'sp4_v_b_25')
// (3, 20, 'local_g0_4')
// (3, 20, 'lutff_0/in_0')
// (3, 20, 'sp4_v_b_12')
// (3, 21, 'sp4_v_b_1')
// (4, 1, 'local_g1_0')
// (4, 1, 'lutff_4/in_3')
// (4, 1, 'sp4_r_v_b_24')
// (4, 1, 'sp4_r_v_b_27')
// (4, 2, 'local_g2_6')
// (4, 2, 'lutff_0/in_2')
// (4, 2, 'sp4_r_v_b_13')
// (4, 2, 'sp4_r_v_b_14')
// (4, 3, 'sp12_h_r_4')
// (4, 3, 'sp4_h_r_20')
// (4, 3, 'sp4_r_v_b_0')
// (4, 3, 'sp4_r_v_b_3')
// (4, 4, 'sp4_r_v_b_43')
// (4, 5, 'sp4_r_v_b_30')
// (4, 6, 'local_g3_3')
// (4, 6, 'lutff_1/in_1')
// (4, 6, 'sp4_h_r_10')
// (4, 6, 'sp4_r_v_b_19')
// (4, 6, 'sp4_v_t_41')
// (4, 7, 'sp4_h_r_43')
// (4, 7, 'sp4_r_v_b_6')
// (4, 7, 'sp4_v_b_41')
// (4, 8, 'sp4_v_b_28')
// (4, 9, 'sp4_v_b_17')
// (4, 10, 'sp4_v_b_4')
// (4, 17, 'sp4_h_r_18')
// (5, 0, 'span4_vert_24')
// (5, 0, 'span4_vert_27')
// (5, 1, 'sp4_v_b_24')
// (5, 1, 'sp4_v_b_27')
// (5, 2, 'sp4_v_b_13')
// (5, 2, 'sp4_v_b_14')
// (5, 3, 'sp12_h_r_7')
// (5, 3, 'sp4_h_r_0')
// (5, 3, 'sp4_h_r_10')
// (5, 3, 'sp4_h_r_33')
// (5, 3, 'sp4_v_b_0')
// (5, 3, 'sp4_v_b_3')
// (5, 3, 'sp4_v_t_43')
// (5, 4, 'sp4_v_b_43')
// (5, 5, 'local_g3_6')
// (5, 5, 'lutff_3/in_0')
// (5, 5, 'sp4_v_b_30')
// (5, 6, 'sp4_h_r_23')
// (5, 6, 'sp4_v_b_19')
// (5, 7, 'sp4_h_l_43')
// (5, 7, 'sp4_h_r_6')
// (5, 7, 'sp4_v_b_6')
// (5, 17, 'sp4_h_r_31')
// (6, 3, 'sp12_h_r_8')
// (6, 3, 'sp4_h_r_13')
// (6, 3, 'sp4_h_r_23')
// (6, 3, 'sp4_h_r_44')
// (6, 6, 'sp4_h_r_34')
// (6, 7, 'sp4_h_r_19')
// (6, 14, 'sp4_r_v_b_42')
// (6, 15, 'sp4_r_v_b_31')
// (6, 16, 'sp4_r_v_b_18')
// (6, 17, 'sp4_h_r_42')
// (6, 17, 'sp4_r_v_b_7')
// (7, 3, 'sp12_h_r_11')
// (7, 3, 'sp4_h_l_44')
// (7, 3, 'sp4_h_r_24')
// (7, 3, 'sp4_h_r_34')
// (7, 3, 'sp4_h_r_9')
// (7, 6, 'sp4_h_r_47')
// (7, 7, 'sp4_h_r_30')
// (7, 7, 'sp4_r_v_b_36')
// (7, 8, 'sp4_r_v_b_25')
// (7, 9, 'sp4_r_v_b_12')
// (7, 10, 'sp4_r_v_b_1')
// (7, 13, 'sp4_h_r_1')
// (7, 13, 'sp4_v_t_42')
// (7, 14, 'sp4_v_b_42')
// (7, 15, 'sp4_v_b_31')
// (7, 16, 'sp4_v_b_18')
// (7, 17, 'sp4_h_l_42')
// (7, 17, 'sp4_v_b_7')
// (8, 3, 'sp12_h_r_12')
// (8, 3, 'sp4_h_r_20')
// (8, 3, 'sp4_h_r_37')
// (8, 3, 'sp4_h_r_47')
// (8, 4, 'local_g1_1')
// (8, 4, 'lutff_0/in_2')
// (8, 4, 'sp4_h_r_1')
// (8, 4, 'sp4_r_v_b_43')
// (8, 5, 'sp4_r_v_b_30')
// (8, 6, 'sp4_h_l_47')
// (8, 6, 'sp4_h_r_7')
// (8, 6, 'sp4_r_v_b_19')
// (8, 6, 'sp4_v_t_36')
// (8, 7, 'sp4_h_r_43')
// (8, 7, 'sp4_r_v_b_6')
// (8, 7, 'sp4_v_b_36')
// (8, 8, 'sp4_v_b_25')
// (8, 9, 'local_g0_4')
// (8, 9, 'lutff_6/in_2')
// (8, 9, 'sp4_v_b_12')
// (8, 10, 'sp4_v_b_1')
// (8, 13, 'local_g0_0')
// (8, 13, 'lutff_2/in_0')
// (8, 13, 'sp12_h_r_0')
// (8, 13, 'sp4_h_r_12')
// (8, 14, 'sp4_r_v_b_44')
// (8, 15, 'sp4_r_v_b_33')
// (8, 16, 'sp4_r_v_b_20')
// (8, 17, 'sp4_r_v_b_9')
// (8, 18, 'sp4_r_v_b_37')
// (8, 19, 'sp4_r_v_b_24')
// (8, 20, 'sp4_r_v_b_13')
// (8, 21, 'sp4_r_v_b_0')
// (9, 3, 'local_g0_7')
// (9, 3, 'lutff_2/in_1')
// (9, 3, 'sp12_h_r_15')
// (9, 3, 'sp4_h_l_37')
// (9, 3, 'sp4_h_l_47')
// (9, 3, 'sp4_h_r_0')
// (9, 3, 'sp4_h_r_33')
// (9, 3, 'sp4_h_r_7')
// (9, 3, 'sp4_v_t_43')
// (9, 4, 'local_g1_4')
// (9, 4, 'lutff_6/in_1')
// (9, 4, 'sp4_h_r_12')
// (9, 4, 'sp4_v_b_43')
// (9, 5, 'sp4_v_b_30')
// (9, 6, 'sp4_h_r_18')
// (9, 6, 'sp4_v_b_19')
// (9, 7, 'sp4_h_l_43')
// (9, 7, 'sp4_v_b_6')
// (9, 13, 'sp12_h_r_3')
// (9, 13, 'sp4_h_r_25')
// (9, 13, 'sp4_h_r_3')
// (9, 13, 'sp4_v_t_44')
// (9, 14, 'sp4_v_b_44')
// (9, 15, 'sp4_v_b_33')
// (9, 16, 'sp4_v_b_20')
// (9, 17, 'sp4_v_b_9')
// (9, 17, 'sp4_v_t_37')
// (9, 18, 'sp4_h_r_9')
// (9, 18, 'sp4_v_b_37')
// (9, 19, 'sp4_v_b_24')
// (9, 20, 'sp4_v_b_13')
// (9, 21, 'local_g1_0')
// (9, 21, 'lutff_7/in_2')
// (9, 21, 'sp4_v_b_0')
// (10, 1, 'local_g0_1')
// (10, 1, 'lutff_7/in_0')
// (10, 1, 'sp4_r_v_b_25')
// (10, 1, 'sp4_r_v_b_34')
// (10, 2, 'local_g3_7')
// (10, 2, 'lutff_5/in_1')
// (10, 2, 'sp4_r_v_b_12')
// (10, 2, 'sp4_r_v_b_23')
// (10, 3, 'sp12_h_r_16')
// (10, 3, 'sp4_h_r_13')
// (10, 3, 'sp4_h_r_18')
// (10, 3, 'sp4_h_r_44')
// (10, 3, 'sp4_r_v_b_1')
// (10, 3, 'sp4_r_v_b_10')
// (10, 4, 'sp4_h_r_25')
// (10, 6, 'sp4_h_r_31')
// (10, 13, 'sp12_h_r_4')
// (10, 13, 'sp4_h_r_14')
// (10, 13, 'sp4_h_r_36')
// (10, 14, 'sp4_r_v_b_46')
// (10, 15, 'sp4_r_v_b_35')
// (10, 16, 'sp4_r_v_b_22')
// (10, 17, 'sp4_r_v_b_11')
// (10, 18, 'local_g1_4')
// (10, 18, 'lutff_5/in_2')
// (10, 18, 'sp4_h_r_20')
// (10, 18, 'sp4_r_v_b_42')
// (10, 19, 'sp4_r_v_b_31')
// (10, 20, 'local_g3_2')
// (10, 20, 'lutff_1/in_0')
// (10, 20, 'sp4_r_v_b_18')
// (10, 21, 'sp4_r_v_b_7')
// (11, 0, 'span4_vert_25')
// (11, 0, 'span4_vert_34')
// (11, 1, 'sp4_v_b_25')
// (11, 1, 'sp4_v_b_34')
// (11, 2, 'sp4_v_b_12')
// (11, 2, 'sp4_v_b_23')
// (11, 3, 'sp12_h_r_19')
// (11, 3, 'sp4_h_l_44')
// (11, 3, 'sp4_h_r_1')
// (11, 3, 'sp4_h_r_24')
// (11, 3, 'sp4_h_r_31')
// (11, 3, 'sp4_h_r_5')
// (11, 3, 'sp4_r_v_b_44')
// (11, 3, 'sp4_v_b_1')
// (11, 3, 'sp4_v_b_10')
// (11, 4, 'sp4_h_r_36')
// (11, 4, 'sp4_r_v_b_33')
// (11, 5, 'sp4_r_v_b_20')
// (11, 6, 'local_g2_1')
// (11, 6, 'lutff_7/in_0')
// (11, 6, 'sp4_h_r_42')
// (11, 6, 'sp4_r_v_b_9')
// (11, 7, 'sp4_r_v_b_47')
// (11, 8, 'sp4_r_v_b_34')
// (11, 9, 'sp4_r_v_b_23')
// (11, 10, 'sp4_r_v_b_10')
// (11, 11, 'sp4_r_v_b_43')
// (11, 12, 'sp4_r_v_b_30')
// (11, 13, 'sp12_h_r_7')
// (11, 13, 'sp4_h_l_36')
// (11, 13, 'sp4_h_r_27')
// (11, 13, 'sp4_h_r_5')
// (11, 13, 'sp4_r_v_b_19')
// (11, 13, 'sp4_v_t_46')
// (11, 14, 'sp4_r_v_b_6')
// (11, 14, 'sp4_v_b_46')
// (11, 15, 'sp4_r_v_b_39')
// (11, 15, 'sp4_v_b_35')
// (11, 16, 'sp4_r_v_b_26')
// (11, 16, 'sp4_v_b_22')
// (11, 17, 'local_g2_7')
// (11, 17, 'lutff_0/in_3')
// (11, 17, 'sp4_r_v_b_15')
// (11, 17, 'sp4_v_b_11')
// (11, 17, 'sp4_v_t_42')
// (11, 18, 'sp4_h_r_33')
// (11, 18, 'sp4_r_v_b_2')
// (11, 18, 'sp4_v_b_42')
// (11, 19, 'sp4_v_b_31')
// (11, 20, 'sp4_v_b_18')
// (11, 21, 'sp4_v_b_7')
// (12, 2, 'sp4_v_t_44')
// (12, 3, 'sp12_h_r_20')
// (12, 3, 'sp4_h_r_12')
// (12, 3, 'sp4_h_r_16')
// (12, 3, 'sp4_h_r_37')
// (12, 3, 'sp4_h_r_42')
// (12, 3, 'sp4_v_b_44')
// (12, 4, 'sp4_h_l_36')
// (12, 4, 'sp4_h_r_5')
// (12, 4, 'sp4_r_v_b_47')
// (12, 4, 'sp4_v_b_33')
// (12, 5, 'sp4_r_v_b_34')
// (12, 5, 'sp4_v_b_20')
// (12, 6, 'sp4_h_l_42')
// (12, 6, 'sp4_h_r_4')
// (12, 6, 'sp4_r_v_b_23')
// (12, 6, 'sp4_v_b_9')
// (12, 6, 'sp4_v_t_47')
// (12, 7, 'sp4_r_v_b_10')
// (12, 7, 'sp4_v_b_47')
// (12, 8, 'sp4_v_b_34')
// (12, 9, 'sp4_v_b_23')
// (12, 10, 'local_g0_2')
// (12, 10, 'lutff_7/in_1')
// (12, 10, 'sp4_v_b_10')
// (12, 10, 'sp4_v_t_43')
// (12, 11, 'sp4_v_b_43')
// (12, 12, 'sp4_v_b_30')
// (12, 13, 'sp12_h_r_8')
// (12, 13, 'sp4_h_r_16')
// (12, 13, 'sp4_h_r_38')
// (12, 13, 'sp4_v_b_19')
// (12, 14, 'sp4_v_b_6')
// (12, 14, 'sp4_v_t_39')
// (12, 15, 'sp4_v_b_39')
// (12, 16, 'sp4_v_b_26')
// (12, 17, 'sp4_v_b_15')
// (12, 18, 'sp4_h_r_44')
// (12, 18, 'sp4_v_b_2')
// (13, 3, 'sp12_h_r_23')
// (13, 3, 'sp4_h_l_37')
// (13, 3, 'sp4_h_l_42')
// (13, 3, 'sp4_h_r_1')
// (13, 3, 'sp4_h_r_25')
// (13, 3, 'sp4_h_r_29')
// (13, 3, 'sp4_h_r_4')
// (13, 3, 'sp4_v_t_47')
// (13, 4, 'sp4_h_r_11')
// (13, 4, 'sp4_h_r_16')
// (13, 4, 'sp4_v_b_47')
// (13, 5, 'local_g3_2')
// (13, 5, 'lutff_5/in_0')
// (13, 5, 'sp4_v_b_34')
// (13, 6, 'sp4_h_r_17')
// (13, 6, 'sp4_v_b_23')
// (13, 7, 'sp4_v_b_10')
// (13, 13, 'sp12_h_r_11')
// (13, 13, 'sp4_h_l_38')
// (13, 13, 'sp4_h_r_29')
// (13, 18, 'sp4_h_l_44')
// (13, 18, 'sp4_h_r_6')
// (14, 1, 'sp4_r_v_b_29')
// (14, 2, 'sp4_r_v_b_16')
// (14, 3, 'local_g1_4')
// (14, 3, 'lutff_1/in_0')
// (14, 3, 'sp12_h_l_23')
// (14, 3, 'sp12_h_r_0')
// (14, 3, 'sp4_h_r_12')
// (14, 3, 'sp4_h_r_17')
// (14, 3, 'sp4_h_r_36')
// (14, 3, 'sp4_h_r_40')
// (14, 3, 'sp4_r_v_b_5')
// (14, 4, 'local_g0_6')
// (14, 4, 'lutff_1/in_3')
// (14, 4, 'sp4_h_r_22')
// (14, 4, 'sp4_h_r_29')
// (14, 4, 'sp4_r_v_b_46')
// (14, 5, 'local_g0_0')
// (14, 5, 'lutff_3/in_1')
// (14, 5, 'sp4_r_v_b_35')
// (14, 6, 'sp4_h_r_28')
// (14, 6, 'sp4_r_v_b_22')
// (14, 7, 'sp4_r_v_b_11')
// (14, 13, 'sp12_h_r_12')
// (14, 13, 'sp4_h_r_40')
// (14, 18, 'sp4_h_r_19')
// (15, 0, 'span4_vert_29')
// (15, 1, 'sp4_v_b_29')
// (15, 2, 'local_g0_0')
// (15, 2, 'lutff_4/in_0')
// (15, 2, 'sp4_v_b_16')
// (15, 3, 'local_g1_3')
// (15, 3, 'lutff_7/in_1')
// (15, 3, 'sp12_h_r_3')
// (15, 3, 'sp4_h_l_36')
// (15, 3, 'sp4_h_l_40')
// (15, 3, 'sp4_h_r_25')
// (15, 3, 'sp4_h_r_28')
// (15, 3, 'sp4_h_r_5')
// (15, 3, 'sp4_v_b_5')
// (15, 3, 'sp4_v_t_46')
// (15, 4, 'sp4_h_r_35')
// (15, 4, 'sp4_h_r_40')
// (15, 4, 'sp4_v_b_46')
// (15, 5, 'sp4_v_b_35')
// (15, 6, 'sp4_h_r_41')
// (15, 6, 'sp4_v_b_22')
// (15, 7, 'sp4_v_b_11')
// (15, 13, 'sp12_h_r_15')
// (15, 13, 'sp4_h_l_40')
// (15, 18, 'sp4_h_r_30')
// (16, 3, 'sp12_h_r_4')
// (16, 3, 'sp4_h_r_16')
// (16, 3, 'sp4_h_r_36')
// (16, 3, 'sp4_h_r_41')
// (16, 4, 'sp4_h_l_40')
// (16, 4, 'sp4_h_r_46')
// (16, 4, 'sp4_h_r_9')
// (16, 6, 'sp4_h_l_41')
// (16, 6, 'sp4_h_r_1')
// (16, 7, 'sp4_r_v_b_40')
// (16, 8, 'sp4_r_v_b_29')
// (16, 9, 'sp4_r_v_b_16')
// (16, 10, 'sp4_r_v_b_5')
// (16, 11, 'sp4_r_v_b_36')
// (16, 12, 'sp4_r_v_b_25')
// (16, 13, 'sp12_h_r_16')
// (16, 13, 'sp4_r_v_b_12')
// (16, 14, 'sp4_r_v_b_1')
// (16, 15, 'sp4_r_v_b_36')
// (16, 16, 'sp4_r_v_b_25')
// (16, 17, 'sp4_r_v_b_12')
// (16, 18, 'sp4_h_r_43')
// (16, 18, 'sp4_r_v_b_1')
// (17, 3, 'sp12_h_r_7')
// (17, 3, 'sp4_h_l_36')
// (17, 3, 'sp4_h_l_41')
// (17, 3, 'sp4_h_r_1')
// (17, 3, 'sp4_h_r_29')
// (17, 4, 'sp4_h_l_46')
// (17, 4, 'sp4_h_r_20')
// (17, 4, 'sp4_h_r_8')
// (17, 6, 'sp4_h_r_12')
// (17, 6, 'sp4_h_r_5')
// (17, 6, 'sp4_v_t_40')
// (17, 7, 'sp4_v_b_40')
// (17, 8, 'sp4_v_b_29')
// (17, 9, 'sp4_v_b_16')
// (17, 10, 'sp4_v_b_5')
// (17, 10, 'sp4_v_t_36')
// (17, 11, 'sp4_v_b_36')
// (17, 12, 'sp4_v_b_25')
// (17, 13, 'sp12_h_r_19')
// (17, 13, 'sp4_v_b_12')
// (17, 14, 'sp4_v_b_1')
// (17, 14, 'sp4_v_t_36')
// (17, 15, 'sp4_v_b_36')
// (17, 16, 'sp4_v_b_25')
// (17, 17, 'sp4_v_b_12')
// (17, 18, 'sp4_h_l_43')
// (17, 18, 'sp4_v_b_1')
// (18, 3, 'sp12_h_r_8')
// (18, 3, 'sp4_h_r_12')
// (18, 3, 'sp4_h_r_40')
// (18, 4, 'sp4_h_r_21')
// (18, 4, 'sp4_h_r_33')
// (18, 6, 'sp4_h_r_16')
// (18, 6, 'sp4_h_r_25')
// (18, 13, 'sp12_h_r_20')
// (19, 1, 'sp4_r_v_b_44')
// (19, 2, 'neigh_op_tnr_2')
// (19, 2, 'sp4_r_v_b_33')
// (19, 3, 'neigh_op_rgt_2')
// (19, 3, 'sp12_h_r_11')
// (19, 3, 'sp4_h_l_40')
// (19, 3, 'sp4_h_r_25')
// (19, 3, 'sp4_h_r_9')
// (19, 3, 'sp4_r_v_b_20')
// (19, 3, 'sp4_r_v_b_36')
// (19, 4, 'neigh_op_bnr_2')
// (19, 4, 'sp4_h_r_32')
// (19, 4, 'sp4_h_r_44')
// (19, 4, 'sp4_r_v_b_25')
// (19, 4, 'sp4_r_v_b_9')
// (19, 5, 'sp4_r_v_b_12')
// (19, 6, 'sp4_h_r_29')
// (19, 6, 'sp4_h_r_36')
// (19, 6, 'sp4_r_v_b_1')
// (19, 13, 'sp12_h_r_23')
// (20, 0, 'span4_vert_44')
// (20, 1, 'sp12_v_t_23')
// (20, 1, 'sp4_r_v_b_45')
// (20, 1, 'sp4_v_b_44')
// (20, 2, 'neigh_op_top_2')
// (20, 2, 'sp12_v_b_23')
// (20, 2, 'sp4_r_v_b_32')
// (20, 2, 'sp4_v_b_33')
// (20, 2, 'sp4_v_t_36')
// (20, 3, 'lutff_2/out')
// (20, 3, 'sp12_h_r_12')
// (20, 3, 'sp12_v_b_20')
// (20, 3, 'sp4_h_r_20')
// (20, 3, 'sp4_h_r_36')
// (20, 3, 'sp4_r_v_b_21')
// (20, 3, 'sp4_r_v_b_37')
// (20, 3, 'sp4_v_b_20')
// (20, 3, 'sp4_v_b_36')
// (20, 4, 'neigh_op_bot_2')
// (20, 4, 'sp12_v_b_19')
// (20, 4, 'sp4_h_l_44')
// (20, 4, 'sp4_h_r_45')
// (20, 4, 'sp4_r_v_b_24')
// (20, 4, 'sp4_r_v_b_8')
// (20, 4, 'sp4_v_b_25')
// (20, 4, 'sp4_v_b_9')
// (20, 5, 'sp12_v_b_16')
// (20, 5, 'sp4_r_v_b_13')
// (20, 5, 'sp4_v_b_12')
// (20, 6, 'sp12_v_b_15')
// (20, 6, 'sp4_h_l_36')
// (20, 6, 'sp4_h_r_40')
// (20, 6, 'sp4_r_v_b_0')
// (20, 6, 'sp4_v_b_1')
// (20, 7, 'sp12_v_b_12')
// (20, 8, 'sp12_v_b_11')
// (20, 9, 'sp12_v_b_8')
// (20, 10, 'sp12_v_b_7')
// (20, 11, 'sp12_v_b_4')
// (20, 12, 'sp12_v_b_3')
// (20, 13, 'sp12_h_l_23')
// (20, 13, 'sp12_v_b_0')
// (21, 0, 'span4_vert_45')
// (21, 1, 'sp4_v_b_45')
// (21, 2, 'neigh_op_tnl_2')
// (21, 2, 'sp4_v_b_32')
// (21, 2, 'sp4_v_t_37')
// (21, 3, 'neigh_op_lft_2')
// (21, 3, 'sp12_h_r_15')
// (21, 3, 'sp4_h_l_36')
// (21, 3, 'sp4_h_r_33')
// (21, 3, 'sp4_v_b_21')
// (21, 3, 'sp4_v_b_37')
// (21, 4, 'neigh_op_bnl_2')
// (21, 4, 'sp4_h_l_45')
// (21, 4, 'sp4_v_b_24')
// (21, 4, 'sp4_v_b_8')
// (21, 5, 'sp4_v_b_13')
// (21, 6, 'sp4_h_l_40')
// (21, 6, 'sp4_v_b_0')
// (22, 3, 'sp12_h_r_16')
// (22, 3, 'sp4_h_r_44')
// (23, 3, 'sp12_h_r_19')
// (23, 3, 'sp4_h_l_44')
// (24, 3, 'sp12_h_r_20')
// (25, 3, 'sp12_h_r_23')

wire n234;
// (1, 8, 'local_g2_3')
// (1, 8, 'lutff_2/in_1')
// (1, 8, 'neigh_op_tnr_3')
// (1, 9, 'neigh_op_rgt_3')
// (1, 10, 'neigh_op_bnr_3')
// (2, 8, 'neigh_op_top_3')
// (2, 9, 'lutff_3/out')
// (2, 10, 'neigh_op_bot_3')
// (3, 8, 'neigh_op_tnl_3')
// (3, 9, 'neigh_op_lft_3')
// (3, 10, 'neigh_op_bnl_3')

reg n235 = 0;
// (1, 8, 'local_g2_7')
// (1, 8, 'lutff_4/in_1')
// (1, 8, 'lutff_7/in_0')
// (1, 8, 'neigh_op_tnr_7')
// (1, 9, 'neigh_op_rgt_7')
// (1, 10, 'local_g1_7')
// (1, 10, 'lutff_0/in_0')
// (1, 10, 'neigh_op_bnr_7')
// (2, 8, 'neigh_op_top_7')
// (2, 9, 'local_g1_7')
// (2, 9, 'lutff_7/in_1')
// (2, 9, 'lutff_7/out')
// (2, 10, 'local_g0_7')
// (2, 10, 'lutff_6/in_3')
// (2, 10, 'neigh_op_bot_7')
// (3, 8, 'neigh_op_tnl_7')
// (3, 9, 'neigh_op_lft_7')
// (3, 10, 'neigh_op_bnl_7')

wire n236;
// (1, 8, 'lutff_2/cout')
// (1, 8, 'lutff_3/in_3')

wire n237;
// (1, 8, 'lutff_3/cout')
// (1, 8, 'lutff_4/in_3')

wire n238;
// (1, 8, 'neigh_op_tnr_1')
// (1, 9, 'neigh_op_rgt_1')
// (1, 10, 'neigh_op_bnr_1')
// (2, 8, 'local_g0_1')
// (2, 8, 'lutff_7/in_0')
// (2, 8, 'neigh_op_top_1')
// (2, 9, 'lutff_1/out')
// (2, 10, 'neigh_op_bot_1')
// (3, 8, 'local_g2_1')
// (3, 8, 'lutff_5/in_0')
// (3, 8, 'neigh_op_tnl_1')
// (3, 9, 'neigh_op_lft_1')
// (3, 10, 'neigh_op_bnl_1')

wire n239;
// (1, 8, 'neigh_op_tnr_2')
// (1, 9, 'neigh_op_rgt_2')
// (1, 10, 'neigh_op_bnr_2')
// (2, 8, 'neigh_op_top_2')
// (2, 9, 'lutff_2/out')
// (2, 10, 'neigh_op_bot_2')
// (3, 8, 'local_g3_2')
// (3, 8, 'lutff_7/in_0')
// (3, 8, 'neigh_op_tnl_2')
// (3, 9, 'neigh_op_lft_2')
// (3, 10, 'neigh_op_bnl_2')

wire n240;
// (1, 8, 'neigh_op_tnr_4')
// (1, 9, 'local_g2_4')
// (1, 9, 'lutff_0/in_0')
// (1, 9, 'lutff_3/in_1')
// (1, 9, 'neigh_op_rgt_4')
// (1, 10, 'neigh_op_bnr_4')
// (2, 8, 'local_g0_4')
// (2, 8, 'local_g1_4')
// (2, 8, 'lutff_2/in_0')
// (2, 8, 'lutff_3/in_0')
// (2, 8, 'lutff_4/in_1')
// (2, 8, 'neigh_op_top_4')
// (2, 9, 'lutff_4/out')
// (2, 10, 'neigh_op_bot_4')
// (3, 8, 'neigh_op_tnl_4')
// (3, 9, 'neigh_op_lft_4')
// (3, 10, 'neigh_op_bnl_4')

wire n241;
// (1, 8, 'neigh_op_tnr_5')
// (1, 9, 'neigh_op_rgt_5')
// (1, 10, 'neigh_op_bnr_5')
// (2, 8, 'neigh_op_top_5')
// (2, 9, 'local_g0_5')
// (2, 9, 'lutff_5/out')
// (2, 9, 'lutff_6/in_3')
// (2, 10, 'neigh_op_bot_5')
// (3, 8, 'neigh_op_tnl_5')
// (3, 9, 'neigh_op_lft_5')
// (3, 10, 'neigh_op_bnl_5')

wire n242;
// (1, 8, 'neigh_op_tnr_6')
// (1, 9, 'neigh_op_rgt_6')
// (1, 10, 'local_g1_6')
// (1, 10, 'lutff_0/in_1')
// (1, 10, 'neigh_op_bnr_6')
// (2, 8, 'neigh_op_top_6')
// (2, 8, 'sp4_r_v_b_40')
// (2, 9, 'lutff_6/out')
// (2, 9, 'sp4_r_v_b_29')
// (2, 10, 'neigh_op_bot_6')
// (2, 10, 'sp4_r_v_b_16')
// (2, 11, 'local_g1_5')
// (2, 11, 'lutff_3/in_3')
// (2, 11, 'sp4_r_v_b_5')
// (3, 7, 'sp4_v_t_40')
// (3, 8, 'neigh_op_tnl_6')
// (3, 8, 'sp4_v_b_40')
// (3, 9, 'neigh_op_lft_6')
// (3, 9, 'sp4_v_b_29')
// (3, 10, 'neigh_op_bnl_6')
// (3, 10, 'sp4_v_b_16')
// (3, 11, 'sp4_v_b_5')

wire n243;
// (1, 8, 'sp4_r_v_b_37')
// (1, 9, 'sp4_r_v_b_24')
// (1, 10, 'sp4_r_v_b_13')
// (1, 11, 'sp4_r_v_b_0')
// (1, 12, 'sp4_r_v_b_37')
// (1, 13, 'sp4_r_v_b_24')
// (1, 14, 'sp4_r_v_b_13')
// (1, 15, 'sp4_r_v_b_0')
// (2, 7, 'sp4_v_t_37')
// (2, 8, 'sp4_v_b_37')
// (2, 9, 'sp4_v_b_24')
// (2, 10, 'local_g1_5')
// (2, 10, 'lutff_5/in_3')
// (2, 10, 'sp4_v_b_13')
// (2, 11, 'local_g0_0')
// (2, 11, 'lutff_0/in_2')
// (2, 11, 'sp4_h_r_0')
// (2, 11, 'sp4_v_b_0')
// (2, 11, 'sp4_v_t_37')
// (2, 12, 'sp4_v_b_37')
// (2, 13, 'local_g3_0')
// (2, 13, 'lutff_2/in_1')
// (2, 13, 'sp4_v_b_24')
// (2, 14, 'sp4_v_b_13')
// (2, 15, 'sp4_v_b_0')
// (3, 10, 'neigh_op_tnr_4')
// (3, 11, 'neigh_op_rgt_4')
// (3, 11, 'sp4_h_r_13')
// (3, 12, 'neigh_op_bnr_4')
// (4, 10, 'neigh_op_top_4')
// (4, 11, 'local_g0_4')
// (4, 11, 'lutff_1/in_3')
// (4, 11, 'lutff_4/out')
// (4, 11, 'sp4_h_r_24')
// (4, 12, 'neigh_op_bot_4')
// (5, 10, 'neigh_op_tnl_4')
// (5, 11, 'neigh_op_lft_4')
// (5, 11, 'sp4_h_r_37')
// (5, 12, 'neigh_op_bnl_4')
// (6, 11, 'sp4_h_l_37')

reg n244 = 0;
// (1, 9, 'neigh_op_tnr_0')
// (1, 9, 'sp4_r_v_b_45')
// (1, 10, 'neigh_op_rgt_0')
// (1, 10, 'sp4_r_v_b_32')
// (1, 11, 'neigh_op_bnr_0')
// (1, 11, 'sp4_r_v_b_21')
// (1, 12, 'local_g2_0')
// (1, 12, 'lutff_1/in_1')
// (1, 12, 'sp4_r_v_b_8')
// (1, 13, 'sp4_r_v_b_45')
// (1, 14, 'local_g2_0')
// (1, 14, 'lutff_1/in_3')
// (1, 14, 'sp4_r_v_b_32')
// (1, 15, 'sp4_r_v_b_21')
// (1, 16, 'sp4_r_v_b_8')
// (2, 8, 'sp4_v_t_45')
// (2, 9, 'neigh_op_top_0')
// (2, 9, 'sp4_v_b_45')
// (2, 10, 'local_g2_0')
// (2, 10, 'lutff_0/in_0')
// (2, 10, 'lutff_0/out')
// (2, 10, 'sp4_v_b_32')
// (2, 11, 'neigh_op_bot_0')
// (2, 11, 'sp4_v_b_21')
// (2, 12, 'sp4_v_b_8')
// (2, 12, 'sp4_v_t_45')
// (2, 13, 'sp4_v_b_45')
// (2, 14, 'sp4_v_b_32')
// (2, 15, 'sp4_v_b_21')
// (2, 16, 'sp4_v_b_8')
// (3, 9, 'neigh_op_tnl_0')
// (3, 10, 'neigh_op_lft_0')
// (3, 11, 'neigh_op_bnl_0')

wire n245;
// (1, 9, 'neigh_op_tnr_2')
// (1, 10, 'neigh_op_rgt_2')
// (1, 11, 'local_g0_2')
// (1, 11, 'lutff_global/cen')
// (1, 11, 'neigh_op_bnr_2')
// (2, 9, 'neigh_op_top_2')
// (2, 10, 'lutff_2/out')
// (2, 11, 'neigh_op_bot_2')
// (3, 9, 'neigh_op_tnl_2')
// (3, 10, 'neigh_op_lft_2')
// (3, 11, 'neigh_op_bnl_2')

reg n246 = 0;
// (1, 9, 'neigh_op_tnr_3')
// (1, 10, 'neigh_op_rgt_3')
// (1, 10, 'sp4_r_v_b_38')
// (1, 11, 'neigh_op_bnr_3')
// (1, 11, 'sp4_r_v_b_27')
// (1, 12, 'local_g2_6')
// (1, 12, 'lutff_2/in_0')
// (1, 12, 'sp4_r_v_b_14')
// (1, 13, 'sp4_r_v_b_3')
// (2, 9, 'neigh_op_top_3')
// (2, 9, 'sp4_v_t_38')
// (2, 10, 'local_g2_3')
// (2, 10, 'lutff_3/in_0')
// (2, 10, 'lutff_3/out')
// (2, 10, 'sp4_v_b_38')
// (2, 11, 'neigh_op_bot_3')
// (2, 11, 'sp4_v_b_27')
// (2, 12, 'sp4_v_b_14')
// (2, 13, 'sp4_v_b_3')
// (3, 9, 'neigh_op_tnl_3')
// (3, 10, 'neigh_op_lft_3')
// (3, 11, 'neigh_op_bnl_3')

reg n247 = 0;
// (1, 9, 'neigh_op_tnr_4')
// (1, 9, 'sp4_r_v_b_37')
// (1, 10, 'neigh_op_rgt_4')
// (1, 10, 'sp4_r_v_b_24')
// (1, 11, 'local_g0_4')
// (1, 11, 'lutff_6/in_2')
// (1, 11, 'neigh_op_bnr_4')
// (1, 11, 'sp4_r_v_b_13')
// (1, 12, 'local_g1_0')
// (1, 12, 'lutff_7/in_2')
// (1, 12, 'sp4_r_v_b_0')
// (2, 8, 'sp4_v_t_37')
// (2, 9, 'neigh_op_top_4')
// (2, 9, 'sp4_v_b_37')
// (2, 10, 'lutff_4/out')
// (2, 10, 'sp4_v_b_24')
// (2, 11, 'neigh_op_bot_4')
// (2, 11, 'sp4_v_b_13')
// (2, 12, 'sp4_v_b_0')
// (3, 9, 'neigh_op_tnl_4')
// (3, 10, 'neigh_op_lft_4')
// (3, 11, 'neigh_op_bnl_4')

wire n248;
// (1, 9, 'neigh_op_tnr_7')
// (1, 10, 'neigh_op_rgt_7')
// (1, 11, 'neigh_op_bnr_7')
// (2, 8, 'sp4_r_v_b_39')
// (2, 9, 'neigh_op_top_7')
// (2, 9, 'sp4_r_v_b_26')
// (2, 10, 'lutff_7/out')
// (2, 10, 'sp4_r_v_b_15')
// (2, 11, 'neigh_op_bot_7')
// (2, 11, 'sp4_r_v_b_2')
// (3, 7, 'sp4_v_t_39')
// (3, 8, 'sp4_v_b_39')
// (3, 9, 'neigh_op_tnl_7')
// (3, 9, 'sp4_v_b_26')
// (3, 10, 'neigh_op_lft_7')
// (3, 10, 'sp4_v_b_15')
// (3, 11, 'neigh_op_bnl_7')
// (3, 11, 'sp4_h_r_8')
// (3, 11, 'sp4_v_b_2')
// (4, 11, 'local_g0_5')
// (4, 11, 'lutff_2/in_1')
// (4, 11, 'sp4_h_r_21')
// (5, 11, 'sp4_h_r_32')
// (6, 11, 'sp4_h_r_45')
// (7, 11, 'sp4_h_l_45')

wire n249;
// (1, 9, 'sp4_r_v_b_39')
// (1, 9, 'sp4_r_v_b_40')
// (1, 10, 'sp4_h_r_5')
// (1, 10, 'sp4_r_v_b_26')
// (1, 10, 'sp4_r_v_b_29')
// (1, 11, 'sp4_r_v_b_15')
// (1, 11, 'sp4_r_v_b_16')
// (1, 12, 'sp4_r_v_b_2')
// (1, 12, 'sp4_r_v_b_5')
// (1, 13, 'local_g2_7')
// (1, 13, 'lutff_5/in_0')
// (1, 13, 'sp4_r_v_b_39')
// (1, 14, 'sp4_r_v_b_26')
// (1, 15, 'sp4_r_v_b_15')
// (1, 16, 'sp4_r_v_b_2')
// (1, 17, 'sp4_r_v_b_39')
// (1, 18, 'sp4_r_v_b_26')
// (1, 19, 'sp4_r_v_b_15')
// (1, 20, 'sp4_r_v_b_2')
// (2, 8, 'sp4_v_t_39')
// (2, 8, 'sp4_v_t_40')
// (2, 9, 'sp4_v_b_39')
// (2, 9, 'sp4_v_b_40')
// (2, 10, 'local_g0_0')
// (2, 10, 'lutff_2/in_2')
// (2, 10, 'lutff_5/in_1')
// (2, 10, 'sp4_h_r_16')
// (2, 10, 'sp4_v_b_26')
// (2, 10, 'sp4_v_b_29')
// (2, 11, 'local_g1_7')
// (2, 11, 'lutff_7/in_3')
// (2, 11, 'sp4_v_b_15')
// (2, 11, 'sp4_v_b_16')
// (2, 12, 'local_g0_2')
// (2, 12, 'local_g0_5')
// (2, 12, 'lutff_3/in_2')
// (2, 12, 'lutff_6/in_0')
// (2, 12, 'sp4_v_b_2')
// (2, 12, 'sp4_v_b_5')
// (2, 12, 'sp4_v_t_39')
// (2, 13, 'sp4_v_b_39')
// (2, 14, 'sp4_v_b_26')
// (2, 15, 'local_g1_7')
// (2, 15, 'lutff_3/in_3')
// (2, 15, 'sp4_v_b_15')
// (2, 16, 'sp4_h_r_2')
// (2, 16, 'sp4_v_b_2')
// (2, 16, 'sp4_v_t_39')
// (2, 17, 'local_g2_7')
// (2, 17, 'lutff_4/in_1')
// (2, 17, 'sp4_v_b_39')
// (2, 18, 'sp4_v_b_26')
// (2, 19, 'sp4_v_b_15')
// (2, 20, 'local_g1_2')
// (2, 20, 'lutff_6/in_3')
// (2, 20, 'sp4_v_b_2')
// (3, 10, 'sp4_h_r_29')
// (3, 12, 'sp4_r_v_b_38')
// (3, 13, 'sp4_r_v_b_27')
// (3, 14, 'local_g2_6')
// (3, 14, 'lutff_5/in_1')
// (3, 14, 'sp4_r_v_b_14')
// (3, 15, 'local_g2_5')
// (3, 15, 'lutff_1/in_2')
// (3, 15, 'neigh_op_tnr_5')
// (3, 15, 'sp4_r_v_b_3')
// (3, 16, 'local_g2_5')
// (3, 16, 'lutff_5/in_2')
// (3, 16, 'neigh_op_rgt_5')
// (3, 16, 'sp4_h_r_15')
// (3, 16, 'sp4_r_v_b_42')
// (3, 17, 'local_g1_5')
// (3, 17, 'lutff_5/in_3')
// (3, 17, 'neigh_op_bnr_5')
// (3, 17, 'sp4_r_v_b_31')
// (3, 18, 'sp4_r_v_b_18')
// (3, 19, 'sp4_r_v_b_7')
// (4, 10, 'sp4_h_r_40')
// (4, 11, 'local_g3_6')
// (4, 11, 'lutff_1/in_0')
// (4, 11, 'sp4_r_v_b_46')
// (4, 11, 'sp4_v_t_38')
// (4, 12, 'sp4_r_v_b_35')
// (4, 12, 'sp4_v_b_38')
// (4, 13, 'sp4_r_v_b_22')
// (4, 13, 'sp4_v_b_27')
// (4, 14, 'local_g0_6')
// (4, 14, 'lutff_0/in_0')
// (4, 14, 'sp4_r_v_b_11')
// (4, 14, 'sp4_v_b_14')
// (4, 15, 'neigh_op_top_5')
// (4, 15, 'sp4_r_v_b_38')
// (4, 15, 'sp4_v_b_3')
// (4, 15, 'sp4_v_t_42')
// (4, 16, 'local_g3_5')
// (4, 16, 'lutff_0/in_0')
// (4, 16, 'lutff_3/in_3')
// (4, 16, 'lutff_5/out')
// (4, 16, 'lutff_7/in_1')
// (4, 16, 'sp4_h_r_26')
// (4, 16, 'sp4_r_v_b_27')
// (4, 16, 'sp4_v_b_42')
// (4, 17, 'neigh_op_bot_5')
// (4, 17, 'sp4_r_v_b_14')
// (4, 17, 'sp4_v_b_31')
// (4, 18, 'sp4_r_v_b_3')
// (4, 18, 'sp4_v_b_18')
// (4, 19, 'local_g1_7')
// (4, 19, 'lutff_5/in_3')
// (4, 19, 'lutff_6/in_0')
// (4, 19, 'sp4_h_r_7')
// (4, 19, 'sp4_v_b_7')
// (5, 10, 'sp4_h_l_40')
// (5, 10, 'sp4_v_t_46')
// (5, 11, 'sp4_v_b_46')
// (5, 12, 'sp4_v_b_35')
// (5, 13, 'sp4_v_b_22')
// (5, 14, 'local_g1_3')
// (5, 14, 'lutff_1/in_3')
// (5, 14, 'lutff_2/in_2')
// (5, 14, 'lutff_5/in_1')
// (5, 14, 'sp4_h_r_3')
// (5, 14, 'sp4_v_b_11')
// (5, 14, 'sp4_v_t_38')
// (5, 15, 'local_g3_5')
// (5, 15, 'lutff_6/in_0')
// (5, 15, 'neigh_op_tnl_5')
// (5, 15, 'sp4_v_b_38')
// (5, 16, 'local_g0_5')
// (5, 16, 'lutff_2/in_1')
// (5, 16, 'neigh_op_lft_5')
// (5, 16, 'sp4_h_r_39')
// (5, 16, 'sp4_v_b_27')
// (5, 17, 'local_g3_5')
// (5, 17, 'lutff_5/in_3')
// (5, 17, 'neigh_op_bnl_5')
// (5, 17, 'sp4_v_b_14')
// (5, 18, 'sp4_h_r_3')
// (5, 18, 'sp4_v_b_3')
// (5, 19, 'sp4_h_r_18')
// (6, 14, 'sp4_h_r_14')
// (6, 16, 'sp4_h_l_39')
// (6, 16, 'sp4_h_r_5')
// (6, 18, 'sp4_h_r_14')
// (6, 19, 'sp4_h_r_31')
// (7, 14, 'sp4_h_r_27')
// (7, 16, 'sp4_h_r_16')
// (7, 18, 'sp4_h_r_27')
// (7, 19, 'sp4_h_r_42')
// (7, 20, 'sp4_r_v_b_42')
// (7, 21, 'local_g0_7')
// (7, 21, 'lutff_5/in_0')
// (7, 21, 'sp4_r_v_b_31')
// (7, 22, 'sp4_r_v_b_18')
// (7, 23, 'sp4_r_v_b_7')
// (8, 11, 'sp4_r_v_b_44')
// (8, 12, 'sp4_r_v_b_33')
// (8, 13, 'sp4_r_v_b_20')
// (8, 14, 'sp4_h_r_38')
// (8, 14, 'sp4_r_v_b_9')
// (8, 16, 'sp4_h_r_29')
// (8, 18, 'sp4_h_r_38')
// (8, 19, 'sp4_h_l_42')
// (8, 19, 'sp4_r_v_b_38')
// (8, 19, 'sp4_v_t_42')
// (8, 20, 'sp4_r_v_b_27')
// (8, 20, 'sp4_v_b_42')
// (8, 21, 'local_g2_6')
// (8, 21, 'lutff_4/in_0')
// (8, 21, 'sp4_r_v_b_14')
// (8, 21, 'sp4_v_b_31')
// (8, 22, 'sp4_r_v_b_3')
// (8, 22, 'sp4_v_b_18')
// (8, 23, 'sp4_v_b_7')
// (9, 10, 'sp4_v_t_44')
// (9, 11, 'local_g2_4')
// (9, 11, 'lutff_6/in_0')
// (9, 11, 'sp4_v_b_44')
// (9, 12, 'sp4_v_b_33')
// (9, 13, 'sp4_r_v_b_40')
// (9, 13, 'sp4_v_b_20')
// (9, 14, 'sp4_h_l_38')
// (9, 14, 'sp4_r_v_b_29')
// (9, 14, 'sp4_v_b_9')
// (9, 15, 'local_g3_0')
// (9, 15, 'lutff_6/in_3')
// (9, 15, 'sp4_r_v_b_16')
// (9, 16, 'sp4_h_r_40')
// (9, 16, 'sp4_r_v_b_5')
// (9, 18, 'sp4_h_l_38')
// (9, 18, 'sp4_v_t_38')
// (9, 19, 'sp4_v_b_38')
// (9, 20, 'sp4_v_b_27')
// (9, 21, 'sp4_v_b_14')
// (9, 22, 'sp4_v_b_3')
// (10, 12, 'sp4_v_t_40')
// (10, 13, 'sp4_v_b_40')
// (10, 14, 'sp4_v_b_29')
// (10, 15, 'sp4_v_b_16')
// (10, 16, 'sp4_h_l_40')
// (10, 16, 'sp4_v_b_5')

wire n250;
// (1, 9, 'sp4_r_v_b_43')
// (1, 10, 'sp4_r_v_b_30')
// (1, 11, 'neigh_op_tnr_3')
// (1, 11, 'sp4_r_v_b_19')
// (1, 12, 'neigh_op_rgt_3')
// (1, 12, 'sp4_r_v_b_6')
// (1, 13, 'neigh_op_bnr_3')
// (2, 8, 'sp4_v_t_43')
// (2, 9, 'sp4_v_b_43')
// (2, 10, 'local_g2_6')
// (2, 10, 'lutff_3/in_3')
// (2, 10, 'sp4_v_b_30')
// (2, 11, 'neigh_op_top_3')
// (2, 11, 'sp4_v_b_19')
// (2, 12, 'lutff_3/out')
// (2, 12, 'sp4_v_b_6')
// (2, 13, 'neigh_op_bot_3')
// (3, 11, 'neigh_op_tnl_3')
// (3, 12, 'neigh_op_lft_3')
// (3, 13, 'neigh_op_bnl_3')

reg n251 = 0;
// (1, 10, 'neigh_op_tnr_0')
// (1, 11, 'neigh_op_rgt_0')
// (1, 12, 'neigh_op_bnr_0')
// (2, 10, 'local_g1_0')
// (2, 10, 'lutff_1/in_0')
// (2, 10, 'neigh_op_top_0')
// (2, 11, 'local_g3_0')
// (2, 11, 'lutff_0/in_1')
// (2, 11, 'lutff_0/out')
// (2, 12, 'neigh_op_bot_0')
// (3, 10, 'neigh_op_tnl_0')
// (3, 11, 'neigh_op_lft_0')
// (3, 12, 'neigh_op_bnl_0')

reg n252 = 0;
// (1, 10, 'neigh_op_tnr_1')
// (1, 10, 'sp4_r_v_b_47')
// (1, 11, 'neigh_op_rgt_1')
// (1, 11, 'sp4_r_v_b_34')
// (1, 12, 'local_g0_1')
// (1, 12, 'lutff_0/in_1')
// (1, 12, 'lutff_4/in_1')
// (1, 12, 'neigh_op_bnr_1')
// (1, 12, 'sp4_r_v_b_23')
// (1, 13, 'sp4_r_v_b_10')
// (1, 14, 'sp4_r_v_b_43')
// (1, 15, 'sp4_r_v_b_30')
// (1, 16, 'sp4_r_v_b_19')
// (1, 17, 'sp4_r_v_b_6')
// (2, 9, 'sp4_v_t_47')
// (2, 10, 'neigh_op_top_1')
// (2, 10, 'sp4_v_b_47')
// (2, 11, 'lutff_1/out')
// (2, 11, 'sp4_v_b_34')
// (2, 12, 'neigh_op_bot_1')
// (2, 12, 'sp4_v_b_23')
// (2, 13, 'sp4_h_r_4')
// (2, 13, 'sp4_v_b_10')
// (2, 13, 'sp4_v_t_43')
// (2, 14, 'local_g3_3')
// (2, 14, 'lutff_7/in_3')
// (2, 14, 'sp4_v_b_43')
// (2, 15, 'sp4_v_b_30')
// (2, 16, 'local_g1_3')
// (2, 16, 'lutff_4/in_0')
// (2, 16, 'lutff_7/in_3')
// (2, 16, 'sp4_v_b_19')
// (2, 17, 'sp4_v_b_6')
// (3, 10, 'neigh_op_tnl_1')
// (3, 11, 'neigh_op_lft_1')
// (3, 12, 'neigh_op_bnl_1')
// (3, 13, 'sp4_h_r_17')
// (4, 13, 'sp4_h_r_28')
// (5, 13, 'sp4_h_r_41')
// (5, 14, 'sp4_r_v_b_41')
// (5, 15, 'sp4_r_v_b_28')
// (5, 16, 'local_g3_1')
// (5, 16, 'lutff_4/in_2')
// (5, 16, 'lutff_6/in_0')
// (5, 16, 'lutff_7/in_3')
// (5, 16, 'sp4_r_v_b_17')
// (5, 17, 'local_g1_4')
// (5, 17, 'lutff_0/in_1')
// (5, 17, 'lutff_4/in_3')
// (5, 17, 'sp4_r_v_b_4')
// (6, 13, 'sp4_h_l_41')
// (6, 13, 'sp4_v_t_41')
// (6, 14, 'sp4_v_b_41')
// (6, 15, 'sp4_v_b_28')
// (6, 16, 'sp4_v_b_17')
// (6, 17, 'sp4_v_b_4')

wire n253;
// (1, 10, 'neigh_op_tnr_2')
// (1, 11, 'neigh_op_rgt_2')
// (1, 12, 'local_g0_2')
// (1, 12, 'lutff_3/in_1')
// (1, 12, 'neigh_op_bnr_2')
// (2, 10, 'local_g1_2')
// (2, 10, 'lutff_3/in_2')
// (2, 10, 'lutff_4/in_3')
// (2, 10, 'neigh_op_top_2')
// (2, 11, 'lutff_2/out')
// (2, 12, 'neigh_op_bot_2')
// (3, 10, 'neigh_op_tnl_2')
// (3, 11, 'neigh_op_lft_2')
// (3, 12, 'neigh_op_bnl_2')

wire n254;
// (1, 10, 'neigh_op_tnr_3')
// (1, 11, 'neigh_op_rgt_3')
// (1, 12, 'neigh_op_bnr_3')
// (2, 10, 'local_g1_3')
// (2, 10, 'lutff_6/in_0')
// (2, 10, 'neigh_op_top_3')
// (2, 11, 'lutff_3/out')
// (2, 12, 'neigh_op_bot_3')
// (3, 10, 'neigh_op_tnl_3')
// (3, 11, 'neigh_op_lft_3')
// (3, 12, 'neigh_op_bnl_3')

wire n255;
// (1, 10, 'neigh_op_tnr_5')
// (1, 11, 'neigh_op_rgt_5')
// (1, 12, 'neigh_op_bnr_5')
// (2, 10, 'neigh_op_top_5')
// (2, 11, 'lutff_5/out')
// (2, 12, 'local_g1_5')
// (2, 12, 'lutff_1/in_3')
// (2, 12, 'neigh_op_bot_5')
// (3, 10, 'neigh_op_tnl_5')
// (3, 11, 'neigh_op_lft_5')
// (3, 12, 'neigh_op_bnl_5')

wire n256;
// (1, 10, 'neigh_op_tnr_6')
// (1, 11, 'neigh_op_rgt_6')
// (1, 12, 'neigh_op_bnr_6')
// (2, 10, 'neigh_op_top_6')
// (2, 11, 'lutff_6/out')
// (2, 12, 'local_g1_6')
// (2, 12, 'lutff_1/in_2')
// (2, 12, 'lutff_3/in_0')
// (2, 12, 'neigh_op_bot_6')
// (3, 10, 'neigh_op_tnl_6')
// (3, 11, 'neigh_op_lft_6')
// (3, 12, 'neigh_op_bnl_6')

wire n257;
// (1, 10, 'sp4_r_v_b_43')
// (1, 11, 'sp4_r_v_b_30')
// (1, 12, 'sp4_r_v_b_19')
// (1, 13, 'sp4_r_v_b_6')
// (1, 14, 'sp4_r_v_b_47')
// (1, 15, 'sp4_r_v_b_34')
// (1, 16, 'neigh_op_tnr_5')
// (1, 16, 'sp4_r_v_b_23')
// (1, 17, 'local_g2_5')
// (1, 17, 'lutff_6/in_1')
// (1, 17, 'neigh_op_rgt_5')
// (1, 17, 'sp4_r_v_b_10')
// (1, 18, 'neigh_op_bnr_5')
// (2, 9, 'sp4_v_t_43')
// (2, 10, 'sp4_r_v_b_42')
// (2, 10, 'sp4_v_b_43')
// (2, 11, 'sp4_r_v_b_31')
// (2, 11, 'sp4_v_b_30')
// (2, 12, 'local_g1_3')
// (2, 12, 'lutff_3/in_1')
// (2, 12, 'sp4_r_v_b_18')
// (2, 12, 'sp4_v_b_19')
// (2, 13, 'sp4_r_v_b_7')
// (2, 13, 'sp4_v_b_6')
// (2, 13, 'sp4_v_t_47')
// (2, 14, 'sp4_r_v_b_46')
// (2, 14, 'sp4_v_b_47')
// (2, 15, 'local_g2_2')
// (2, 15, 'lutff_1/in_3')
// (2, 15, 'lutff_4/in_0')
// (2, 15, 'sp4_r_v_b_35')
// (2, 15, 'sp4_v_b_34')
// (2, 16, 'neigh_op_top_5')
// (2, 16, 'sp4_r_v_b_22')
// (2, 16, 'sp4_v_b_23')
// (2, 17, 'local_g2_5')
// (2, 17, 'lutff_4/in_3')
// (2, 17, 'lutff_5/out')
// (2, 17, 'sp4_r_v_b_11')
// (2, 17, 'sp4_v_b_10')
// (2, 18, 'neigh_op_bot_5')
// (3, 9, 'sp4_v_t_42')
// (3, 10, 'sp4_v_b_42')
// (3, 11, 'sp4_v_b_31')
// (3, 12, 'local_g0_2')
// (3, 12, 'lutff_6/in_0')
// (3, 12, 'sp4_v_b_18')
// (3, 13, 'sp4_v_b_7')
// (3, 13, 'sp4_v_t_46')
// (3, 14, 'sp4_v_b_46')
// (3, 15, 'sp4_v_b_35')
// (3, 16, 'neigh_op_tnl_5')
// (3, 16, 'sp4_v_b_22')
// (3, 17, 'local_g0_5')
// (3, 17, 'lutff_5/in_0')
// (3, 17, 'lutff_7/in_2')
// (3, 17, 'neigh_op_lft_5')
// (3, 17, 'sp4_v_b_11')
// (3, 18, 'neigh_op_bnl_5')

wire n258;
// (1, 10, 'sp4_r_v_b_45')
// (1, 11, 'local_g0_3')
// (1, 11, 'lutff_2/in_1')
// (1, 11, 'sp4_r_v_b_32')
// (1, 12, 'sp4_r_v_b_21')
// (1, 13, 'sp4_r_v_b_8')
// (1, 14, 'sp4_r_v_b_37')
// (1, 15, 'sp4_r_v_b_24')
// (1, 16, 'sp4_r_v_b_13')
// (1, 17, 'sp4_r_v_b_0')
// (2, 9, 'sp4_v_t_45')
// (2, 10, 'local_g2_5')
// (2, 10, 'lutff_7/in_2')
// (2, 10, 'sp4_v_b_45')
// (2, 11, 'sp4_v_b_32')
// (2, 12, 'sp4_v_b_21')
// (2, 13, 'sp4_v_b_8')
// (2, 13, 'sp4_v_t_37')
// (2, 14, 'sp4_v_b_37')
// (2, 15, 'local_g2_0')
// (2, 15, 'lutff_4/in_2')
// (2, 15, 'sp4_v_b_24')
// (2, 16, 'local_g0_5')
// (2, 16, 'lutff_6/in_3')
// (2, 16, 'sp4_v_b_13')
// (2, 17, 'sp4_h_r_0')
// (2, 17, 'sp4_v_b_0')
// (3, 10, 'sp4_r_v_b_41')
// (3, 11, 'sp4_r_v_b_28')
// (3, 12, 'local_g3_1')
// (3, 12, 'lutff_1/in_3')
// (3, 12, 'sp4_r_v_b_17')
// (3, 13, 'sp4_r_v_b_4')
// (3, 14, 'sp4_r_v_b_45')
// (3, 15, 'sp4_r_v_b_32')
// (3, 16, 'neigh_op_tnr_4')
// (3, 16, 'sp4_r_v_b_21')
// (3, 17, 'neigh_op_rgt_4')
// (3, 17, 'sp4_h_r_13')
// (3, 17, 'sp4_r_v_b_8')
// (3, 18, 'neigh_op_bnr_4')
// (4, 9, 'sp4_v_t_41')
// (4, 10, 'sp4_v_b_41')
// (4, 11, 'sp4_v_b_28')
// (4, 12, 'sp4_v_b_17')
// (4, 13, 'sp4_v_b_4')
// (4, 13, 'sp4_v_t_45')
// (4, 14, 'sp4_r_v_b_44')
// (4, 14, 'sp4_v_b_45')
// (4, 15, 'sp4_r_v_b_33')
// (4, 15, 'sp4_v_b_32')
// (4, 16, 'neigh_op_top_4')
// (4, 16, 'sp4_r_v_b_20')
// (4, 16, 'sp4_r_v_b_36')
// (4, 16, 'sp4_v_b_21')
// (4, 17, 'lutff_4/out')
// (4, 17, 'sp4_h_r_24')
// (4, 17, 'sp4_r_v_b_25')
// (4, 17, 'sp4_r_v_b_9')
// (4, 17, 'sp4_v_b_8')
// (4, 18, 'neigh_op_bot_4')
// (4, 18, 'sp4_r_v_b_12')
// (4, 19, 'sp4_r_v_b_1')
// (5, 13, 'sp4_h_r_9')
// (5, 13, 'sp4_v_t_44')
// (5, 14, 'sp4_v_b_44')
// (5, 15, 'sp4_h_r_1')
// (5, 15, 'sp4_v_b_33')
// (5, 15, 'sp4_v_t_36')
// (5, 16, 'neigh_op_tnl_4')
// (5, 16, 'sp4_v_b_20')
// (5, 16, 'sp4_v_b_36')
// (5, 17, 'neigh_op_lft_4')
// (5, 17, 'sp4_h_r_37')
// (5, 17, 'sp4_v_b_25')
// (5, 17, 'sp4_v_b_9')
// (5, 18, 'neigh_op_bnl_4')
// (5, 18, 'sp4_v_b_12')
// (5, 19, 'sp4_v_b_1')
// (6, 13, 'sp4_h_r_20')
// (6, 15, 'sp4_h_r_12')
// (6, 17, 'sp4_h_l_37')
// (7, 13, 'sp4_h_r_33')
// (7, 15, 'sp4_h_r_25')
// (8, 10, 'sp4_r_v_b_44')
// (8, 11, 'sp4_r_v_b_33')
// (8, 12, 'sp4_r_v_b_20')
// (8, 13, 'sp4_h_r_44')
// (8, 13, 'sp4_r_v_b_9')
// (8, 15, 'sp4_h_r_36')
// (9, 9, 'sp4_v_t_44')
// (9, 10, 'sp4_v_b_44')
// (9, 11, 'local_g2_1')
// (9, 11, 'lutff_6/in_1')
// (9, 11, 'sp4_v_b_33')
// (9, 12, 'sp4_v_b_20')
// (9, 13, 'sp4_h_l_44')
// (9, 13, 'sp4_v_b_9')
// (9, 15, 'sp4_h_l_36')
// (9, 15, 'sp4_h_r_9')
// (10, 15, 'sp4_h_r_20')
// (11, 15, 'local_g2_1')
// (11, 15, 'lutff_4/in_3')
// (11, 15, 'sp4_h_r_33')
// (12, 15, 'sp4_h_r_44')
// (13, 15, 'sp4_h_l_44')

wire n259;
// (1, 10, 'sp4_r_v_b_46')
// (1, 11, 'sp4_r_v_b_35')
// (1, 12, 'sp4_r_v_b_22')
// (1, 13, 'sp4_r_v_b_11')
// (2, 9, 'sp4_v_t_46')
// (2, 10, 'sp4_v_b_46')
// (2, 11, 'local_g2_3')
// (2, 11, 'lutff_6/in_1')
// (2, 11, 'sp4_v_b_35')
// (2, 12, 'sp4_v_b_22')
// (2, 13, 'sp4_h_r_6')
// (2, 13, 'sp4_v_b_11')
// (3, 12, 'local_g2_7')
// (3, 12, 'lutff_6/in_3')
// (3, 12, 'neigh_op_tnr_7')
// (3, 13, 'neigh_op_rgt_7')
// (3, 13, 'sp4_h_r_19')
// (3, 14, 'neigh_op_bnr_7')
// (4, 12, 'neigh_op_top_7')
// (4, 13, 'lutff_7/out')
// (4, 13, 'sp4_h_r_30')
// (4, 14, 'neigh_op_bot_7')
// (5, 12, 'neigh_op_tnl_7')
// (5, 13, 'neigh_op_lft_7')
// (5, 13, 'sp4_h_r_43')
// (5, 14, 'neigh_op_bnl_7')
// (6, 13, 'sp4_h_l_43')

wire n260;
// (1, 11, 'local_g2_2')
// (1, 11, 'lutff_3/in_1')
// (1, 11, 'neigh_op_tnr_2')
// (1, 12, 'local_g3_2')
// (1, 12, 'lutff_4/in_3')
// (1, 12, 'neigh_op_rgt_2')
// (1, 13, 'neigh_op_bnr_2')
// (2, 11, 'local_g1_2')
// (2, 11, 'lutff_1/in_0')
// (2, 11, 'lutff_6/in_3')
// (2, 11, 'neigh_op_top_2')
// (2, 12, 'lutff_2/out')
// (2, 13, 'neigh_op_bot_2')
// (3, 11, 'local_g3_2')
// (3, 11, 'lutff_7/in_2')
// (3, 11, 'neigh_op_tnl_2')
// (3, 12, 'neigh_op_lft_2')
// (3, 13, 'neigh_op_bnl_2')

reg n261 = 0;
// (1, 11, 'neigh_op_tnr_1')
// (1, 12, 'local_g2_1')
// (1, 12, 'local_g3_1')
// (1, 12, 'lutff_2/in_3')
// (1, 12, 'lutff_4/in_0')
// (1, 12, 'neigh_op_rgt_1')
// (1, 13, 'neigh_op_bnr_1')
// (2, 9, 'sp12_v_t_22')
// (2, 10, 'sp12_v_b_22')
// (2, 11, 'neigh_op_top_1')
// (2, 11, 'sp12_v_b_21')
// (2, 12, 'local_g1_1')
// (2, 12, 'lutff_1/in_1')
// (2, 12, 'lutff_1/out')
// (2, 12, 'sp12_v_b_18')
// (2, 12, 'sp4_h_r_2')
// (2, 13, 'neigh_op_bot_1')
// (2, 13, 'sp12_v_b_17')
// (2, 14, 'sp12_v_b_14')
// (2, 15, 'sp12_v_b_13')
// (2, 16, 'sp12_v_b_10')
// (2, 17, 'sp12_v_b_9')
// (2, 18, 'sp12_v_b_6')
// (2, 19, 'sp12_v_b_5')
// (2, 20, 'sp12_v_b_2')
// (2, 21, 'sp12_h_r_1')
// (2, 21, 'sp12_v_b_1')
// (3, 11, 'neigh_op_tnl_1')
// (3, 12, 'neigh_op_lft_1')
// (3, 12, 'sp4_h_r_15')
// (3, 13, 'neigh_op_bnl_1')
// (3, 21, 'sp12_h_r_2')
// (4, 12, 'sp4_h_r_26')
// (4, 21, 'sp12_h_r_5')
// (5, 12, 'local_g2_7')
// (5, 12, 'lutff_2/in_1')
// (5, 12, 'sp4_h_r_39')
// (5, 13, 'sp4_r_v_b_39')
// (5, 14, 'sp4_r_v_b_26')
// (5, 15, 'local_g2_7')
// (5, 15, 'lutff_0/in_1')
// (5, 15, 'sp4_r_v_b_15')
// (5, 16, 'sp4_r_v_b_2')
// (5, 21, 'sp12_h_r_6')
// (6, 12, 'sp4_h_l_39')
// (6, 12, 'sp4_h_r_5')
// (6, 12, 'sp4_v_t_39')
// (6, 13, 'sp4_v_b_39')
// (6, 14, 'sp4_v_b_26')
// (6, 15, 'sp4_v_b_15')
// (6, 16, 'sp4_v_b_2')
// (6, 21, 'sp12_h_r_9')
// (7, 12, 'sp4_h_r_16')
// (7, 21, 'sp12_h_r_10')
// (8, 12, 'sp4_h_r_29')
// (8, 21, 'sp12_h_r_13')
// (9, 9, 'sp4_r_v_b_46')
// (9, 10, 'sp4_r_v_b_35')
// (9, 11, 'sp4_r_v_b_22')
// (9, 12, 'sp4_h_r_40')
// (9, 12, 'sp4_r_v_b_11')
// (9, 21, 'sp12_h_r_14')
// (10, 8, 'sp4_v_t_46')
// (10, 9, 'sp4_v_b_46')
// (10, 10, 'sp4_v_b_35')
// (10, 11, 'local_g0_6')
// (10, 11, 'lutff_5/in_1')
// (10, 11, 'sp4_v_b_22')
// (10, 12, 'sp4_h_l_40')
// (10, 12, 'sp4_v_b_11')
// (10, 21, 'sp12_h_r_17')
// (11, 21, 'local_g0_2')
// (11, 21, 'lutff_6/in_2')
// (11, 21, 'sp12_h_r_18')
// (12, 21, 'sp12_h_r_21')
// (13, 21, 'sp12_h_r_22')
// (14, 21, 'sp12_h_l_22')

wire n262;
// (1, 11, 'neigh_op_tnr_4')
// (1, 12, 'neigh_op_rgt_4')
// (1, 13, 'neigh_op_bnr_4')
// (2, 11, 'neigh_op_top_4')
// (2, 12, 'local_g3_4')
// (2, 12, 'lutff_4/out')
// (2, 12, 'lutff_5/in_0')
// (2, 13, 'neigh_op_bot_4')
// (3, 11, 'neigh_op_tnl_4')
// (3, 12, 'neigh_op_lft_4')
// (3, 13, 'neigh_op_bnl_4')

wire n263;
// (1, 11, 'neigh_op_tnr_7')
// (1, 12, 'neigh_op_rgt_7')
// (1, 13, 'local_g0_7')
// (1, 13, 'lutff_7/in_0')
// (1, 13, 'neigh_op_bnr_7')
// (2, 11, 'neigh_op_top_7')
// (2, 12, 'lutff_7/out')
// (2, 13, 'neigh_op_bot_7')
// (3, 11, 'neigh_op_tnl_7')
// (3, 12, 'neigh_op_lft_7')
// (3, 13, 'neigh_op_bnl_7')

reg n264 = 0;
// (1, 11, 'sp4_h_r_1')
// (1, 12, 'sp4_h_r_1')
// (1, 18, 'sp4_h_r_1')
// (2, 11, 'local_g0_4')
// (2, 11, 'lutff_5/in_3')
// (2, 11, 'sp4_h_r_12')
// (2, 12, 'local_g0_4')
// (2, 12, 'lutff_7/in_3')
// (2, 12, 'sp4_h_r_12')
// (2, 12, 'sp4_r_v_b_44')
// (2, 13, 'sp4_r_v_b_33')
// (2, 14, 'sp4_r_v_b_20')
// (2, 15, 'local_g2_1')
// (2, 15, 'lutff_7/in_0')
// (2, 15, 'sp4_r_v_b_9')
// (2, 18, 'local_g0_4')
// (2, 18, 'lutff_7/in_3')
// (2, 18, 'sp4_h_r_12')
// (3, 9, 'sp4_r_v_b_44')
// (3, 10, 'neigh_op_tnr_2')
// (3, 10, 'sp4_r_v_b_33')
// (3, 11, 'local_g1_1')
// (3, 11, 'lutff_7/in_3')
// (3, 11, 'neigh_op_rgt_2')
// (3, 11, 'sp4_h_r_25')
// (3, 11, 'sp4_h_r_9')
// (3, 11, 'sp4_r_v_b_20')
// (3, 11, 'sp4_v_t_44')
// (3, 12, 'neigh_op_bnr_2')
// (3, 12, 'sp4_h_r_25')
// (3, 12, 'sp4_r_v_b_9')
// (3, 12, 'sp4_v_b_44')
// (3, 13, 'sp4_r_v_b_40')
// (3, 13, 'sp4_v_b_33')
// (3, 14, 'sp4_r_v_b_29')
// (3, 14, 'sp4_v_b_20')
// (3, 15, 'sp4_r_v_b_16')
// (3, 15, 'sp4_v_b_9')
// (3, 16, 'sp4_r_v_b_5')
// (3, 18, 'sp4_h_r_25')
// (4, 8, 'sp4_v_t_44')
// (4, 9, 'sp4_r_v_b_45')
// (4, 9, 'sp4_v_b_44')
// (4, 10, 'neigh_op_top_2')
// (4, 10, 'sp4_r_v_b_32')
// (4, 10, 'sp4_v_b_33')
// (4, 11, 'lutff_2/out')
// (4, 11, 'sp4_h_r_20')
// (4, 11, 'sp4_h_r_36')
// (4, 11, 'sp4_h_r_4')
// (4, 11, 'sp4_r_v_b_21')
// (4, 11, 'sp4_r_v_b_37')
// (4, 11, 'sp4_v_b_20')
// (4, 12, 'neigh_op_bot_2')
// (4, 12, 'sp4_h_r_36')
// (4, 12, 'sp4_r_v_b_24')
// (4, 12, 'sp4_r_v_b_8')
// (4, 12, 'sp4_v_b_9')
// (4, 12, 'sp4_v_t_40')
// (4, 13, 'sp4_r_v_b_13')
// (4, 13, 'sp4_r_v_b_46')
// (4, 13, 'sp4_v_b_40')
// (4, 14, 'sp4_r_v_b_0')
// (4, 14, 'sp4_r_v_b_35')
// (4, 14, 'sp4_v_b_29')
// (4, 15, 'sp4_r_v_b_22')
// (4, 15, 'sp4_r_v_b_45')
// (4, 15, 'sp4_v_b_16')
// (4, 16, 'local_g0_5')
// (4, 16, 'lutff_4/in_1')
// (4, 16, 'sp4_r_v_b_11')
// (4, 16, 'sp4_r_v_b_32')
// (4, 16, 'sp4_v_b_5')
// (4, 17, 'sp4_r_v_b_21')
// (4, 18, 'sp4_h_r_36')
// (4, 18, 'sp4_r_v_b_8')
// (5, 8, 'sp4_v_t_45')
// (5, 9, 'sp4_v_b_45')
// (5, 10, 'neigh_op_tnl_2')
// (5, 10, 'sp4_v_b_32')
// (5, 10, 'sp4_v_t_37')
// (5, 11, 'neigh_op_lft_2')
// (5, 11, 'sp4_h_l_36')
// (5, 11, 'sp4_h_r_17')
// (5, 11, 'sp4_h_r_33')
// (5, 11, 'sp4_v_b_21')
// (5, 11, 'sp4_v_b_37')
// (5, 12, 'neigh_op_bnl_2')
// (5, 12, 'sp4_h_l_36')
// (5, 12, 'sp4_v_b_24')
// (5, 12, 'sp4_v_b_8')
// (5, 12, 'sp4_v_t_46')
// (5, 13, 'sp4_v_b_13')
// (5, 13, 'sp4_v_b_46')
// (5, 14, 'sp4_v_b_0')
// (5, 14, 'sp4_v_b_35')
// (5, 14, 'sp4_v_t_45')
// (5, 15, 'local_g1_6')
// (5, 15, 'lutff_3/in_0')
// (5, 15, 'sp4_v_b_22')
// (5, 15, 'sp4_v_b_45')
// (5, 16, 'sp4_h_r_5')
// (5, 16, 'sp4_v_b_11')
// (5, 16, 'sp4_v_b_32')
// (5, 17, 'sp4_v_b_21')
// (5, 18, 'sp4_h_l_36')
// (5, 18, 'sp4_v_b_8')
// (6, 11, 'sp4_h_r_28')
// (6, 11, 'sp4_h_r_44')
// (6, 16, 'sp4_h_r_16')
// (7, 11, 'sp4_h_l_44')
// (7, 11, 'sp4_h_r_41')
// (7, 12, 'sp4_r_v_b_41')
// (7, 13, 'sp4_r_v_b_28')
// (7, 14, 'sp4_r_v_b_17')
// (7, 15, 'sp4_r_v_b_4')
// (7, 16, 'sp4_h_r_29')
// (8, 11, 'sp4_h_l_41')
// (8, 11, 'sp4_h_r_4')
// (8, 11, 'sp4_v_t_41')
// (8, 12, 'sp4_v_b_41')
// (8, 13, 'sp4_v_b_28')
// (8, 14, 'sp4_v_b_17')
// (8, 15, 'sp4_h_r_10')
// (8, 15, 'sp4_v_b_4')
// (8, 16, 'sp4_h_r_40')
// (9, 11, 'sp4_h_r_17')
// (9, 15, 'sp4_h_r_23')
// (9, 16, 'sp4_h_l_40')
// (9, 16, 'sp4_h_r_5')
// (10, 11, 'sp4_h_r_28')
// (10, 15, 'sp4_h_r_34')
// (10, 16, 'sp4_h_r_16')
// (11, 11, 'sp4_h_r_41')
// (11, 12, 'sp4_r_v_b_44')
// (11, 13, 'sp4_r_v_b_33')
// (11, 14, 'sp4_r_v_b_20')
// (11, 15, 'local_g3_7')
// (11, 15, 'lutff_3/in_3')
// (11, 15, 'sp4_h_r_47')
// (11, 15, 'sp4_r_v_b_9')
// (11, 16, 'local_g3_5')
// (11, 16, 'lutff_5/in_3')
// (11, 16, 'sp4_h_r_29')
// (11, 16, 'sp4_r_v_b_44')
// (11, 17, 'sp4_r_v_b_33')
// (11, 18, 'local_g3_4')
// (11, 18, 'lutff_5/in_0')
// (11, 18, 'sp4_r_v_b_20')
// (11, 19, 'sp4_r_v_b_9')
// (12, 11, 'sp4_h_l_41')
// (12, 11, 'sp4_v_t_44')
// (12, 12, 'sp4_v_b_44')
// (12, 13, 'sp4_v_b_33')
// (12, 14, 'sp4_v_b_20')
// (12, 15, 'sp4_h_l_47')
// (12, 15, 'sp4_v_b_9')
// (12, 15, 'sp4_v_t_44')
// (12, 16, 'sp4_h_r_40')
// (12, 16, 'sp4_v_b_44')
// (12, 17, 'sp4_v_b_33')
// (12, 18, 'sp4_v_b_20')
// (12, 19, 'sp4_v_b_9')
// (13, 16, 'sp4_h_l_40')

wire n265;
// (1, 11, 'sp4_h_r_11')
// (2, 11, 'sp4_h_r_22')
// (3, 10, 'neigh_op_tnr_7')
// (3, 11, 'neigh_op_rgt_7')
// (3, 11, 'sp4_h_r_35')
// (3, 12, 'neigh_op_bnr_7')
// (4, 10, 'neigh_op_top_7')
// (4, 11, 'lutff_7/out')
// (4, 11, 'sp4_h_r_46')
// (4, 12, 'neigh_op_bot_7')
// (4, 12, 'sp4_r_v_b_46')
// (4, 13, 'sp4_r_v_b_35')
// (4, 14, 'sp4_r_v_b_22')
// (4, 15, 'local_g2_3')
// (4, 15, 'lutff_1/in_2')
// (4, 15, 'sp4_r_v_b_11')
// (5, 10, 'neigh_op_tnl_7')
// (5, 11, 'neigh_op_lft_7')
// (5, 11, 'sp4_h_l_46')
// (5, 11, 'sp4_v_t_46')
// (5, 12, 'neigh_op_bnl_7')
// (5, 12, 'sp4_v_b_46')
// (5, 13, 'sp4_v_b_35')
// (5, 14, 'sp4_v_b_22')
// (5, 15, 'sp4_v_b_11')

reg n266 = 0;
// (1, 11, 'sp4_r_v_b_36')
// (1, 12, 'sp4_r_v_b_25')
// (1, 13, 'local_g2_4')
// (1, 13, 'lutff_4/in_0')
// (1, 13, 'sp4_r_v_b_12')
// (1, 14, 'sp4_r_v_b_1')
// (1, 15, 'sp4_h_r_9')
// (2, 10, 'sp4_v_t_36')
// (2, 11, 'sp4_v_b_36')
// (2, 12, 'sp4_v_b_25')
// (2, 13, 'sp4_v_b_12')
// (2, 14, 'sp4_h_r_1')
// (2, 14, 'sp4_v_b_1')
// (2, 15, 'local_g0_4')
// (2, 15, 'lutff_0/in_2')
// (2, 15, 'sp4_h_r_20')
// (3, 14, 'sp4_h_r_12')
// (3, 15, 'sp4_h_r_33')
// (4, 11, 'sp4_r_v_b_41')
// (4, 12, 'sp4_r_v_b_28')
// (4, 12, 'sp4_r_v_b_44')
// (4, 13, 'local_g2_2')
// (4, 13, 'lutff_5/in_1')
// (4, 13, 'neigh_op_tnr_2')
// (4, 13, 'sp4_r_v_b_17')
// (4, 13, 'sp4_r_v_b_33')
// (4, 14, 'neigh_op_rgt_2')
// (4, 14, 'sp4_h_r_25')
// (4, 14, 'sp4_r_v_b_20')
// (4, 14, 'sp4_r_v_b_36')
// (4, 14, 'sp4_r_v_b_4')
// (4, 15, 'neigh_op_bnr_2')
// (4, 15, 'sp4_h_r_44')
// (4, 15, 'sp4_r_v_b_25')
// (4, 15, 'sp4_r_v_b_9')
// (4, 16, 'local_g2_4')
// (4, 16, 'lutff_4/in_0')
// (4, 16, 'sp4_r_v_b_12')
// (4, 17, 'sp4_r_v_b_1')
// (5, 10, 'sp4_v_t_41')
// (5, 11, 'sp4_v_b_41')
// (5, 11, 'sp4_v_t_44')
// (5, 12, 'local_g2_4')
// (5, 12, 'lutff_6/in_0')
// (5, 12, 'sp4_v_b_28')
// (5, 12, 'sp4_v_b_44')
// (5, 13, 'local_g1_2')
// (5, 13, 'lutff_6/in_3')
// (5, 13, 'neigh_op_top_2')
// (5, 13, 'sp4_v_b_17')
// (5, 13, 'sp4_v_b_33')
// (5, 13, 'sp4_v_t_36')
// (5, 14, 'local_g3_2')
// (5, 14, 'lutff_2/in_1')
// (5, 14, 'lutff_2/out')
// (5, 14, 'sp4_h_r_36')
// (5, 14, 'sp4_v_b_20')
// (5, 14, 'sp4_v_b_36')
// (5, 14, 'sp4_v_b_4')
// (5, 15, 'neigh_op_bot_2')
// (5, 15, 'sp4_h_l_44')
// (5, 15, 'sp4_v_b_25')
// (5, 15, 'sp4_v_b_9')
// (5, 16, 'local_g0_4')
// (5, 16, 'lutff_5/in_1')
// (5, 16, 'sp4_v_b_12')
// (5, 17, 'sp4_v_b_1')
// (6, 13, 'neigh_op_tnl_2')
// (6, 14, 'neigh_op_lft_2')
// (6, 14, 'sp4_h_l_36')
// (6, 15, 'neigh_op_bnl_2')

wire n267;
// (1, 11, 'sp4_r_v_b_37')
// (1, 12, 'local_g0_0')
// (1, 12, 'lutff_7/in_1')
// (1, 12, 'sp4_r_v_b_24')
// (1, 13, 'neigh_op_tnr_0')
// (1, 13, 'sp4_r_v_b_13')
// (1, 14, 'neigh_op_rgt_0')
// (1, 14, 'sp4_r_v_b_0')
// (1, 15, 'neigh_op_bnr_0')
// (2, 10, 'sp12_v_t_23')
// (2, 10, 'sp4_v_t_37')
// (2, 11, 'sp12_v_b_23')
// (2, 11, 'sp4_v_b_37')
// (2, 12, 'sp12_v_b_20')
// (2, 12, 'sp4_v_b_24')
// (2, 13, 'neigh_op_top_0')
// (2, 13, 'sp12_v_b_19')
// (2, 13, 'sp4_r_v_b_44')
// (2, 13, 'sp4_v_b_13')
// (2, 14, 'local_g3_0')
// (2, 14, 'lutff_0/out')
// (2, 14, 'lutff_3/in_2')
// (2, 14, 'sp12_v_b_16')
// (2, 14, 'sp4_r_v_b_33')
// (2, 14, 'sp4_v_b_0')
// (2, 15, 'neigh_op_bot_0')
// (2, 15, 'sp12_v_b_15')
// (2, 15, 'sp4_r_v_b_20')
// (2, 16, 'sp12_v_b_12')
// (2, 16, 'sp4_r_v_b_9')
// (2, 17, 'local_g3_3')
// (2, 17, 'lutff_3/in_1')
// (2, 17, 'sp12_v_b_11')
// (2, 18, 'sp12_v_b_8')
// (2, 19, 'sp12_v_b_7')
// (2, 20, 'sp12_v_b_4')
// (2, 21, 'local_g2_3')
// (2, 21, 'lutff_6/in_1')
// (2, 21, 'sp12_v_b_3')
// (2, 22, 'sp12_v_b_0')
// (3, 12, 'sp4_v_t_44')
// (3, 13, 'neigh_op_tnl_0')
// (3, 13, 'sp4_v_b_44')
// (3, 14, 'neigh_op_lft_0')
// (3, 14, 'sp4_v_b_33')
// (3, 15, 'neigh_op_bnl_0')
// (3, 15, 'sp4_v_b_20')
// (3, 16, 'sp4_h_r_9')
// (3, 16, 'sp4_v_b_9')
// (4, 16, 'sp4_h_r_20')
// (5, 16, 'local_g2_1')
// (5, 16, 'lutff_0/in_3')
// (5, 16, 'sp4_h_r_33')
// (6, 16, 'sp4_h_r_44')
// (7, 16, 'sp4_h_l_44')

wire n268;
// (1, 11, 'sp4_r_v_b_38')
// (1, 12, 'neigh_op_tnr_7')
// (1, 12, 'sp4_r_v_b_27')
// (1, 13, 'neigh_op_rgt_7')
// (1, 13, 'sp4_h_r_3')
// (1, 13, 'sp4_r_v_b_14')
// (1, 14, 'neigh_op_bnr_7')
// (1, 14, 'sp4_r_v_b_3')
// (1, 15, 'sp4_r_v_b_43')
// (1, 16, 'sp4_r_v_b_30')
// (1, 17, 'sp4_r_v_b_19')
// (1, 18, 'sp4_r_v_b_6')
// (2, 10, 'sp4_v_t_38')
// (2, 11, 'sp4_r_v_b_39')
// (2, 11, 'sp4_v_b_38')
// (2, 12, 'neigh_op_top_7')
// (2, 12, 'sp4_r_v_b_26')
// (2, 12, 'sp4_v_b_27')
// (2, 13, 'lutff_7/out')
// (2, 13, 'sp4_h_r_14')
// (2, 13, 'sp4_r_v_b_15')
// (2, 13, 'sp4_r_v_b_47')
// (2, 13, 'sp4_v_b_14')
// (2, 14, 'local_g0_7')
// (2, 14, 'lutff_6/in_3')
// (2, 14, 'neigh_op_bot_7')
// (2, 14, 'sp4_r_v_b_2')
// (2, 14, 'sp4_r_v_b_34')
// (2, 14, 'sp4_v_b_3')
// (2, 14, 'sp4_v_t_43')
// (2, 15, 'sp4_r_v_b_23')
// (2, 15, 'sp4_r_v_b_39')
// (2, 15, 'sp4_v_b_43')
// (2, 16, 'sp4_r_v_b_10')
// (2, 16, 'sp4_r_v_b_26')
// (2, 16, 'sp4_v_b_30')
// (2, 17, 'local_g1_3')
// (2, 17, 'lutff_5/in_1')
// (2, 17, 'sp4_r_v_b_15')
// (2, 17, 'sp4_v_b_19')
// (2, 18, 'local_g0_6')
// (2, 18, 'lutff_2/in_0')
// (2, 18, 'sp4_r_v_b_2')
// (2, 18, 'sp4_v_b_6')
// (3, 10, 'sp4_v_t_39')
// (3, 11, 'sp4_v_b_39')
// (3, 12, 'neigh_op_tnl_7')
// (3, 12, 'sp4_v_b_26')
// (3, 12, 'sp4_v_t_47')
// (3, 13, 'neigh_op_lft_7')
// (3, 13, 'sp4_h_r_27')
// (3, 13, 'sp4_v_b_15')
// (3, 13, 'sp4_v_b_47')
// (3, 14, 'neigh_op_bnl_7')
// (3, 14, 'sp4_v_b_2')
// (3, 14, 'sp4_v_b_34')
// (3, 14, 'sp4_v_t_39')
// (3, 15, 'sp4_v_b_23')
// (3, 15, 'sp4_v_b_39')
// (3, 16, 'sp4_h_r_10')
// (3, 16, 'sp4_v_b_10')
// (3, 16, 'sp4_v_b_26')
// (3, 17, 'sp4_v_b_15')
// (3, 18, 'local_g0_2')
// (3, 18, 'lutff_6/in_0')
// (3, 18, 'sp4_v_b_2')
// (4, 13, 'sp4_h_r_38')
// (4, 14, 'sp4_r_v_b_45')
// (4, 15, 'sp4_r_v_b_32')
// (4, 16, 'sp4_h_r_23')
// (4, 16, 'sp4_r_v_b_21')
// (4, 17, 'local_g2_0')
// (4, 17, 'lutff_3/in_1')
// (4, 17, 'sp4_r_v_b_8')
// (5, 13, 'sp4_h_l_38')
// (5, 13, 'sp4_v_t_45')
// (5, 14, 'sp4_v_b_45')
// (5, 15, 'sp4_v_b_32')
// (5, 16, 'local_g3_2')
// (5, 16, 'lutff_6/in_3')
// (5, 16, 'sp4_h_r_34')
// (5, 16, 'sp4_v_b_21')
// (5, 17, 'local_g1_0')
// (5, 17, 'lutff_3/in_0')
// (5, 17, 'sp4_v_b_8')
// (6, 16, 'sp4_h_r_47')
// (7, 16, 'sp4_h_l_47')

wire n269;
// (1, 11, 'sp4_r_v_b_45')
// (1, 12, 'sp4_r_v_b_32')
// (1, 13, 'neigh_op_tnr_4')
// (1, 13, 'sp4_r_v_b_21')
// (1, 14, 'neigh_op_rgt_4')
// (1, 14, 'sp4_r_v_b_8')
// (1, 15, 'neigh_op_bnr_4')
// (2, 10, 'sp4_v_t_45')
// (2, 11, 'sp4_v_b_45')
// (2, 12, 'sp4_v_b_32')
// (2, 13, 'neigh_op_top_4')
// (2, 13, 'sp4_v_b_21')
// (2, 14, 'local_g0_2')
// (2, 14, 'lutff_4/out')
// (2, 14, 'lutff_global/cen')
// (2, 14, 'sp4_h_r_2')
// (2, 14, 'sp4_v_b_8')
// (2, 15, 'neigh_op_bot_4')
// (3, 13, 'neigh_op_tnl_4')
// (3, 14, 'neigh_op_lft_4')
// (3, 14, 'sp4_h_r_15')
// (3, 15, 'neigh_op_bnl_4')
// (4, 14, 'sp4_h_r_26')
// (5, 14, 'sp4_h_r_39')
// (6, 14, 'sp4_h_l_39')

wire n270;
// (1, 12, 'local_g0_6')
// (1, 12, 'lutff_5/in_1')
// (1, 12, 'sp4_h_r_6')
// (2, 12, 'sp4_h_r_19')
// (3, 10, 'neigh_op_tnr_1')
// (3, 11, 'neigh_op_rgt_1')
// (3, 12, 'neigh_op_bnr_1')
// (3, 12, 'sp4_h_r_30')
// (4, 9, 'sp4_r_v_b_43')
// (4, 10, 'neigh_op_top_1')
// (4, 10, 'sp4_r_v_b_30')
// (4, 11, 'local_g2_1')
// (4, 11, 'lutff_1/out')
// (4, 11, 'lutff_6/in_3')
// (4, 11, 'sp4_r_v_b_19')
// (4, 12, 'neigh_op_bot_1')
// (4, 12, 'sp4_h_r_43')
// (4, 12, 'sp4_r_v_b_6')
// (5, 8, 'sp4_v_t_43')
// (5, 9, 'sp4_v_b_43')
// (5, 10, 'neigh_op_tnl_1')
// (5, 10, 'sp4_v_b_30')
// (5, 11, 'neigh_op_lft_1')
// (5, 11, 'sp4_v_b_19')
// (5, 12, 'neigh_op_bnl_1')
// (5, 12, 'sp4_h_l_43')
// (5, 12, 'sp4_v_b_6')

reg n271 = 0;
// (1, 12, 'local_g1_1')
// (1, 12, 'lutff_6/in_0')
// (1, 12, 'sp4_h_r_9')
// (1, 13, 'sp4_h_r_5')
// (1, 14, 'sp4_h_r_10')
// (2, 12, 'sp4_h_r_20')
// (2, 13, 'local_g1_0')
// (2, 13, 'lutff_5/in_0')
// (2, 13, 'sp4_h_r_16')
// (2, 14, 'local_g1_7')
// (2, 14, 'lutff_2/in_2')
// (2, 14, 'sp4_h_r_23')
// (3, 11, 'local_g3_6')
// (3, 11, 'lutff_6/in_3')
// (3, 11, 'neigh_op_tnr_6')
// (3, 11, 'sp4_r_v_b_41')
// (3, 12, 'neigh_op_rgt_6')
// (3, 12, 'sp4_h_r_33')
// (3, 12, 'sp4_r_v_b_28')
// (3, 13, 'neigh_op_bnr_6')
// (3, 13, 'sp4_h_r_29')
// (3, 13, 'sp4_r_v_b_17')
// (3, 14, 'local_g1_4')
// (3, 14, 'lutff_7/in_0')
// (3, 14, 'sp4_h_r_34')
// (3, 14, 'sp4_r_v_b_4')
// (4, 10, 'sp4_r_v_b_37')
// (4, 10, 'sp4_v_t_41')
// (4, 11, 'neigh_op_top_6')
// (4, 11, 'sp4_r_v_b_24')
// (4, 11, 'sp4_r_v_b_40')
// (4, 11, 'sp4_v_b_41')
// (4, 12, 'local_g1_6')
// (4, 12, 'lutff_0/in_1')
// (4, 12, 'lutff_6/in_3')
// (4, 12, 'lutff_6/out')
// (4, 12, 'sp4_h_r_44')
// (4, 12, 'sp4_r_v_b_13')
// (4, 12, 'sp4_r_v_b_29')
// (4, 12, 'sp4_r_v_b_45')
// (4, 12, 'sp4_v_b_28')
// (4, 13, 'neigh_op_bot_6')
// (4, 13, 'sp4_h_r_40')
// (4, 13, 'sp4_r_v_b_0')
// (4, 13, 'sp4_r_v_b_16')
// (4, 13, 'sp4_r_v_b_32')
// (4, 13, 'sp4_v_b_17')
// (4, 14, 'sp4_h_r_47')
// (4, 14, 'sp4_r_v_b_21')
// (4, 14, 'sp4_r_v_b_5')
// (4, 14, 'sp4_v_b_4')
// (4, 15, 'local_g2_0')
// (4, 15, 'lutff_7/in_3')
// (4, 15, 'sp4_r_v_b_8')
// (5, 9, 'sp4_v_t_37')
// (5, 10, 'sp4_v_b_37')
// (5, 10, 'sp4_v_t_40')
// (5, 11, 'neigh_op_tnl_6')
// (5, 11, 'sp4_v_b_24')
// (5, 11, 'sp4_v_b_40')
// (5, 11, 'sp4_v_t_45')
// (5, 12, 'local_g0_6')
// (5, 12, 'lutff_5/in_1')
// (5, 12, 'neigh_op_lft_6')
// (5, 12, 'sp4_h_l_44')
// (5, 12, 'sp4_v_b_13')
// (5, 12, 'sp4_v_b_29')
// (5, 12, 'sp4_v_b_45')
// (5, 13, 'local_g2_6')
// (5, 13, 'lutff_3/in_3')
// (5, 13, 'lutff_4/in_0')
// (5, 13, 'lutff_7/in_3')
// (5, 13, 'neigh_op_bnl_6')
// (5, 13, 'sp4_h_l_40')
// (5, 13, 'sp4_v_b_0')
// (5, 13, 'sp4_v_b_16')
// (5, 13, 'sp4_v_b_32')
// (5, 14, 'sp4_h_l_47')
// (5, 14, 'sp4_v_b_21')
// (5, 14, 'sp4_v_b_5')
// (5, 15, 'sp4_v_b_8')

wire n272;
// (1, 12, 'local_g3_4')
// (1, 12, 'lutff_0/in_3')
// (1, 12, 'neigh_op_tnr_4')
// (1, 13, 'neigh_op_rgt_4')
// (1, 14, 'neigh_op_bnr_4')
// (2, 6, 'sp4_r_v_b_44')
// (2, 7, 'local_g0_2')
// (2, 7, 'lutff_6/in_0')
// (2, 7, 'sp4_r_v_b_33')
// (2, 8, 'sp4_r_v_b_20')
// (2, 9, 'sp4_r_v_b_9')
// (2, 10, 'sp4_r_v_b_44')
// (2, 11, 'local_g2_1')
// (2, 11, 'lutff_5/in_2')
// (2, 11, 'sp4_r_v_b_33')
// (2, 12, 'local_g1_4')
// (2, 12, 'lutff_4/in_3')
// (2, 12, 'neigh_op_top_4')
// (2, 12, 'sp4_r_v_b_20')
// (2, 13, 'lutff_4/out')
// (2, 13, 'sp4_r_v_b_9')
// (2, 14, 'neigh_op_bot_4')
// (3, 5, 'sp4_v_t_44')
// (3, 6, 'sp4_v_b_44')
// (3, 7, 'sp4_v_b_33')
// (3, 8, 'sp4_v_b_20')
// (3, 9, 'sp4_v_b_9')
// (3, 9, 'sp4_v_t_44')
// (3, 10, 'sp4_v_b_44')
// (3, 11, 'sp4_v_b_33')
// (3, 12, 'neigh_op_tnl_4')
// (3, 12, 'sp4_v_b_20')
// (3, 13, 'neigh_op_lft_4')
// (3, 13, 'sp4_v_b_9')
// (3, 14, 'neigh_op_bnl_4')

wire n273;
// (1, 12, 'neigh_op_tnr_1')
// (1, 13, 'local_g3_1')
// (1, 13, 'lutff_6/in_2')
// (1, 13, 'lutff_7/in_1')
// (1, 13, 'neigh_op_rgt_1')
// (1, 14, 'neigh_op_bnr_1')
// (2, 12, 'neigh_op_top_1')
// (2, 13, 'lutff_1/out')
// (2, 14, 'neigh_op_bot_1')
// (3, 12, 'neigh_op_tnl_1')
// (3, 13, 'neigh_op_lft_1')
// (3, 14, 'neigh_op_bnl_1')

wire n274;
// (1, 12, 'neigh_op_tnr_2')
// (1, 13, 'neigh_op_rgt_2')
// (1, 13, 'sp4_h_r_9')
// (1, 13, 'sp4_r_v_b_36')
// (1, 14, 'neigh_op_bnr_2')
// (1, 14, 'sp4_r_v_b_25')
// (1, 15, 'sp4_r_v_b_12')
// (1, 16, 'sp4_r_v_b_1')
// (2, 12, 'neigh_op_top_2')
// (2, 12, 'sp4_h_r_1')
// (2, 12, 'sp4_v_t_36')
// (2, 13, 'local_g3_2')
// (2, 13, 'lutff_2/out')
// (2, 13, 'lutff_5/in_2')
// (2, 13, 'sp4_h_r_20')
// (2, 13, 'sp4_v_b_36')
// (2, 14, 'neigh_op_bot_2')
// (2, 14, 'sp4_v_b_25')
// (2, 15, 'sp4_v_b_12')
// (2, 16, 'sp4_v_b_1')
// (3, 12, 'local_g3_2')
// (3, 12, 'lutff_2/in_1')
// (3, 12, 'neigh_op_tnl_2')
// (3, 12, 'sp4_h_r_12')
// (3, 13, 'neigh_op_lft_2')
// (3, 13, 'sp4_h_r_33')
// (3, 14, 'neigh_op_bnl_2')
// (4, 10, 'sp4_r_v_b_44')
// (4, 11, 'sp4_r_v_b_33')
// (4, 12, 'local_g3_1')
// (4, 12, 'local_g3_4')
// (4, 12, 'lutff_2/in_0')
// (4, 12, 'lutff_3/in_0')
// (4, 12, 'lutff_4/in_0')
// (4, 12, 'lutff_5/in_0')
// (4, 12, 'lutff_6/in_1')
// (4, 12, 'sp4_h_r_25')
// (4, 12, 'sp4_r_v_b_20')
// (4, 13, 'sp4_h_r_44')
// (4, 13, 'sp4_r_v_b_9')
// (5, 9, 'sp4_v_t_44')
// (5, 10, 'sp4_v_b_44')
// (5, 11, 'sp4_v_b_33')
// (5, 12, 'sp4_h_r_36')
// (5, 12, 'sp4_v_b_20')
// (5, 13, 'sp4_h_l_44')
// (5, 13, 'sp4_v_b_9')
// (6, 12, 'sp4_h_l_36')

wire n275;
// (1, 12, 'neigh_op_tnr_6')
// (1, 13, 'neigh_op_rgt_6')
// (1, 14, 'neigh_op_bnr_6')
// (2, 12, 'neigh_op_top_6')
// (2, 12, 'sp4_r_v_b_40')
// (2, 13, 'lutff_6/out')
// (2, 13, 'sp4_r_v_b_29')
// (2, 14, 'neigh_op_bot_6')
// (2, 14, 'sp4_r_v_b_16')
// (2, 15, 'sp4_r_v_b_5')
// (3, 11, 'sp4_v_t_40')
// (3, 12, 'neigh_op_tnl_6')
// (3, 12, 'sp4_v_b_40')
// (3, 13, 'neigh_op_lft_6')
// (3, 13, 'sp4_v_b_29')
// (3, 14, 'neigh_op_bnl_6')
// (3, 14, 'sp4_v_b_16')
// (3, 15, 'sp4_h_r_11')
// (3, 15, 'sp4_v_b_5')
// (4, 15, 'local_g1_6')
// (4, 15, 'lutff_6/in_3')
// (4, 15, 'sp4_h_r_22')
// (5, 15, 'sp4_h_r_35')
// (6, 15, 'sp4_h_r_46')
// (7, 15, 'sp4_h_l_46')

wire n276;
// (1, 12, 'sp4_r_v_b_41')
// (1, 13, 'sp4_r_v_b_28')
// (1, 14, 'neigh_op_tnr_2')
// (1, 14, 'sp4_r_v_b_17')
// (1, 15, 'neigh_op_rgt_2')
// (1, 15, 'sp4_r_v_b_4')
// (1, 16, 'neigh_op_bnr_2')
// (2, 11, 'sp4_v_t_41')
// (2, 12, 'sp4_v_b_41')
// (2, 13, 'local_g3_4')
// (2, 13, 'lutff_6/in_3')
// (2, 13, 'sp4_v_b_28')
// (2, 14, 'neigh_op_top_2')
// (2, 14, 'sp4_v_b_17')
// (2, 15, 'lutff_2/out')
// (2, 15, 'sp4_v_b_4')
// (2, 16, 'neigh_op_bot_2')
// (3, 14, 'neigh_op_tnl_2')
// (3, 15, 'neigh_op_lft_2')
// (3, 16, 'neigh_op_bnl_2')

reg n277 = 0;
// (1, 12, 'sp4_r_v_b_46')
// (1, 13, 'sp4_r_v_b_35')
// (1, 14, 'sp4_r_v_b_22')
// (1, 15, 'sp4_r_v_b_11')
// (2, 11, 'sp4_v_t_46')
// (2, 12, 'sp4_h_r_10')
// (2, 12, 'sp4_v_b_46')
// (2, 13, 'sp4_v_b_35')
// (2, 14, 'local_g0_6')
// (2, 14, 'lutff_3/in_3')
// (2, 14, 'sp4_v_b_22')
// (2, 15, 'sp4_h_r_11')
// (2, 15, 'sp4_v_b_11')
// (3, 12, 'local_g1_7')
// (3, 12, 'lutff_4/in_0')
// (3, 12, 'sp4_h_r_23')
// (3, 12, 'sp4_r_v_b_41')
// (3, 13, 'sp4_r_v_b_28')
// (3, 14, 'sp4_r_v_b_17')
// (3, 15, 'sp4_h_r_22')
// (3, 15, 'sp4_r_v_b_4')
// (3, 20, 'local_g1_1')
// (3, 20, 'lutff_4/in_2')
// (3, 20, 'sp4_h_r_9')
// (3, 21, 'local_g0_7')
// (3, 21, 'lutff_0/in_3')
// (3, 21, 'lutff_3/in_2')
// (3, 21, 'lutff_6/in_1')
// (3, 21, 'sp4_h_r_7')
// (4, 11, 'sp4_v_t_41')
// (4, 12, 'sp4_h_r_34')
// (4, 12, 'sp4_v_b_41')
// (4, 13, 'sp4_v_b_28')
// (4, 14, 'local_g0_1')
// (4, 14, 'lutff_7/in_0')
// (4, 14, 'sp4_v_b_17')
// (4, 15, 'sp4_h_r_35')
// (4, 15, 'sp4_h_r_4')
// (4, 15, 'sp4_v_b_4')
// (4, 20, 'sp4_h_r_20')
// (4, 21, 'sp4_h_r_18')
// (5, 12, 'sp4_h_r_47')
// (5, 15, 'sp4_h_r_17')
// (5, 15, 'sp4_h_r_46')
// (5, 20, 'sp4_h_r_33')
// (5, 21, 'sp4_h_r_31')
// (6, 11, 'sp4_h_r_2')
// (6, 12, 'sp4_h_l_47')
// (6, 12, 'sp4_h_r_10')
// (6, 15, 'sp4_h_l_46')
// (6, 15, 'sp4_h_r_28')
// (6, 15, 'sp4_h_r_8')
// (6, 20, 'sp4_h_r_44')
// (6, 21, 'sp4_h_r_42')
// (7, 11, 'local_g1_7')
// (7, 11, 'lutff_6/in_0')
// (7, 11, 'sp4_h_r_15')
// (7, 12, 'sp4_h_r_23')
// (7, 15, 'sp4_h_r_21')
// (7, 15, 'sp4_h_r_41')
// (7, 16, 'sp4_r_v_b_47')
// (7, 17, 'sp4_r_v_b_34')
// (7, 18, 'sp4_r_v_b_23')
// (7, 19, 'sp4_r_v_b_10')
// (7, 20, 'sp4_h_l_44')
// (7, 20, 'sp4_h_r_6')
// (7, 21, 'local_g0_3')
// (7, 21, 'lutff_4/in_1')
// (7, 21, 'sp4_h_l_42')
// (7, 21, 'sp4_h_r_11')
// (8, 11, 'sp4_h_r_26')
// (8, 12, 'sp4_h_r_34')
// (8, 15, 'sp4_h_l_41')
// (8, 15, 'sp4_h_r_32')
// (8, 15, 'sp4_v_t_47')
// (8, 16, 'sp4_v_b_47')
// (8, 17, 'sp4_v_b_34')
// (8, 18, 'sp4_v_b_23')
// (8, 19, 'sp4_h_r_10')
// (8, 19, 'sp4_v_b_10')
// (8, 20, 'sp4_h_r_19')
// (8, 21, 'sp4_h_r_22')
// (9, 11, 'sp4_h_r_39')
// (9, 12, 'sp4_h_r_47')
// (9, 12, 'sp4_r_v_b_39')
// (9, 13, 'sp4_r_v_b_26')
// (9, 13, 'sp4_r_v_b_47')
// (9, 14, 'sp4_r_v_b_15')
// (9, 14, 'sp4_r_v_b_34')
// (9, 15, 'sp4_h_r_45')
// (9, 15, 'sp4_r_v_b_2')
// (9, 15, 'sp4_r_v_b_23')
// (9, 16, 'sp4_r_v_b_10')
// (9, 16, 'sp4_r_v_b_39')
// (9, 17, 'local_g0_2')
// (9, 17, 'lutff_4/in_0')
// (9, 17, 'lutff_5/in_3')
// (9, 17, 'sp4_r_v_b_26')
// (9, 17, 'sp4_r_v_b_42')
// (9, 18, 'neigh_op_tnr_1')
// (9, 18, 'sp4_r_v_b_15')
// (9, 18, 'sp4_r_v_b_31')
// (9, 19, 'neigh_op_rgt_1')
// (9, 19, 'sp4_h_r_23')
// (9, 19, 'sp4_r_v_b_18')
// (9, 19, 'sp4_r_v_b_2')
// (9, 20, 'neigh_op_bnr_1')
// (9, 20, 'sp4_h_r_30')
// (9, 20, 'sp4_r_v_b_7')
// (9, 21, 'sp4_h_r_35')
// (10, 11, 'sp4_h_l_39')
// (10, 11, 'sp4_h_r_2')
// (10, 11, 'sp4_v_t_39')
// (10, 12, 'sp4_h_l_47')
// (10, 12, 'sp4_v_b_39')
// (10, 12, 'sp4_v_t_47')
// (10, 13, 'sp4_v_b_26')
// (10, 13, 'sp4_v_b_47')
// (10, 14, 'sp4_v_b_15')
// (10, 14, 'sp4_v_b_34')
// (10, 15, 'sp4_h_l_45')
// (10, 15, 'sp4_v_b_2')
// (10, 15, 'sp4_v_b_23')
// (10, 15, 'sp4_v_t_39')
// (10, 16, 'sp4_r_v_b_38')
// (10, 16, 'sp4_v_b_10')
// (10, 16, 'sp4_v_b_39')
// (10, 16, 'sp4_v_t_42')
// (10, 17, 'sp4_r_v_b_27')
// (10, 17, 'sp4_r_v_b_43')
// (10, 17, 'sp4_v_b_26')
// (10, 17, 'sp4_v_b_42')
// (10, 18, 'neigh_op_top_1')
// (10, 18, 'sp4_r_v_b_14')
// (10, 18, 'sp4_r_v_b_30')
// (10, 18, 'sp4_r_v_b_46')
// (10, 18, 'sp4_v_b_15')
// (10, 18, 'sp4_v_b_31')
// (10, 19, 'local_g1_1')
// (10, 19, 'lutff_1/out')
// (10, 19, 'lutff_3/in_1')
// (10, 19, 'sp4_h_r_34')
// (10, 19, 'sp4_r_v_b_19')
// (10, 19, 'sp4_r_v_b_3')
// (10, 19, 'sp4_r_v_b_35')
// (10, 19, 'sp4_v_b_18')
// (10, 19, 'sp4_v_b_2')
// (10, 20, 'neigh_op_bot_1')
// (10, 20, 'sp4_h_r_43')
// (10, 20, 'sp4_r_v_b_22')
// (10, 20, 'sp4_r_v_b_6')
// (10, 20, 'sp4_v_b_7')
// (10, 21, 'sp4_h_r_46')
// (10, 21, 'sp4_r_v_b_11')
// (11, 11, 'local_g1_7')
// (11, 11, 'lutff_5/in_1')
// (11, 11, 'sp4_h_r_15')
// (11, 15, 'sp4_v_t_38')
// (11, 16, 'sp4_v_b_38')
// (11, 16, 'sp4_v_t_43')
// (11, 17, 'local_g3_3')
// (11, 17, 'lutff_2/in_0')
// (11, 17, 'sp4_v_b_27')
// (11, 17, 'sp4_v_b_43')
// (11, 17, 'sp4_v_t_46')
// (11, 18, 'neigh_op_tnl_1')
// (11, 18, 'sp4_v_b_14')
// (11, 18, 'sp4_v_b_30')
// (11, 18, 'sp4_v_b_46')
// (11, 19, 'neigh_op_lft_1')
// (11, 19, 'sp4_h_r_47')
// (11, 19, 'sp4_v_b_19')
// (11, 19, 'sp4_v_b_3')
// (11, 19, 'sp4_v_b_35')
// (11, 20, 'neigh_op_bnl_1')
// (11, 20, 'sp4_h_l_43')
// (11, 20, 'sp4_v_b_22')
// (11, 20, 'sp4_v_b_6')
// (11, 21, 'sp4_h_l_46')
// (11, 21, 'sp4_v_b_11')
// (12, 11, 'sp4_h_r_26')
// (12, 19, 'sp4_h_l_47')
// (13, 11, 'sp4_h_r_39')
// (14, 11, 'sp4_h_l_39')

wire n278;
// (1, 13, 'local_g0_4')
// (1, 13, 'lutff_4/in_2')
// (1, 13, 'sp4_h_r_4')
// (2, 12, 'neigh_op_tnr_6')
// (2, 13, 'neigh_op_rgt_6')
// (2, 13, 'sp4_h_r_17')
// (2, 14, 'neigh_op_bnr_6')
// (3, 12, 'neigh_op_top_6')
// (3, 13, 'lutff_6/out')
// (3, 13, 'sp4_h_r_28')
// (3, 14, 'neigh_op_bot_6')
// (4, 12, 'neigh_op_tnl_6')
// (4, 13, 'neigh_op_lft_6')
// (4, 13, 'sp4_h_r_41')
// (4, 14, 'neigh_op_bnl_6')
// (5, 13, 'sp4_h_l_41')

wire n279;
// (1, 13, 'lutff_1/cout')
// (1, 13, 'lutff_2/in_3')

reg n280 = 0;
// (1, 13, 'neigh_op_tnr_1')
// (1, 14, 'neigh_op_rgt_1')
// (1, 14, 'sp4_h_r_7')
// (1, 15, 'neigh_op_bnr_1')
// (2, 12, 'sp4_r_v_b_43')
// (2, 13, 'neigh_op_top_1')
// (2, 13, 'sp4_r_v_b_30')
// (2, 13, 'sp4_r_v_b_46')
// (2, 14, 'lutff_1/out')
// (2, 14, 'sp4_h_r_18')
// (2, 14, 'sp4_r_v_b_19')
// (2, 14, 'sp4_r_v_b_35')
// (2, 15, 'neigh_op_bot_1')
// (2, 15, 'sp4_r_v_b_22')
// (2, 15, 'sp4_r_v_b_6')
// (2, 16, 'sp4_r_v_b_11')
// (2, 16, 'sp4_r_v_b_44')
// (2, 17, 'sp4_r_v_b_33')
// (2, 18, 'sp4_r_v_b_20')
// (2, 19, 'sp4_r_v_b_9')
// (3, 11, 'sp4_v_t_43')
// (3, 12, 'sp4_v_b_43')
// (3, 12, 'sp4_v_t_46')
// (3, 13, 'neigh_op_tnl_1')
// (3, 13, 'sp4_v_b_30')
// (3, 13, 'sp4_v_b_46')
// (3, 14, 'neigh_op_lft_1')
// (3, 14, 'sp4_h_r_31')
// (3, 14, 'sp4_v_b_19')
// (3, 14, 'sp4_v_b_35')
// (3, 15, 'local_g2_1')
// (3, 15, 'lutff_2/in_3')
// (3, 15, 'neigh_op_bnl_1')
// (3, 15, 'sp4_v_b_22')
// (3, 15, 'sp4_v_b_6')
// (3, 15, 'sp4_v_t_44')
// (3, 16, 'sp4_h_r_11')
// (3, 16, 'sp4_v_b_11')
// (3, 16, 'sp4_v_b_44')
// (3, 17, 'sp4_v_b_33')
// (3, 18, 'sp4_v_b_20')
// (3, 19, 'sp4_h_r_3')
// (3, 19, 'sp4_v_b_9')
// (4, 11, 'sp4_r_v_b_36')
// (4, 12, 'sp4_r_v_b_25')
// (4, 13, 'local_g2_4')
// (4, 13, 'lutff_6/in_0')
// (4, 13, 'sp4_r_v_b_12')
// (4, 14, 'sp4_h_r_42')
// (4, 14, 'sp4_r_v_b_1')
// (4, 16, 'local_g1_6')
// (4, 16, 'lutff_5/in_2')
// (4, 16, 'sp4_h_r_22')
// (4, 19, 'sp4_h_r_14')
// (5, 10, 'sp4_v_t_36')
// (5, 11, 'sp4_v_b_36')
// (5, 12, 'sp4_v_b_25')
// (5, 13, 'sp4_v_b_12')
// (5, 14, 'sp4_h_l_42')
// (5, 14, 'sp4_v_b_1')
// (5, 16, 'sp4_h_r_35')
// (5, 19, 'local_g2_3')
// (5, 19, 'lutff_1/in_0')
// (5, 19, 'sp4_h_r_27')
// (6, 16, 'sp4_h_r_46')
// (6, 19, 'sp4_h_r_38')
// (7, 16, 'sp4_h_l_46')
// (7, 19, 'sp4_h_l_38')

wire n281;
// (1, 13, 'neigh_op_tnr_2')
// (1, 14, 'local_g3_2')
// (1, 14, 'lutff_5/in_0')
// (1, 14, 'neigh_op_rgt_2')
// (1, 15, 'neigh_op_bnr_2')
// (2, 13, 'neigh_op_top_2')
// (2, 14, 'local_g2_2')
// (2, 14, 'lutff_2/out')
// (2, 14, 'lutff_3/in_1')
// (2, 14, 'lutff_6/in_2')
// (2, 15, 'neigh_op_bot_2')
// (3, 13, 'neigh_op_tnl_2')
// (3, 14, 'neigh_op_lft_2')
// (3, 15, 'neigh_op_bnl_2')

wire n282;
// (1, 13, 'neigh_op_tnr_3')
// (1, 14, 'neigh_op_rgt_3')
// (1, 15, 'neigh_op_bnr_3')
// (2, 11, 'sp4_r_v_b_42')
// (2, 12, 'local_g0_7')
// (2, 12, 'lutff_6/in_1')
// (2, 12, 'sp4_r_v_b_31')
// (2, 13, 'local_g0_3')
// (2, 13, 'lutff_4/in_1')
// (2, 13, 'neigh_op_top_3')
// (2, 13, 'sp4_r_v_b_18')
// (2, 14, 'lutff_3/out')
// (2, 14, 'sp4_r_v_b_39')
// (2, 14, 'sp4_r_v_b_7')
// (2, 15, 'local_g0_3')
// (2, 15, 'lutff_4/in_3')
// (2, 15, 'neigh_op_bot_3')
// (2, 15, 'sp4_r_v_b_26')
// (2, 16, 'sp4_r_v_b_15')
// (2, 17, 'sp4_r_v_b_2')
// (3, 10, 'sp4_v_t_42')
// (3, 11, 'sp4_v_b_42')
// (3, 12, 'sp4_v_b_31')
// (3, 13, 'neigh_op_tnl_3')
// (3, 13, 'sp4_v_b_18')
// (3, 13, 'sp4_v_t_39')
// (3, 14, 'neigh_op_lft_3')
// (3, 14, 'sp4_v_b_39')
// (3, 14, 'sp4_v_b_7')
// (3, 15, 'neigh_op_bnl_3')
// (3, 15, 'sp4_v_b_26')
// (3, 16, 'local_g0_7')
// (3, 16, 'lutff_6/in_3')
// (3, 16, 'sp4_v_b_15')
// (3, 17, 'sp4_v_b_2')

wire n283;
// (1, 13, 'neigh_op_tnr_5')
// (1, 14, 'neigh_op_rgt_5')
// (1, 15, 'neigh_op_bnr_5')
// (2, 11, 'sp4_r_v_b_46')
// (2, 12, 'sp4_r_v_b_35')
// (2, 13, 'neigh_op_top_5')
// (2, 13, 'sp4_r_v_b_22')
// (2, 14, 'lutff_5/out')
// (2, 14, 'sp4_r_v_b_11')
// (2, 15, 'neigh_op_bot_5')
// (3, 10, 'sp4_v_t_46')
// (3, 11, 'sp4_v_b_46')
// (3, 12, 'local_g2_3')
// (3, 12, 'lutff_1/in_2')
// (3, 12, 'sp4_v_b_35')
// (3, 13, 'neigh_op_tnl_5')
// (3, 13, 'sp4_v_b_22')
// (3, 14, 'neigh_op_lft_5')
// (3, 14, 'sp4_v_b_11')
// (3, 15, 'neigh_op_bnl_5')

wire n284;
// (1, 13, 'neigh_op_tnr_7')
// (1, 14, 'neigh_op_rgt_7')
// (1, 15, 'neigh_op_bnr_7')
// (2, 13, 'neigh_op_top_7')
// (2, 14, 'lutff_7/out')
// (2, 15, 'neigh_op_bot_7')
// (3, 13, 'neigh_op_tnl_7')
// (3, 14, 'local_g0_7')
// (3, 14, 'lutff_7/in_2')
// (3, 14, 'neigh_op_lft_7')
// (3, 15, 'neigh_op_bnl_7')

wire n285;
// (1, 14, 'local_g1_6')
// (1, 14, 'lutff_6/in_1')
// (1, 14, 'sp4_h_r_6')
// (2, 13, 'neigh_op_tnr_7')
// (2, 14, 'neigh_op_rgt_7')
// (2, 14, 'sp4_h_r_19')
// (2, 15, 'neigh_op_bnr_7')
// (3, 13, 'neigh_op_top_7')
// (3, 14, 'lutff_7/out')
// (3, 14, 'sp4_h_r_30')
// (3, 15, 'neigh_op_bot_7')
// (4, 13, 'neigh_op_tnl_7')
// (4, 14, 'neigh_op_lft_7')
// (4, 14, 'sp4_h_r_43')
// (4, 15, 'neigh_op_bnl_7')
// (5, 14, 'sp4_h_l_43')

wire n286;
// (1, 14, 'neigh_op_tnr_0')
// (1, 15, 'neigh_op_rgt_0')
// (1, 16, 'neigh_op_bnr_0')
// (2, 14, 'neigh_op_top_0')
// (2, 15, 'lutff_0/out')
// (2, 15, 'sp4_h_r_0')
// (2, 16, 'neigh_op_bot_0')
// (3, 14, 'neigh_op_tnl_0')
// (3, 15, 'neigh_op_lft_0')
// (3, 15, 'sp4_h_r_13')
// (3, 16, 'neigh_op_bnl_0')
// (4, 15, 'local_g3_0')
// (4, 15, 'lutff_1/in_0')
// (4, 15, 'lutff_4/in_1')
// (4, 15, 'sp4_h_r_24')
// (5, 15, 'sp4_h_r_37')
// (6, 15, 'sp4_h_l_37')

wire n287;
// (1, 14, 'neigh_op_tnr_1')
// (1, 15, 'neigh_op_rgt_1')
// (1, 16, 'neigh_op_bnr_1')
// (2, 14, 'neigh_op_top_1')
// (2, 15, 'local_g1_1')
// (2, 15, 'lutff_1/out')
// (2, 15, 'lutff_6/in_2')
// (2, 16, 'neigh_op_bot_1')
// (3, 14, 'neigh_op_tnl_1')
// (3, 15, 'local_g0_1')
// (3, 15, 'lutff_0/in_1')
// (3, 15, 'lutff_5/in_2')
// (3, 15, 'neigh_op_lft_1')
// (3, 16, 'local_g3_1')
// (3, 16, 'lutff_0/in_0')
// (3, 16, 'neigh_op_bnl_1')

reg n288 = 0;
// (1, 14, 'neigh_op_tnr_3')
// (1, 15, 'neigh_op_rgt_3')
// (1, 15, 'sp4_r_v_b_38')
// (1, 16, 'neigh_op_bnr_3')
// (1, 16, 'sp4_r_v_b_27')
// (1, 17, 'local_g2_6')
// (1, 17, 'lutff_5/in_1')
// (1, 17, 'sp4_r_v_b_14')
// (1, 18, 'sp4_r_v_b_3')
// (2, 14, 'local_g0_3')
// (2, 14, 'lutff_2/in_1')
// (2, 14, 'lutff_7/in_0')
// (2, 14, 'neigh_op_top_3')
// (2, 14, 'sp4_v_t_38')
// (2, 15, 'local_g2_3')
// (2, 15, 'lutff_3/out')
// (2, 15, 'lutff_4/in_1')
// (2, 15, 'sp4_v_b_38')
// (2, 16, 'neigh_op_bot_3')
// (2, 16, 'sp4_v_b_27')
// (2, 17, 'sp4_v_b_14')
// (2, 18, 'sp4_v_b_3')
// (3, 14, 'local_g2_3')
// (3, 14, 'lutff_4/in_1')
// (3, 14, 'neigh_op_tnl_3')
// (3, 15, 'local_g0_3')
// (3, 15, 'lutff_3/in_0')
// (3, 15, 'neigh_op_lft_3')
// (3, 16, 'neigh_op_bnl_3')

wire n289;
// (1, 14, 'neigh_op_tnr_4')
// (1, 15, 'neigh_op_rgt_4')
// (1, 16, 'neigh_op_bnr_4')
// (2, 14, 'neigh_op_top_4')
// (2, 15, 'local_g3_4')
// (2, 15, 'lutff_3/in_2')
// (2, 15, 'lutff_4/out')
// (2, 16, 'neigh_op_bot_4')
// (3, 14, 'neigh_op_tnl_4')
// (3, 15, 'neigh_op_lft_4')
// (3, 16, 'neigh_op_bnl_4')

reg n290 = 0;
// (1, 14, 'neigh_op_tnr_6')
// (1, 15, 'neigh_op_rgt_6')
// (1, 16, 'neigh_op_bnr_6')
// (2, 14, 'neigh_op_top_6')
// (2, 15, 'local_g0_6')
// (2, 15, 'local_g3_6')
// (2, 15, 'lutff_6/in_1')
// (2, 15, 'lutff_6/out')
// (2, 15, 'lutff_7/in_3')
// (2, 16, 'neigh_op_bot_6')
// (3, 14, 'neigh_op_tnl_6')
// (3, 15, 'neigh_op_lft_6')
// (3, 16, 'neigh_op_bnl_6')

wire n291;
// (1, 14, 'sp4_r_v_b_38')
// (1, 15, 'neigh_op_tnr_7')
// (1, 15, 'sp4_r_v_b_27')
// (1, 16, 'neigh_op_rgt_7')
// (1, 16, 'sp4_r_v_b_14')
// (1, 17, 'neigh_op_bnr_7')
// (1, 17, 'sp4_r_v_b_3')
// (2, 13, 'sp4_v_t_38')
// (2, 14, 'sp4_v_b_38')
// (2, 15, 'neigh_op_top_7')
// (2, 15, 'sp4_v_b_27')
// (2, 16, 'lutff_7/out')
// (2, 16, 'sp4_v_b_14')
// (2, 17, 'neigh_op_bot_7')
// (2, 17, 'sp4_h_r_9')
// (2, 17, 'sp4_v_b_3')
// (3, 15, 'neigh_op_tnl_7')
// (3, 16, 'neigh_op_lft_7')
// (3, 17, 'neigh_op_bnl_7')
// (3, 17, 'sp4_h_r_20')
// (4, 17, 'local_g2_1')
// (4, 17, 'lutff_3/in_0')
// (4, 17, 'sp4_h_r_33')
// (5, 17, 'sp4_h_r_44')
// (6, 17, 'sp4_h_l_44')

wire n292;
// (1, 15, 'neigh_op_tnr_0')
// (1, 16, 'neigh_op_rgt_0')
// (1, 17, 'neigh_op_bnr_0')
// (2, 14, 'sp4_r_v_b_41')
// (2, 15, 'neigh_op_top_0')
// (2, 15, 'sp4_r_v_b_28')
// (2, 16, 'lutff_0/out')
// (2, 16, 'sp4_r_v_b_17')
// (2, 17, 'neigh_op_bot_0')
// (2, 17, 'sp4_r_v_b_4')
// (3, 13, 'sp4_v_t_41')
// (3, 14, 'sp4_v_b_41')
// (3, 15, 'neigh_op_tnl_0')
// (3, 15, 'sp4_v_b_28')
// (3, 16, 'neigh_op_lft_0')
// (3, 16, 'sp4_v_b_17')
// (3, 17, 'neigh_op_bnl_0')
// (3, 17, 'sp4_h_r_10')
// (3, 17, 'sp4_h_r_4')
// (3, 17, 'sp4_v_b_4')
// (4, 17, 'local_g1_1')
// (4, 17, 'lutff_4/in_0')
// (4, 17, 'sp4_h_r_17')
// (4, 17, 'sp4_h_r_23')
// (5, 17, 'local_g2_2')
// (5, 17, 'lutff_0/in_0')
// (5, 17, 'sp4_h_r_28')
// (5, 17, 'sp4_h_r_34')
// (6, 17, 'sp4_h_r_41')
// (6, 17, 'sp4_h_r_47')
// (7, 17, 'sp4_h_l_41')
// (7, 17, 'sp4_h_l_47')

wire n293;
// (1, 15, 'neigh_op_tnr_1')
// (1, 16, 'neigh_op_rgt_1')
// (1, 17, 'neigh_op_bnr_1')
// (2, 15, 'neigh_op_top_1')
// (2, 16, 'local_g1_1')
// (2, 16, 'lutff_0/in_0')
// (2, 16, 'lutff_1/out')
// (2, 16, 'lutff_4/in_2')
// (2, 16, 'lutff_7/in_1')
// (2, 17, 'neigh_op_bot_1')
// (3, 15, 'neigh_op_tnl_1')
// (3, 16, 'neigh_op_lft_1')
// (3, 17, 'neigh_op_bnl_1')

reg n294 = 0;
// (1, 15, 'neigh_op_tnr_3')
// (1, 16, 'local_g2_3')
// (1, 16, 'local_g3_3')
// (1, 16, 'lutff_0/in_1')
// (1, 16, 'lutff_1/in_3')
// (1, 16, 'neigh_op_rgt_3')
// (1, 17, 'neigh_op_bnr_3')
// (2, 15, 'neigh_op_top_3')
// (2, 16, 'local_g2_3')
// (2, 16, 'local_g3_3')
// (2, 16, 'lutff_0/in_2')
// (2, 16, 'lutff_3/in_1')
// (2, 16, 'lutff_3/out')
// (2, 16, 'lutff_4/in_3')
// (2, 17, 'neigh_op_bot_3')
// (3, 15, 'neigh_op_tnl_3')
// (3, 16, 'neigh_op_lft_3')
// (3, 17, 'neigh_op_bnl_3')

wire n295;
// (1, 15, 'neigh_op_tnr_4')
// (1, 16, 'neigh_op_rgt_4')
// (1, 17, 'neigh_op_bnr_4')
// (2, 15, 'neigh_op_top_4')
// (2, 16, 'lutff_4/out')
// (2, 17, 'local_g1_4')
// (2, 17, 'lutff_5/in_2')
// (2, 17, 'neigh_op_bot_4')
// (3, 15, 'neigh_op_tnl_4')
// (3, 16, 'neigh_op_lft_4')
// (3, 17, 'local_g3_4')
// (3, 17, 'lutff_3/in_0')
// (3, 17, 'neigh_op_bnl_4')

reg n296 = 0;
// (1, 15, 'sp4_r_v_b_36')
// (1, 16, 'sp4_r_v_b_25')
// (1, 17, 'sp4_r_v_b_12')
// (1, 18, 'sp4_r_v_b_1')
// (2, 14, 'sp4_h_r_7')
// (2, 14, 'sp4_v_t_36')
// (2, 15, 'local_g2_4')
// (2, 15, 'lutff_2/in_0')
// (2, 15, 'sp4_v_b_36')
// (2, 16, 'sp4_v_b_25')
// (2, 17, 'sp4_v_b_12')
// (2, 18, 'sp4_v_b_1')
// (3, 14, 'sp4_h_r_18')
// (4, 13, 'neigh_op_tnr_5')
// (4, 14, 'neigh_op_rgt_5')
// (4, 14, 'sp4_h_r_31')
// (4, 15, 'neigh_op_bnr_5')
// (5, 13, 'neigh_op_top_5')
// (5, 14, 'local_g1_5')
// (5, 14, 'local_g2_5')
// (5, 14, 'lutff_4/in_0')
// (5, 14, 'lutff_5/in_2')
// (5, 14, 'lutff_5/out')
// (5, 14, 'sp4_h_r_42')
// (5, 15, 'local_g0_5')
// (5, 15, 'lutff_1/in_0')
// (5, 15, 'neigh_op_bot_5')
// (6, 13, 'neigh_op_tnl_5')
// (6, 14, 'neigh_op_lft_5')
// (6, 14, 'sp4_h_l_42')
// (6, 15, 'neigh_op_bnl_5')

reg n297 = 0;
// (1, 15, 'sp4_r_v_b_45')
// (1, 16, 'sp4_r_v_b_32')
// (1, 17, 'sp4_r_v_b_21')
// (1, 18, 'sp4_r_v_b_8')
// (2, 14, 'local_g0_0')
// (2, 14, 'lutff_5/in_1')
// (2, 14, 'sp4_h_r_8')
// (2, 14, 'sp4_v_t_45')
// (2, 15, 'local_g3_5')
// (2, 15, 'lutff_2/in_2')
// (2, 15, 'sp4_v_b_45')
// (2, 16, 'sp4_v_b_32')
// (2, 17, 'sp4_v_b_21')
// (2, 18, 'sp4_v_b_8')
// (3, 11, 'sp4_r_v_b_37')
// (3, 12, 'sp4_r_v_b_24')
// (3, 13, 'neigh_op_tnr_0')
// (3, 13, 'sp4_r_v_b_13')
// (3, 14, 'neigh_op_rgt_0')
// (3, 14, 'sp4_h_r_21')
// (3, 14, 'sp4_r_v_b_0')
// (3, 15, 'neigh_op_bnr_0')
// (4, 10, 'sp4_v_t_37')
// (4, 11, 'local_g2_5')
// (4, 11, 'lutff_3/in_0')
// (4, 11, 'sp4_v_b_37')
// (4, 12, 'sp4_v_b_24')
// (4, 13, 'neigh_op_top_0')
// (4, 13, 'sp4_v_b_13')
// (4, 14, 'local_g1_0')
// (4, 14, 'lutff_0/in_1')
// (4, 14, 'lutff_0/out')
// (4, 14, 'lutff_1/in_2')
// (4, 14, 'sp4_h_r_32')
// (4, 14, 'sp4_v_b_0')
// (4, 15, 'neigh_op_bot_0')
// (5, 13, 'neigh_op_tnl_0')
// (5, 14, 'neigh_op_lft_0')
// (5, 14, 'sp4_h_r_45')
// (5, 15, 'neigh_op_bnl_0')
// (6, 14, 'sp4_h_l_45')

wire n298;
// (1, 16, 'lutff_1/cout')
// (1, 16, 'lutff_2/in_3')

wire n299;
// (1, 16, 'neigh_op_tnr_2')
// (1, 17, 'neigh_op_rgt_2')
// (1, 18, 'neigh_op_bnr_2')
// (2, 16, 'neigh_op_top_2')
// (2, 17, 'lutff_2/out')
// (2, 17, 'sp4_h_r_4')
// (2, 18, 'neigh_op_bot_2')
// (3, 16, 'neigh_op_tnl_2')
// (3, 17, 'neigh_op_lft_2')
// (3, 17, 'sp4_h_r_17')
// (3, 18, 'neigh_op_bnl_2')
// (4, 17, 'local_g3_4')
// (4, 17, 'lutff_7/in_0')
// (4, 17, 'sp4_h_r_28')
// (5, 17, 'sp4_h_r_41')
// (6, 17, 'sp4_h_l_41')

reg n300 = 0;
// (1, 16, 'neigh_op_tnr_3')
// (1, 17, 'neigh_op_rgt_3')
// (1, 17, 'sp4_r_v_b_38')
// (1, 18, 'neigh_op_bnr_3')
// (1, 18, 'sp4_r_v_b_27')
// (1, 19, 'sp4_r_v_b_14')
// (1, 20, 'sp4_r_v_b_3')
// (2, 16, 'neigh_op_top_3')
// (2, 16, 'sp4_v_t_38')
// (2, 17, 'local_g2_3')
// (2, 17, 'lutff_3/in_2')
// (2, 17, 'lutff_3/out')
// (2, 17, 'sp4_v_b_38')
// (2, 18, 'local_g1_3')
// (2, 18, 'lutff_0/in_2')
// (2, 18, 'lutff_1/in_3')
// (2, 18, 'lutff_3/in_1')
// (2, 18, 'neigh_op_bot_3')
// (2, 18, 'sp4_v_b_27')
// (2, 19, 'local_g0_6')
// (2, 19, 'lutff_5/in_1')
// (2, 19, 'sp4_v_b_14')
// (2, 20, 'sp4_v_b_3')
// (3, 16, 'neigh_op_tnl_3')
// (3, 17, 'local_g0_3')
// (3, 17, 'lutff_3/in_2')
// (3, 17, 'neigh_op_lft_3')
// (3, 18, 'local_g3_3')
// (3, 18, 'lutff_3/in_1')
// (3, 18, 'neigh_op_bnl_3')

wire n301;
// (1, 16, 'neigh_op_tnr_6')
// (1, 17, 'neigh_op_rgt_6')
// (1, 18, 'local_g0_6')
// (1, 18, 'lutff_0/in_2')
// (1, 18, 'neigh_op_bnr_6')
// (2, 16, 'neigh_op_top_6')
// (2, 17, 'lutff_6/out')
// (2, 18, 'local_g1_6')
// (2, 18, 'lutff_2/in_3')
// (2, 18, 'neigh_op_bot_6')
// (3, 16, 'neigh_op_tnl_6')
// (3, 17, 'neigh_op_lft_6')
// (3, 18, 'local_g3_6')
// (3, 18, 'lutff_4/in_3')
// (3, 18, 'neigh_op_bnl_6')

wire n302;
// (1, 16, 'neigh_op_tnr_7')
// (1, 17, 'neigh_op_rgt_7')
// (1, 17, 'sp4_h_r_3')
// (1, 18, 'neigh_op_bnr_7')
// (2, 16, 'neigh_op_top_7')
// (2, 17, 'lutff_7/out')
// (2, 17, 'sp4_h_r_14')
// (2, 18, 'neigh_op_bot_7')
// (3, 16, 'neigh_op_tnl_7')
// (3, 17, 'neigh_op_lft_7')
// (3, 17, 'sp4_h_r_27')
// (3, 18, 'neigh_op_bnl_7')
// (4, 17, 'sp4_h_r_38')
// (5, 17, 'sp4_h_l_38')
// (5, 17, 'sp4_h_r_11')
// (6, 17, 'sp4_h_r_22')
// (7, 17, 'local_g3_3')
// (7, 17, 'lutff_1/in_1')
// (7, 17, 'lutff_2/in_2')
// (7, 17, 'lutff_4/in_0')
// (7, 17, 'sp4_h_r_35')
// (8, 17, 'sp4_h_r_46')
// (9, 17, 'sp4_h_l_46')

reg n303 = 0;
// (1, 16, 'sp4_h_r_2')
// (2, 15, 'neigh_op_tnr_5')
// (2, 16, 'neigh_op_rgt_5')
// (2, 16, 'sp4_h_r_15')
// (2, 16, 'sp4_r_v_b_42')
// (2, 17, 'neigh_op_bnr_5')
// (2, 17, 'sp4_r_v_b_31')
// (2, 18, 'local_g3_2')
// (2, 18, 'lutff_7/in_0')
// (2, 18, 'sp4_r_v_b_18')
// (2, 19, 'sp4_r_v_b_7')
// (3, 15, 'local_g0_5')
// (3, 15, 'lutff_2/in_1')
// (3, 15, 'lutff_6/in_3')
// (3, 15, 'neigh_op_top_5')
// (3, 15, 'sp4_v_t_42')
// (3, 16, 'local_g0_5')
// (3, 16, 'local_g3_5')
// (3, 16, 'lutff_1/in_2')
// (3, 16, 'lutff_2/in_2')
// (3, 16, 'lutff_5/in_0')
// (3, 16, 'lutff_5/out')
// (3, 16, 'sp4_h_r_26')
// (3, 16, 'sp4_r_v_b_43')
// (3, 16, 'sp4_v_b_42')
// (3, 17, 'neigh_op_bot_5')
// (3, 17, 'sp4_r_v_b_30')
// (3, 17, 'sp4_v_b_31')
// (3, 18, 'sp4_r_v_b_19')
// (3, 18, 'sp4_v_b_18')
// (3, 19, 'sp4_r_v_b_6')
// (3, 19, 'sp4_v_b_7')
// (4, 13, 'sp4_r_v_b_39')
// (4, 14, 'sp4_r_v_b_26')
// (4, 15, 'local_g3_5')
// (4, 15, 'lutff_0/in_2')
// (4, 15, 'neigh_op_tnl_5')
// (4, 15, 'sp4_r_v_b_15')
// (4, 15, 'sp4_v_t_43')
// (4, 16, 'neigh_op_lft_5')
// (4, 16, 'sp4_h_r_39')
// (4, 16, 'sp4_r_v_b_2')
// (4, 16, 'sp4_v_b_43')
// (4, 17, 'neigh_op_bnl_5')
// (4, 17, 'sp4_v_b_30')
// (4, 18, 'sp4_v_b_19')
// (4, 19, 'sp4_h_r_6')
// (4, 19, 'sp4_v_b_6')
// (5, 12, 'sp4_v_t_39')
// (5, 13, 'sp4_v_b_39')
// (5, 14, 'sp4_v_b_26')
// (5, 15, 'local_g1_7')
// (5, 15, 'lutff_3/in_3')
// (5, 15, 'sp4_v_b_15')
// (5, 16, 'sp4_h_l_39')
// (5, 16, 'sp4_v_b_2')
// (5, 19, 'local_g1_3')
// (5, 19, 'lutff_1/in_1')
// (5, 19, 'sp4_h_r_19')
// (6, 19, 'sp4_h_r_30')
// (7, 19, 'sp4_h_r_43')
// (8, 19, 'sp4_h_l_43')

reg n304 = 0;
// (1, 16, 'sp4_h_r_4')
// (2, 10, 'local_g2_4')
// (2, 10, 'lutff_7/in_3')
// (2, 10, 'sp4_r_v_b_36')
// (2, 11, 'local_g1_1')
// (2, 11, 'lutff_5/in_1')
// (2, 11, 'sp4_r_v_b_25')
// (2, 12, 'sp4_r_v_b_12')
// (2, 13, 'sp4_r_v_b_1')
// (2, 14, 'sp4_r_v_b_36')
// (2, 15, 'neigh_op_tnr_6')
// (2, 15, 'sp4_r_v_b_25')
// (2, 16, 'neigh_op_rgt_6')
// (2, 16, 'sp4_h_r_1')
// (2, 16, 'sp4_h_r_17')
// (2, 16, 'sp4_r_v_b_12')
// (2, 17, 'neigh_op_bnr_6')
// (2, 17, 'sp4_r_v_b_1')
// (3, 9, 'sp4_v_t_36')
// (3, 10, 'sp4_v_b_36')
// (3, 11, 'sp4_v_b_25')
// (3, 12, 'sp4_v_b_12')
// (3, 13, 'sp4_v_b_1')
// (3, 13, 'sp4_v_t_36')
// (3, 14, 'sp4_v_b_36')
// (3, 15, 'neigh_op_top_6')
// (3, 15, 'sp4_r_v_b_40')
// (3, 15, 'sp4_v_b_25')
// (3, 16, 'local_g2_6')
// (3, 16, 'lutff_6/in_2')
// (3, 16, 'lutff_6/out')
// (3, 16, 'sp4_h_r_12')
// (3, 16, 'sp4_h_r_28')
// (3, 16, 'sp4_r_v_b_29')
// (3, 16, 'sp4_v_b_12')
// (3, 17, 'neigh_op_bot_6')
// (3, 17, 'sp4_r_v_b_16')
// (3, 17, 'sp4_v_b_1')
// (3, 18, 'sp4_r_v_b_5')
// (4, 14, 'sp4_h_r_10')
// (4, 14, 'sp4_v_t_40')
// (4, 15, 'neigh_op_tnl_6')
// (4, 15, 'sp4_v_b_40')
// (4, 16, 'neigh_op_lft_6')
// (4, 16, 'sp4_h_r_25')
// (4, 16, 'sp4_h_r_41')
// (4, 16, 'sp4_v_b_29')
// (4, 17, 'neigh_op_bnl_6')
// (4, 17, 'sp4_r_v_b_44')
// (4, 17, 'sp4_v_b_16')
// (4, 18, 'sp4_r_v_b_33')
// (4, 18, 'sp4_v_b_5')
// (4, 19, 'sp4_r_v_b_20')
// (4, 20, 'sp4_r_v_b_9')
// (5, 14, 'sp4_h_r_23')
// (5, 16, 'local_g3_4')
// (5, 16, 'lutff_4/in_1')
// (5, 16, 'sp4_h_l_41')
// (5, 16, 'sp4_h_r_36')
// (5, 16, 'sp4_v_t_44')
// (5, 17, 'local_g2_4')
// (5, 17, 'lutff_0/in_2')
// (5, 17, 'lutff_4/in_0')
// (5, 17, 'sp4_v_b_44')
// (5, 18, 'sp4_v_b_33')
// (5, 19, 'sp4_v_b_20')
// (5, 20, 'sp4_v_b_9')
// (6, 14, 'sp4_h_r_34')
// (6, 16, 'sp4_h_l_36')
// (7, 14, 'local_g2_7')
// (7, 14, 'lutff_0/in_3')
// (7, 14, 'lutff_4/in_3')
// (7, 14, 'lutff_6/in_3')
// (7, 14, 'sp4_h_r_47')
// (8, 14, 'sp4_h_l_47')

wire n305;
// (1, 16, 'sp4_r_v_b_36')
// (1, 17, 'neigh_op_tnr_6')
// (1, 17, 'sp4_r_v_b_25')
// (1, 18, 'neigh_op_rgt_6')
// (1, 18, 'sp4_r_v_b_12')
// (1, 19, 'neigh_op_bnr_6')
// (1, 19, 'sp4_r_v_b_1')
// (2, 15, 'sp4_h_r_1')
// (2, 15, 'sp4_v_t_36')
// (2, 16, 'sp4_v_b_36')
// (2, 17, 'neigh_op_top_6')
// (2, 17, 'sp4_v_b_25')
// (2, 18, 'lutff_6/out')
// (2, 18, 'sp4_v_b_12')
// (2, 19, 'neigh_op_bot_6')
// (2, 19, 'sp4_v_b_1')
// (3, 15, 'local_g1_4')
// (3, 15, 'lutff_7/in_0')
// (3, 15, 'sp4_h_r_12')
// (3, 17, 'neigh_op_tnl_6')
// (3, 18, 'neigh_op_lft_6')
// (3, 19, 'neigh_op_bnl_6')
// (4, 15, 'sp4_h_r_25')
// (5, 15, 'sp4_h_r_36')
// (6, 15, 'sp4_h_l_36')

wire n306;
// (1, 16, 'sp4_r_v_b_43')
// (1, 17, 'local_g1_6')
// (1, 17, 'lutff_5/in_2')
// (1, 17, 'sp4_r_v_b_30')
// (1, 18, 'neigh_op_tnr_3')
// (1, 18, 'sp4_r_v_b_19')
// (1, 19, 'neigh_op_rgt_3')
// (1, 19, 'sp4_r_v_b_6')
// (1, 20, 'neigh_op_bnr_3')
// (2, 15, 'sp4_v_t_43')
// (2, 16, 'sp4_v_b_43')
// (2, 17, 'sp4_v_b_30')
// (2, 18, 'local_g0_3')
// (2, 18, 'lutff_4/in_3')
// (2, 18, 'neigh_op_top_3')
// (2, 18, 'sp4_v_b_19')
// (2, 19, 'lutff_3/out')
// (2, 19, 'sp4_v_b_6')
// (2, 20, 'local_g1_3')
// (2, 20, 'lutff_5/in_3')
// (2, 20, 'neigh_op_bot_3')
// (3, 18, 'neigh_op_tnl_3')
// (3, 19, 'neigh_op_lft_3')
// (3, 20, 'neigh_op_bnl_3')

wire n307;
// (1, 17, 'local_g3_5')
// (1, 17, 'lutff_2/in_0')
// (1, 17, 'lutff_4/in_2')
// (1, 17, 'lutff_7/in_1')
// (1, 17, 'neigh_op_tnr_5')
// (1, 18, 'local_g3_5')
// (1, 18, 'lutff_5/in_3')
// (1, 18, 'neigh_op_rgt_5')
// (1, 19, 'neigh_op_bnr_5')
// (2, 17, 'local_g1_5')
// (2, 17, 'lutff_3/in_3')
// (2, 17, 'neigh_op_top_5')
// (2, 18, 'lutff_5/out')
// (2, 19, 'local_g0_5')
// (2, 19, 'local_g1_5')
// (2, 19, 'lutff_1/in_0')
// (2, 19, 'lutff_2/in_2')
// (2, 19, 'lutff_5/in_3')
// (2, 19, 'lutff_6/in_0')
// (2, 19, 'neigh_op_bot_5')
// (3, 17, 'neigh_op_tnl_5')
// (3, 18, 'neigh_op_lft_5')
// (3, 19, 'neigh_op_bnl_5')

wire n308;
// (1, 17, 'lutff_1/cout')
// (1, 17, 'lutff_2/in_3')

reg n309 = 0;
// (1, 17, 'neigh_op_tnr_0')
// (1, 18, 'neigh_op_rgt_0')
// (1, 19, 'neigh_op_bnr_0')
// (2, 17, 'neigh_op_top_0')
// (2, 18, 'local_g1_0')
// (2, 18, 'lutff_0/in_1')
// (2, 18, 'lutff_0/out')
// (2, 18, 'sp4_h_r_0')
// (2, 19, 'neigh_op_bot_0')
// (3, 17, 'neigh_op_tnl_0')
// (3, 18, 'local_g0_0')
// (3, 18, 'local_g1_5')
// (3, 18, 'lutff_0/in_2')
// (3, 18, 'lutff_1/in_3')
// (3, 18, 'lutff_6/in_2')
// (3, 18, 'neigh_op_lft_0')
// (3, 18, 'sp4_h_r_13')
// (3, 19, 'neigh_op_bnl_0')
// (4, 18, 'sp4_h_r_24')
// (5, 18, 'sp4_h_r_37')
// (6, 18, 'sp4_h_l_37')

wire n310;
// (1, 17, 'neigh_op_tnr_1')
// (1, 18, 'neigh_op_rgt_1')
// (1, 18, 'sp4_h_r_7')
// (1, 19, 'neigh_op_bnr_1')
// (2, 16, 'sp4_r_v_b_43')
// (2, 17, 'neigh_op_top_1')
// (2, 17, 'sp4_r_v_b_30')
// (2, 18, 'local_g0_2')
// (2, 18, 'lutff_1/out')
// (2, 18, 'lutff_global/cen')
// (2, 18, 'sp4_h_r_18')
// (2, 18, 'sp4_r_v_b_19')
// (2, 19, 'neigh_op_bot_1')
// (2, 19, 'sp4_r_v_b_6')
// (3, 15, 'sp4_v_t_43')
// (3, 16, 'sp4_v_b_43')
// (3, 17, 'neigh_op_tnl_1')
// (3, 17, 'sp4_v_b_30')
// (3, 18, 'local_g1_3')
// (3, 18, 'lutff_global/cen')
// (3, 18, 'neigh_op_lft_1')
// (3, 18, 'sp4_h_r_31')
// (3, 18, 'sp4_v_b_19')
// (3, 19, 'neigh_op_bnl_1')
// (3, 19, 'sp4_v_b_6')
// (4, 18, 'sp4_h_r_42')
// (5, 18, 'sp4_h_l_42')

wire n311;
// (1, 17, 'neigh_op_tnr_2')
// (1, 18, 'neigh_op_rgt_2')
// (1, 19, 'neigh_op_bnr_2')
// (2, 17, 'neigh_op_top_2')
// (2, 18, 'local_g2_2')
// (2, 18, 'lutff_1/in_1')
// (2, 18, 'lutff_2/out')
// (2, 19, 'neigh_op_bot_2')
// (3, 17, 'neigh_op_tnl_2')
// (3, 18, 'neigh_op_lft_2')
// (3, 19, 'neigh_op_bnl_2')

reg n312 = 0;
// (1, 17, 'neigh_op_tnr_3')
// (1, 18, 'neigh_op_rgt_3')
// (1, 19, 'neigh_op_bnr_3')
// (2, 17, 'neigh_op_top_3')
// (2, 18, 'lutff_3/out')
// (2, 19, 'neigh_op_bot_3')
// (3, 17, 'neigh_op_tnl_3')
// (3, 18, 'local_g0_3')
// (3, 18, 'lutff_1/in_2')
// (3, 18, 'lutff_5/in_2')
// (3, 18, 'neigh_op_lft_3')
// (3, 19, 'neigh_op_bnl_3')

wire n313;
// (1, 17, 'neigh_op_tnr_4')
// (1, 18, 'neigh_op_rgt_4')
// (1, 19, 'neigh_op_bnr_4')
// (2, 17, 'neigh_op_top_4')
// (2, 18, 'lutff_4/out')
// (2, 19, 'neigh_op_bot_4')
// (3, 17, 'local_g2_4')
// (3, 17, 'lutff_3/in_3')
// (3, 17, 'neigh_op_tnl_4')
// (3, 18, 'neigh_op_lft_4')
// (3, 19, 'neigh_op_bnl_4')

wire n314;
// (1, 17, 'neigh_op_tnr_7')
// (1, 18, 'neigh_op_rgt_7')
// (1, 19, 'neigh_op_bnr_7')
// (2, 17, 'neigh_op_top_7')
// (2, 18, 'local_g2_7')
// (2, 18, 'lutff_6/in_3')
// (2, 18, 'lutff_7/out')
// (2, 19, 'neigh_op_bot_7')
// (3, 17, 'neigh_op_tnl_7')
// (3, 18, 'neigh_op_lft_7')
// (3, 19, 'neigh_op_bnl_7')

reg n315 = 0;
// (1, 17, 'sp4_h_r_11')
// (2, 17, 'local_g0_6')
// (2, 17, 'lutff_2/in_0')
// (2, 17, 'sp4_h_r_22')
// (3, 16, 'neigh_op_tnr_7')
// (3, 17, 'neigh_op_rgt_7')
// (3, 17, 'sp4_h_r_35')
// (3, 18, 'neigh_op_bnr_7')
// (4, 16, 'neigh_op_top_7')
// (4, 17, 'local_g3_7')
// (4, 17, 'lutff_1/in_3')
// (4, 17, 'lutff_7/out')
// (4, 17, 'sp4_h_r_46')
// (4, 18, 'neigh_op_bot_7')
// (5, 16, 'neigh_op_tnl_7')
// (5, 17, 'neigh_op_lft_7')
// (5, 17, 'sp4_h_l_46')
// (5, 18, 'neigh_op_bnl_7')

reg n316 = 0;
// (1, 17, 'sp4_h_r_7')
// (2, 17, 'local_g1_2')
// (2, 17, 'lutff_0/in_1')
// (2, 17, 'sp4_h_r_18')
// (3, 16, 'neigh_op_tnr_5')
// (3, 17, 'local_g2_5')
// (3, 17, 'lutff_6/in_3')
// (3, 17, 'neigh_op_rgt_5')
// (3, 17, 'sp4_h_r_31')
// (3, 18, 'neigh_op_bnr_5')
// (4, 16, 'neigh_op_top_5')
// (4, 17, 'local_g0_5')
// (4, 17, 'lutff_1/in_0')
// (4, 17, 'lutff_5/in_0')
// (4, 17, 'lutff_5/out')
// (4, 17, 'sp4_h_r_42')
// (4, 18, 'neigh_op_bot_5')
// (5, 16, 'neigh_op_tnl_5')
// (5, 17, 'neigh_op_lft_5')
// (5, 17, 'sp4_h_l_42')
// (5, 18, 'neigh_op_bnl_5')

wire n317;
// (1, 17, 'sp4_h_r_9')
// (2, 17, 'sp4_h_r_20')
// (3, 16, 'neigh_op_tnr_6')
// (3, 17, 'neigh_op_rgt_6')
// (3, 17, 'sp4_h_r_33')
// (3, 18, 'neigh_op_bnr_6')
// (4, 14, 'sp4_r_v_b_38')
// (4, 15, 'sp4_r_v_b_27')
// (4, 16, 'neigh_op_top_6')
// (4, 16, 'sp4_r_v_b_14')
// (4, 17, 'local_g1_3')
// (4, 17, 'lutff_6/out')
// (4, 17, 'lutff_global/cen')
// (4, 17, 'sp4_h_r_44')
// (4, 17, 'sp4_r_v_b_3')
// (4, 18, 'neigh_op_bot_6')
// (5, 13, 'sp4_v_t_38')
// (5, 14, 'sp4_v_b_38')
// (5, 15, 'sp4_v_b_27')
// (5, 16, 'neigh_op_tnl_6')
// (5, 16, 'sp4_v_b_14')
// (5, 17, 'neigh_op_lft_6')
// (5, 17, 'sp4_h_l_44')
// (5, 17, 'sp4_v_b_3')
// (5, 18, 'neigh_op_bnl_6')

reg n318 = 0;
// (1, 17, 'sp4_r_v_b_43')
// (1, 18, 'sp4_r_v_b_30')
// (1, 19, 'local_g2_3')
// (1, 19, 'lutff_3/in_2')
// (1, 19, 'neigh_op_tnr_3')
// (1, 19, 'sp4_r_v_b_19')
// (1, 20, 'neigh_op_rgt_3')
// (1, 20, 'sp4_r_v_b_6')
// (1, 21, 'neigh_op_bnr_3')
// (2, 16, 'sp4_v_t_43')
// (2, 17, 'sp4_r_v_b_42')
// (2, 17, 'sp4_v_b_43')
// (2, 18, 'local_g2_6')
// (2, 18, 'local_g3_6')
// (2, 18, 'lutff_0/in_0')
// (2, 18, 'lutff_1/in_0')
// (2, 18, 'lutff_3/in_3')
// (2, 18, 'lutff_6/in_1')
// (2, 18, 'sp4_r_v_b_31')
// (2, 18, 'sp4_v_b_30')
// (2, 19, 'neigh_op_top_3')
// (2, 19, 'sp4_r_v_b_18')
// (2, 19, 'sp4_v_b_19')
// (2, 20, 'local_g0_3')
// (2, 20, 'local_g3_3')
// (2, 20, 'lutff_1/in_0')
// (2, 20, 'lutff_2/in_0')
// (2, 20, 'lutff_3/out')
// (2, 20, 'sp4_r_v_b_7')
// (2, 20, 'sp4_v_b_6')
// (2, 21, 'neigh_op_bot_3')
// (3, 16, 'sp4_v_t_42')
// (3, 17, 'sp4_v_b_42')
// (3, 18, 'local_g3_7')
// (3, 18, 'lutff_3/in_3')
// (3, 18, 'sp4_v_b_31')
// (3, 19, 'neigh_op_tnl_3')
// (3, 19, 'sp4_v_b_18')
// (3, 20, 'local_g1_3')
// (3, 20, 'lutff_1/in_3')
// (3, 20, 'neigh_op_lft_3')
// (3, 20, 'sp4_v_b_7')
// (3, 21, 'neigh_op_bnl_3')

reg n319 = 0;
// (1, 18, 'neigh_op_tnr_1')
// (1, 19, 'neigh_op_rgt_1')
// (1, 20, 'neigh_op_bnr_1')
// (2, 18, 'neigh_op_top_1')
// (2, 19, 'local_g1_1')
// (2, 19, 'lutff_1/in_1')
// (2, 19, 'lutff_1/out')
// (2, 19, 'lutff_7/in_1')
// (2, 20, 'neigh_op_bot_1')
// (3, 18, 'neigh_op_tnl_1')
// (3, 19, 'neigh_op_lft_1')
// (3, 20, 'neigh_op_bnl_1')

reg n320 = 0;
// (1, 18, 'neigh_op_tnr_2')
// (1, 19, 'neigh_op_rgt_2')
// (1, 20, 'neigh_op_bnr_2')
// (2, 18, 'neigh_op_top_2')
// (2, 19, 'local_g1_2')
// (2, 19, 'lutff_2/in_1')
// (2, 19, 'lutff_2/out')
// (2, 19, 'lutff_7/in_2')
// (2, 20, 'neigh_op_bot_2')
// (3, 18, 'neigh_op_tnl_2')
// (3, 19, 'neigh_op_lft_2')
// (3, 20, 'neigh_op_bnl_2')

wire n321;
// (1, 18, 'neigh_op_tnr_4')
// (1, 19, 'neigh_op_rgt_4')
// (1, 20, 'neigh_op_bnr_4')
// (2, 18, 'neigh_op_top_4')
// (2, 19, 'lutff_4/out')
// (2, 20, 'neigh_op_bot_4')
// (3, 18, 'neigh_op_tnl_4')
// (3, 19, 'local_g0_4')
// (3, 19, 'lutff_6/in_2')
// (3, 19, 'neigh_op_lft_4')
// (3, 20, 'neigh_op_bnl_4')

wire n322;
// (1, 18, 'neigh_op_tnr_5')
// (1, 19, 'neigh_op_rgt_5')
// (1, 20, 'neigh_op_bnr_5')
// (2, 18, 'neigh_op_top_5')
// (2, 19, 'local_g0_2')
// (2, 19, 'lutff_5/out')
// (2, 19, 'lutff_global/cen')
// (2, 19, 'sp4_h_r_10')
// (2, 20, 'neigh_op_bot_5')
// (3, 18, 'neigh_op_tnl_5')
// (3, 19, 'neigh_op_lft_5')
// (3, 19, 'sp4_h_r_23')
// (3, 20, 'neigh_op_bnl_5')
// (4, 19, 'sp4_h_r_34')
// (5, 19, 'sp4_h_r_47')
// (6, 19, 'sp4_h_l_47')

reg n323 = 0;
// (1, 18, 'neigh_op_tnr_6')
// (1, 19, 'neigh_op_rgt_6')
// (1, 20, 'neigh_op_bnr_6')
// (2, 18, 'neigh_op_top_6')
// (2, 19, 'local_g1_6')
// (2, 19, 'local_g2_6')
// (2, 19, 'lutff_0/in_1')
// (2, 19, 'lutff_1/in_3')
// (2, 19, 'lutff_6/in_3')
// (2, 19, 'lutff_6/out')
// (2, 19, 'lutff_7/in_0')
// (2, 20, 'neigh_op_bot_6')
// (3, 18, 'neigh_op_tnl_6')
// (3, 19, 'neigh_op_lft_6')
// (3, 20, 'neigh_op_bnl_6')

reg n324 = 0;
// (1, 18, 'sp4_r_v_b_39')
// (1, 19, 'sp4_r_v_b_26')
// (1, 20, 'neigh_op_tnr_1')
// (1, 20, 'sp4_r_v_b_15')
// (1, 21, 'neigh_op_rgt_1')
// (1, 21, 'sp4_r_v_b_2')
// (1, 22, 'neigh_op_bnr_1')
// (2, 17, 'sp4_v_t_39')
// (2, 18, 'sp4_v_b_39')
// (2, 19, 'local_g3_2')
// (2, 19, 'lutff_3/in_2')
// (2, 19, 'sp4_v_b_26')
// (2, 20, 'neigh_op_top_1')
// (2, 20, 'sp4_v_b_15')
// (2, 21, 'local_g1_1')
// (2, 21, 'lutff_1/in_1')
// (2, 21, 'lutff_1/out')
// (2, 21, 'sp4_v_b_2')
// (2, 22, 'neigh_op_bot_1')
// (3, 20, 'neigh_op_tnl_1')
// (3, 21, 'neigh_op_lft_1')
// (3, 22, 'neigh_op_bnl_1')

reg n325 = 0;
// (1, 18, 'sp4_r_v_b_41')
// (1, 19, 'sp4_r_v_b_28')
// (1, 20, 'neigh_op_tnr_2')
// (1, 20, 'sp4_r_v_b_17')
// (1, 21, 'neigh_op_rgt_2')
// (1, 21, 'sp4_r_v_b_4')
// (1, 22, 'neigh_op_bnr_2')
// (2, 17, 'sp4_v_t_41')
// (2, 18, 'sp4_v_b_41')
// (2, 19, 'local_g2_4')
// (2, 19, 'lutff_3/in_3')
// (2, 19, 'sp4_v_b_28')
// (2, 20, 'neigh_op_top_2')
// (2, 20, 'sp4_v_b_17')
// (2, 21, 'local_g0_2')
// (2, 21, 'lutff_2/in_0')
// (2, 21, 'lutff_2/out')
// (2, 21, 'sp4_v_b_4')
// (2, 22, 'neigh_op_bot_2')
// (3, 20, 'neigh_op_tnl_2')
// (3, 21, 'neigh_op_lft_2')
// (3, 22, 'neigh_op_bnl_2')

wire n326;
// (1, 19, 'lutff_1/cout')
// (1, 19, 'lutff_2/in_3')

reg n327 = 0;
// (1, 19, 'neigh_op_tnr_0')
// (1, 20, 'neigh_op_rgt_0')
// (1, 21, 'neigh_op_bnr_0')
// (2, 19, 'local_g0_0')
// (2, 19, 'lutff_4/in_0')
// (2, 19, 'neigh_op_top_0')
// (2, 20, 'local_g1_0')
// (2, 20, 'lutff_0/in_3')
// (2, 20, 'lutff_0/out')
// (2, 21, 'neigh_op_bot_0')
// (3, 19, 'neigh_op_tnl_0')
// (3, 20, 'neigh_op_lft_0')
// (3, 21, 'neigh_op_bnl_0')

wire n328;
// (1, 19, 'neigh_op_tnr_2')
// (1, 20, 'neigh_op_rgt_2')
// (1, 21, 'neigh_op_bnr_2')
// (2, 19, 'neigh_op_top_2')
// (2, 20, 'local_g3_2')
// (2, 20, 'lutff_2/out')
// (2, 20, 'lutff_3/in_0')
// (2, 21, 'neigh_op_bot_2')
// (3, 19, 'neigh_op_tnl_2')
// (3, 20, 'neigh_op_lft_2')
// (3, 21, 'neigh_op_bnl_2')

reg n329 = 0;
// (1, 19, 'neigh_op_tnr_6')
// (1, 20, 'local_g2_6')
// (1, 20, 'local_g3_6')
// (1, 20, 'lutff_4/in_3')
// (1, 20, 'lutff_5/in_2')
// (1, 20, 'lutff_6/in_0')
// (1, 20, 'lutff_7/in_3')
// (1, 20, 'neigh_op_rgt_6')
// (1, 21, 'neigh_op_bnr_6')
// (2, 19, 'neigh_op_top_6')
// (2, 20, 'local_g1_6')
// (2, 20, 'lutff_6/in_1')
// (2, 20, 'lutff_6/out')
// (2, 21, 'neigh_op_bot_6')
// (3, 19, 'neigh_op_tnl_6')
// (3, 20, 'neigh_op_lft_6')
// (3, 21, 'neigh_op_bnl_6')

wire n330;
// (1, 19, 'neigh_op_tnr_7')
// (1, 20, 'neigh_op_rgt_7')
// (1, 21, 'neigh_op_bnr_7')
// (2, 19, 'neigh_op_top_7')
// (2, 20, 'lutff_7/out')
// (2, 21, 'neigh_op_bot_7')
// (3, 19, 'neigh_op_tnl_7')
// (3, 20, 'local_g0_7')
// (3, 20, 'lutff_1/in_0')
// (3, 20, 'neigh_op_lft_7')
// (3, 21, 'neigh_op_bnl_7')

reg n331 = 0;
// (1, 19, 'sp4_r_v_b_46')
// (1, 20, 'neigh_op_tnr_3')
// (1, 20, 'sp4_r_v_b_35')
// (1, 21, 'neigh_op_rgt_3')
// (1, 21, 'sp4_r_v_b_22')
// (1, 22, 'neigh_op_bnr_3')
// (1, 22, 'sp4_r_v_b_11')
// (2, 18, 'sp4_v_t_46')
// (2, 19, 'local_g3_6')
// (2, 19, 'lutff_3/in_0')
// (2, 19, 'sp4_v_b_46')
// (2, 20, 'neigh_op_top_3')
// (2, 20, 'sp4_v_b_35')
// (2, 21, 'local_g1_3')
// (2, 21, 'lutff_0/in_2')
// (2, 21, 'lutff_1/in_3')
// (2, 21, 'lutff_3/in_3')
// (2, 21, 'lutff_3/out')
// (2, 21, 'sp4_v_b_22')
// (2, 22, 'neigh_op_bot_3')
// (2, 22, 'sp4_v_b_11')
// (3, 20, 'neigh_op_tnl_3')
// (3, 21, 'neigh_op_lft_3')
// (3, 22, 'neigh_op_bnl_3')

wire n332;
// (1, 20, 'lutff_1/cout')
// (1, 20, 'lutff_2/in_3')

wire n333;
// (1, 20, 'neigh_op_tnr_6')
// (1, 21, 'neigh_op_rgt_6')
// (1, 22, 'neigh_op_bnr_6')
// (2, 20, 'neigh_op_top_6')
// (2, 21, 'lutff_6/out')
// (2, 22, 'neigh_op_bot_6')
// (3, 20, 'neigh_op_tnl_6')
// (3, 21, 'local_g0_6')
// (3, 21, 'lutff_0/in_0')
// (3, 21, 'lutff_2/in_0')
// (3, 21, 'neigh_op_lft_6')
// (3, 22, 'neigh_op_bnl_6')

reg n334 = 0;
// (1, 20, 'sp4_h_r_2')
// (2, 19, 'neigh_op_tnr_5')
// (2, 20, 'neigh_op_rgt_5')
// (2, 20, 'sp4_h_r_15')
// (2, 21, 'neigh_op_bnr_5')
// (3, 11, 'sp4_r_v_b_38')
// (3, 12, 'sp4_r_v_b_27')
// (3, 13, 'sp4_r_v_b_14')
// (3, 14, 'sp4_r_v_b_3')
// (3, 15, 'sp4_r_v_b_38')
// (3, 16, 'sp4_r_v_b_27')
// (3, 17, 'sp4_r_v_b_14')
// (3, 17, 'sp4_r_v_b_46')
// (3, 18, 'sp4_r_v_b_3')
// (3, 18, 'sp4_r_v_b_35')
// (3, 19, 'local_g1_5')
// (3, 19, 'lutff_3/in_1')
// (3, 19, 'neigh_op_top_5')
// (3, 19, 'sp4_r_v_b_22')
// (3, 19, 'sp4_r_v_b_38')
// (3, 20, 'lutff_5/out')
// (3, 20, 'sp4_h_r_10')
// (3, 20, 'sp4_h_r_26')
// (3, 20, 'sp4_r_v_b_11')
// (3, 20, 'sp4_r_v_b_27')
// (3, 21, 'neigh_op_bot_5')
// (3, 21, 'sp4_r_v_b_14')
// (3, 22, 'sp4_r_v_b_3')
// (4, 10, 'sp4_h_r_3')
// (4, 10, 'sp4_v_t_38')
// (4, 11, 'sp4_v_b_38')
// (4, 12, 'sp4_v_b_27')
// (4, 13, 'sp4_v_b_14')
// (4, 14, 'sp4_v_b_3')
// (4, 14, 'sp4_v_t_38')
// (4, 15, 'sp4_v_b_38')
// (4, 16, 'sp4_h_r_11')
// (4, 16, 'sp4_v_b_27')
// (4, 16, 'sp4_v_t_46')
// (4, 17, 'sp4_v_b_14')
// (4, 17, 'sp4_v_b_46')
// (4, 18, 'sp4_h_r_8')
// (4, 18, 'sp4_v_b_3')
// (4, 18, 'sp4_v_b_35')
// (4, 18, 'sp4_v_t_38')
// (4, 19, 'local_g3_5')
// (4, 19, 'lutff_1/in_1')
// (4, 19, 'neigh_op_tnl_5')
// (4, 19, 'sp4_v_b_22')
// (4, 19, 'sp4_v_b_38')
// (4, 20, 'neigh_op_lft_5')
// (4, 20, 'sp4_h_r_23')
// (4, 20, 'sp4_h_r_39')
// (4, 20, 'sp4_v_b_11')
// (4, 20, 'sp4_v_b_27')
// (4, 21, 'local_g2_5')
// (4, 21, 'lutff_7/in_2')
// (4, 21, 'neigh_op_bnl_5')
// (4, 21, 'sp4_v_b_14')
// (4, 22, 'sp4_v_b_3')
// (5, 10, 'sp4_h_r_14')
// (5, 16, 'sp4_h_r_22')
// (5, 18, 'sp4_h_r_21')
// (5, 20, 'sp4_h_l_39')
// (5, 20, 'sp4_h_r_10')
// (5, 20, 'sp4_h_r_34')
// (6, 10, 'sp4_h_r_27')
// (6, 16, 'sp4_h_r_35')
// (6, 18, 'sp4_h_r_32')
// (6, 20, 'sp4_h_r_23')
// (6, 20, 'sp4_h_r_47')
// (7, 10, 'sp4_h_r_38')
// (7, 16, 'local_g3_6')
// (7, 16, 'lutff_2/in_3')
// (7, 16, 'sp4_h_r_46')
// (7, 18, 'sp4_h_r_45')
// (7, 20, 'sp4_h_l_47')
// (7, 20, 'sp4_h_r_10')
// (7, 20, 'sp4_h_r_34')
// (8, 10, 'sp4_h_l_38')
// (8, 10, 'sp4_h_r_11')
// (8, 13, 'sp4_r_v_b_36')
// (8, 14, 'sp4_r_v_b_25')
// (8, 15, 'sp4_r_v_b_12')
// (8, 16, 'sp4_h_l_46')
// (8, 16, 'sp4_r_v_b_1')
// (8, 17, 'sp4_r_v_b_47')
// (8, 18, 'local_g1_3')
// (8, 18, 'lutff_4/in_2')
// (8, 18, 'sp4_h_l_45')
// (8, 18, 'sp4_h_r_11')
// (8, 18, 'sp4_r_v_b_34')
// (8, 19, 'sp4_r_v_b_23')
// (8, 20, 'sp4_h_r_23')
// (8, 20, 'sp4_h_r_47')
// (8, 20, 'sp4_r_v_b_10')
// (9, 10, 'sp4_h_r_22')
// (9, 12, 'sp4_v_t_36')
// (9, 13, 'sp4_v_b_36')
// (9, 14, 'sp4_v_b_25')
// (9, 15, 'local_g1_4')
// (9, 15, 'lutff_7/in_0')
// (9, 15, 'sp4_v_b_12')
// (9, 16, 'sp4_v_b_1')
// (9, 16, 'sp4_v_t_47')
// (9, 17, 'sp4_v_b_47')
// (9, 18, 'sp4_h_r_22')
// (9, 18, 'sp4_v_b_34')
// (9, 19, 'local_g0_7')
// (9, 19, 'lutff_6/in_1')
// (9, 19, 'sp4_v_b_23')
// (9, 20, 'sp4_h_l_47')
// (9, 20, 'sp4_h_r_34')
// (9, 20, 'sp4_v_b_10')
// (10, 10, 'local_g2_3')
// (10, 10, 'lutff_4/in_3')
// (10, 10, 'sp4_h_r_35')
// (10, 17, 'sp4_r_v_b_41')
// (10, 18, 'sp4_h_r_35')
// (10, 18, 'sp4_r_v_b_28')
// (10, 19, 'local_g3_1')
// (10, 19, 'lutff_4/in_2')
// (10, 19, 'sp4_r_v_b_17')
// (10, 20, 'sp4_h_r_47')
// (10, 20, 'sp4_r_v_b_4')
// (11, 10, 'sp4_h_r_46')
// (11, 16, 'sp4_v_t_41')
// (11, 17, 'sp4_v_b_41')
// (11, 18, 'sp4_h_r_46')
// (11, 18, 'sp4_v_b_28')
// (11, 19, 'sp4_v_b_17')
// (11, 20, 'sp4_h_l_47')
// (11, 20, 'sp4_v_b_4')
// (12, 10, 'sp4_h_l_46')
// (12, 18, 'sp4_h_l_46')

wire n335;
// (1, 21, 'local_g1_2')
// (1, 21, 'lutff_7/in_0')
// (1, 21, 'sp4_h_r_10')
// (2, 20, 'neigh_op_tnr_1')
// (2, 21, 'neigh_op_rgt_1')
// (2, 21, 'sp4_h_r_23')
// (2, 22, 'neigh_op_bnr_1')
// (3, 20, 'neigh_op_top_1')
// (3, 21, 'lutff_1/out')
// (3, 21, 'sp4_h_r_34')
// (3, 22, 'neigh_op_bot_1')
// (4, 20, 'neigh_op_tnl_1')
// (4, 21, 'neigh_op_lft_1')
// (4, 21, 'sp4_h_r_47')
// (4, 22, 'neigh_op_bnl_1')
// (5, 21, 'sp4_h_l_47')

wire n336;
// (1, 21, 'lutff_1/cout')
// (1, 21, 'lutff_2/in_3')

wire n337;
// (1, 21, 'lutff_2/cout')
// (1, 21, 'lutff_3/in_3')

wire n338;
// (2, 0, 'logic_op_tnr_0')
// (2, 1, 'neigh_op_rgt_0')
// (2, 2, 'neigh_op_bnr_0')
// (3, 0, 'logic_op_top_0')
// (3, 1, 'local_g3_0')
// (3, 1, 'lutff_0/out')
// (3, 1, 'lutff_3/in_2')
// (3, 2, 'neigh_op_bot_0')
// (4, 0, 'logic_op_tnl_0')
// (4, 1, 'neigh_op_lft_0')
// (4, 2, 'neigh_op_bnl_0')

reg n339 = 0;
// (2, 0, 'logic_op_tnr_1')
// (2, 1, 'neigh_op_rgt_1')
// (2, 2, 'neigh_op_bnr_1')
// (3, 0, 'logic_op_top_1')
// (3, 1, 'local_g1_1')
// (3, 1, 'lutff_1/out')
// (3, 1, 'lutff_2/in_0')
// (3, 2, 'neigh_op_bot_1')
// (4, 0, 'logic_op_tnl_1')
// (4, 1, 'neigh_op_lft_1')
// (4, 2, 'neigh_op_bnl_1')

wire n340;
// (2, 0, 'logic_op_tnr_2')
// (2, 1, 'neigh_op_rgt_2')
// (2, 2, 'neigh_op_bnr_2')
// (3, 0, 'logic_op_top_2')
// (3, 1, 'local_g3_2')
// (3, 1, 'lutff_2/out')
// (3, 1, 'lutff_3/in_0')
// (3, 2, 'neigh_op_bot_2')
// (4, 0, 'logic_op_tnl_2')
// (4, 1, 'neigh_op_lft_2')
// (4, 2, 'neigh_op_bnl_2')

wire n341;
// (2, 0, 'logic_op_tnr_3')
// (2, 1, 'neigh_op_rgt_3')
// (2, 2, 'neigh_op_bnr_3')
// (3, 0, 'logic_op_top_3')
// (3, 1, 'lutff_3/out')
// (3, 2, 'local_g0_3')
// (3, 2, 'lutff_6/in_1')
// (3, 2, 'neigh_op_bot_3')
// (4, 0, 'logic_op_tnl_3')
// (4, 1, 'neigh_op_lft_3')
// (4, 2, 'neigh_op_bnl_3')

reg n342 = 0;
// (2, 0, 'logic_op_tnr_4')
// (2, 1, 'neigh_op_rgt_4')
// (2, 2, 'neigh_op_bnr_4')
// (3, 0, 'logic_op_top_4')
// (3, 1, 'local_g2_4')
// (3, 1, 'lutff_0/in_2')
// (3, 1, 'lutff_4/out')
// (3, 2, 'neigh_op_bot_4')
// (4, 0, 'logic_op_tnl_4')
// (4, 1, 'neigh_op_lft_4')
// (4, 2, 'neigh_op_bnl_4')

reg n343 = 0;
// (2, 0, 'logic_op_tnr_5')
// (2, 1, 'neigh_op_rgt_5')
// (2, 2, 'neigh_op_bnr_5')
// (3, 0, 'logic_op_top_5')
// (3, 1, 'local_g0_5')
// (3, 1, 'lutff_0/in_3')
// (3, 1, 'lutff_5/out')
// (3, 2, 'neigh_op_bot_5')
// (4, 0, 'logic_op_tnl_5')
// (4, 1, 'neigh_op_lft_5')
// (4, 2, 'neigh_op_bnl_5')

reg n344 = 0;
// (2, 0, 'logic_op_tnr_6')
// (2, 1, 'neigh_op_rgt_6')
// (2, 2, 'neigh_op_bnr_6')
// (3, 0, 'logic_op_top_6')
// (3, 1, 'lutff_6/out')
// (3, 2, 'local_g1_6')
// (3, 2, 'lutff_2/in_1')
// (3, 2, 'neigh_op_bot_6')
// (4, 0, 'logic_op_tnl_6')
// (4, 1, 'neigh_op_lft_6')
// (4, 2, 'neigh_op_bnl_6')

reg n345 = 0;
// (2, 0, 'logic_op_tnr_7')
// (2, 1, 'neigh_op_rgt_7')
// (2, 2, 'neigh_op_bnr_7')
// (3, 0, 'logic_op_top_7')
// (3, 1, 'local_g2_7')
// (3, 1, 'lutff_2/in_3')
// (3, 1, 'lutff_7/out')
// (3, 2, 'neigh_op_bot_7')
// (4, 0, 'logic_op_tnl_7')
// (4, 1, 'neigh_op_lft_7')
// (4, 2, 'neigh_op_bnl_7')

wire n346;
// (2, 1, 'neigh_op_tnr_0')
// (2, 2, 'neigh_op_rgt_0')
// (2, 3, 'neigh_op_bnr_0')
// (3, 1, 'neigh_op_top_0')
// (3, 2, 'local_g2_0')
// (3, 2, 'lutff_0/out')
// (3, 2, 'lutff_7/in_3')
// (3, 3, 'neigh_op_bot_0')
// (4, 1, 'neigh_op_tnl_0')
// (4, 2, 'neigh_op_lft_0')
// (4, 3, 'neigh_op_bnl_0')

reg n347 = 0;
// (2, 1, 'neigh_op_tnr_1')
// (2, 2, 'neigh_op_rgt_1')
// (2, 3, 'neigh_op_bnr_1')
// (3, 1, 'neigh_op_top_1')
// (3, 2, 'local_g2_1')
// (3, 2, 'lutff_1/out')
// (3, 2, 'lutff_4/in_3')
// (3, 3, 'neigh_op_bot_1')
// (4, 1, 'neigh_op_tnl_1')
// (4, 2, 'neigh_op_lft_1')
// (4, 3, 'neigh_op_bnl_1')

wire n348;
// (2, 1, 'neigh_op_tnr_2')
// (2, 2, 'neigh_op_rgt_2')
// (2, 3, 'neigh_op_bnr_2')
// (3, 1, 'neigh_op_top_2')
// (3, 2, 'local_g2_2')
// (3, 2, 'lutff_2/out')
// (3, 2, 'lutff_6/in_0')
// (3, 3, 'neigh_op_bot_2')
// (4, 1, 'neigh_op_tnl_2')
// (4, 2, 'neigh_op_lft_2')
// (4, 3, 'neigh_op_bnl_2')

reg n349 = 0;
// (2, 1, 'neigh_op_tnr_3')
// (2, 2, 'neigh_op_rgt_3')
// (2, 3, 'neigh_op_bnr_3')
// (3, 1, 'neigh_op_top_3')
// (3, 2, 'local_g2_3')
// (3, 2, 'lutff_3/out')
// (3, 2, 'lutff_4/in_1')
// (3, 3, 'neigh_op_bot_3')
// (4, 1, 'neigh_op_tnl_3')
// (4, 2, 'neigh_op_lft_3')
// (4, 3, 'neigh_op_bnl_3')

wire n350;
// (2, 1, 'neigh_op_tnr_4')
// (2, 2, 'neigh_op_rgt_4')
// (2, 3, 'neigh_op_bnr_4')
// (3, 1, 'neigh_op_top_4')
// (3, 2, 'local_g2_4')
// (3, 2, 'lutff_4/out')
// (3, 2, 'lutff_6/in_2')
// (3, 3, 'neigh_op_bot_4')
// (4, 1, 'neigh_op_tnl_4')
// (4, 2, 'neigh_op_lft_4')
// (4, 3, 'neigh_op_bnl_4')

reg n351 = 0;
// (2, 1, 'neigh_op_tnr_5')
// (2, 2, 'neigh_op_rgt_5')
// (2, 3, 'neigh_op_bnr_5')
// (3, 1, 'neigh_op_top_5')
// (3, 2, 'local_g2_5')
// (3, 2, 'lutff_2/in_3')
// (3, 2, 'lutff_5/out')
// (3, 3, 'neigh_op_bot_5')
// (4, 1, 'neigh_op_tnl_5')
// (4, 2, 'neigh_op_lft_5')
// (4, 3, 'neigh_op_bnl_5')

wire n352;
// (2, 1, 'neigh_op_tnr_6')
// (2, 2, 'neigh_op_rgt_6')
// (2, 3, 'neigh_op_bnr_6')
// (3, 1, 'neigh_op_top_6')
// (3, 2, 'local_g2_6')
// (3, 2, 'lutff_6/out')
// (3, 2, 'lutff_7/in_1')
// (3, 3, 'neigh_op_bot_6')
// (4, 1, 'neigh_op_tnl_6')
// (4, 2, 'neigh_op_lft_6')
// (4, 3, 'neigh_op_bnl_6')

wire n353;
// (2, 1, 'neigh_op_tnr_7')
// (2, 2, 'neigh_op_rgt_7')
// (2, 3, 'neigh_op_bnr_7')
// (3, 1, 'neigh_op_top_7')
// (3, 2, 'lutff_7/out')
// (3, 3, 'neigh_op_bot_7')
// (4, 1, 'neigh_op_tnl_7')
// (4, 2, 'local_g1_7')
// (4, 2, 'lutff_7/in_3')
// (4, 2, 'neigh_op_lft_7')
// (4, 3, 'neigh_op_bnl_7')

reg n354 = 0;
// (2, 2, 'local_g1_5')
// (2, 2, 'lutff_6/in_0')
// (2, 2, 'sp4_h_r_5')
// (2, 7, 'sp4_h_r_2')
// (3, 1, 'sp4_r_v_b_13')
// (3, 1, 'sp4_r_v_b_20')
// (3, 2, 'local_g1_0')
// (3, 2, 'lutff_5/in_2')
// (3, 2, 'sp4_h_r_16')
// (3, 2, 'sp4_r_v_b_0')
// (3, 2, 'sp4_r_v_b_9')
// (3, 3, 'local_g3_4')
// (3, 3, 'lutff_0/in_3')
// (3, 3, 'sp4_r_v_b_44')
// (3, 3, 'sp4_r_v_b_46')
// (3, 4, 'sp4_r_v_b_33')
// (3, 4, 'sp4_r_v_b_35')
// (3, 5, 'sp4_r_v_b_20')
// (3, 5, 'sp4_r_v_b_22')
// (3, 6, 'sp4_r_v_b_11')
// (3, 6, 'sp4_r_v_b_9')
// (3, 7, 'local_g0_7')
// (3, 7, 'lutff_5/in_2')
// (3, 7, 'sp4_h_r_15')
// (3, 7, 'sp4_r_v_b_44')
// (3, 8, 'sp4_r_v_b_33')
// (3, 9, 'sp4_r_v_b_20')
// (3, 10, 'local_g2_1')
// (3, 10, 'lutff_1/in_2')
// (3, 10, 'sp4_r_v_b_9')
// (4, 0, 'span4_vert_13')
// (4, 0, 'span4_vert_20')
// (4, 1, 'local_g1_4')
// (4, 1, 'lutff_0/in_1')
// (4, 1, 'sp4_v_b_13')
// (4, 1, 'sp4_v_b_20')
// (4, 2, 'sp4_h_r_29')
// (4, 2, 'sp4_v_b_0')
// (4, 2, 'sp4_v_b_9')
// (4, 2, 'sp4_v_t_44')
// (4, 2, 'sp4_v_t_46')
// (4, 3, 'local_g3_6')
// (4, 3, 'lutff_6/in_3')
// (4, 3, 'sp4_v_b_44')
// (4, 3, 'sp4_v_b_46')
// (4, 4, 'sp4_v_b_33')
// (4, 4, 'sp4_v_b_35')
// (4, 5, 'local_g1_4')
// (4, 5, 'lutff_1/in_2')
// (4, 5, 'sp4_v_b_20')
// (4, 5, 'sp4_v_b_22')
// (4, 6, 'sp4_h_r_6')
// (4, 6, 'sp4_h_r_9')
// (4, 6, 'sp4_v_b_11')
// (4, 6, 'sp4_v_b_9')
// (4, 6, 'sp4_v_t_44')
// (4, 7, 'sp4_h_r_26')
// (4, 7, 'sp4_v_b_44')
// (4, 8, 'sp4_v_b_33')
// (4, 9, 'sp4_v_b_20')
// (4, 10, 'sp4_v_b_9')
// (5, 2, 'sp4_h_r_40')
// (5, 4, 'sp4_r_v_b_46')
// (5, 5, 'sp4_r_v_b_35')
// (5, 6, 'sp4_h_r_19')
// (5, 6, 'sp4_h_r_20')
// (5, 6, 'sp4_r_v_b_22')
// (5, 7, 'local_g2_3')
// (5, 7, 'lutff_1/in_2')
// (5, 7, 'sp4_h_r_39')
// (5, 7, 'sp4_r_v_b_11')
// (5, 17, 'sp4_r_v_b_44')
// (5, 18, 'sp4_r_v_b_33')
// (5, 19, 'sp4_r_v_b_20')
// (5, 20, 'local_g2_1')
// (5, 20, 'lutff_5/in_2')
// (5, 20, 'sp4_r_v_b_9')
// (6, 2, 'sp4_h_l_40')
// (6, 2, 'sp4_h_r_2')
// (6, 3, 'sp4_v_t_46')
// (6, 4, 'sp4_v_b_46')
// (6, 5, 'sp4_v_b_35')
// (6, 6, 'sp4_h_r_30')
// (6, 6, 'sp4_h_r_33')
// (6, 6, 'sp4_v_b_22')
// (6, 7, 'sp4_h_l_39')
// (6, 7, 'sp4_h_r_6')
// (6, 7, 'sp4_v_b_11')
// (6, 16, 'sp4_h_r_3')
// (6, 16, 'sp4_v_t_44')
// (6, 17, 'sp4_v_b_44')
// (6, 18, 'sp4_v_b_33')
// (6, 19, 'sp4_v_b_20')
// (6, 20, 'sp4_v_b_9')
// (7, 2, 'sp4_h_r_15')
// (7, 3, 'sp4_r_v_b_43')
// (7, 4, 'sp4_r_v_b_30')
// (7, 5, 'sp4_r_v_b_19')
// (7, 6, 'sp4_h_r_43')
// (7, 6, 'sp4_h_r_44')
// (7, 6, 'sp4_r_v_b_6')
// (7, 7, 'sp4_h_r_19')
// (7, 7, 'sp4_r_v_b_37')
// (7, 8, 'sp4_r_v_b_24')
// (7, 9, 'sp4_r_v_b_13')
// (7, 10, 'sp4_r_v_b_0')
// (7, 11, 'sp4_r_v_b_37')
// (7, 11, 'sp4_r_v_b_46')
// (7, 12, 'sp4_r_v_b_24')
// (7, 12, 'sp4_r_v_b_35')
// (7, 13, 'sp4_r_v_b_13')
// (7, 13, 'sp4_r_v_b_22')
// (7, 14, 'sp4_r_v_b_0')
// (7, 14, 'sp4_r_v_b_11')
// (7, 15, 'sp4_r_v_b_46')
// (7, 16, 'sp4_h_r_14')
// (7, 16, 'sp4_r_v_b_35')
// (7, 17, 'sp4_r_v_b_22')
// (7, 18, 'sp4_r_v_b_11')
// (7, 19, 'sp4_r_v_b_42')
// (7, 20, 'sp4_r_v_b_31')
// (7, 21, 'local_g3_2')
// (7, 21, 'lutff_6/in_1')
// (7, 21, 'sp4_r_v_b_18')
// (7, 22, 'sp4_r_v_b_7')
// (8, 2, 'sp4_h_r_26')
// (8, 2, 'sp4_v_t_43')
// (8, 3, 'sp4_r_v_b_42')
// (8, 3, 'sp4_v_b_43')
// (8, 4, 'sp4_r_v_b_31')
// (8, 4, 'sp4_v_b_30')
// (8, 5, 'local_g0_3')
// (8, 5, 'lutff_1/in_2')
// (8, 5, 'sp4_r_v_b_18')
// (8, 5, 'sp4_v_b_19')
// (8, 6, 'sp4_h_l_43')
// (8, 6, 'sp4_h_l_44')
// (8, 6, 'sp4_h_r_6')
// (8, 6, 'sp4_r_v_b_7')
// (8, 6, 'sp4_v_b_6')
// (8, 6, 'sp4_v_t_37')
// (8, 7, 'sp4_h_r_30')
// (8, 7, 'sp4_v_b_37')
// (8, 8, 'local_g3_0')
// (8, 8, 'lutff_4/in_1')
// (8, 8, 'sp4_v_b_24')
// (8, 9, 'sp4_v_b_13')
// (8, 10, 'sp4_h_r_5')
// (8, 10, 'sp4_v_b_0')
// (8, 10, 'sp4_v_t_37')
// (8, 10, 'sp4_v_t_46')
// (8, 11, 'sp4_v_b_37')
// (8, 11, 'sp4_v_b_46')
// (8, 12, 'sp4_v_b_24')
// (8, 12, 'sp4_v_b_35')
// (8, 13, 'local_g0_5')
// (8, 13, 'lutff_0/in_3')
// (8, 13, 'sp4_v_b_13')
// (8, 13, 'sp4_v_b_22')
// (8, 14, 'sp4_h_r_9')
// (8, 14, 'sp4_v_b_0')
// (8, 14, 'sp4_v_b_11')
// (8, 14, 'sp4_v_t_46')
// (8, 15, 'sp4_v_b_46')
// (8, 16, 'sp4_h_r_27')
// (8, 16, 'sp4_v_b_35')
// (8, 17, 'sp4_v_b_22')
// (8, 18, 'sp4_v_b_11')
// (8, 18, 'sp4_v_t_42')
// (8, 19, 'sp4_v_b_42')
// (8, 20, 'sp4_v_b_31')
// (8, 21, 'sp4_v_b_18')
// (8, 22, 'sp4_v_b_7')
// (9, 1, 'local_g3_5')
// (9, 1, 'lutff_3/in_3')
// (9, 1, 'sp4_r_v_b_21')
// (9, 2, 'sp4_h_r_39')
// (9, 2, 'sp4_r_v_b_8')
// (9, 2, 'sp4_v_t_42')
// (9, 3, 'sp4_v_b_42')
// (9, 4, 'sp4_v_b_31')
// (9, 5, 'local_g1_2')
// (9, 5, 'lutff_3/in_0')
// (9, 5, 'sp4_v_b_18')
// (9, 6, 'sp4_h_r_19')
// (9, 6, 'sp4_h_r_2')
// (9, 6, 'sp4_v_b_7')
// (9, 7, 'sp4_h_r_43')
// (9, 10, 'sp4_h_r_16')
// (9, 14, 'local_g1_4')
// (9, 14, 'lutff_5/in_2')
// (9, 14, 'sp4_h_r_20')
// (9, 16, 'sp4_h_r_38')
// (10, 0, 'span4_vert_21')
// (10, 1, 'sp4_v_b_21')
// (10, 2, 'sp4_h_l_39')
// (10, 2, 'sp4_h_r_11')
// (10, 2, 'sp4_h_r_8')
// (10, 2, 'sp4_v_b_8')
// (10, 3, 'sp4_h_r_4')
// (10, 6, 'sp4_h_r_15')
// (10, 6, 'sp4_h_r_3')
// (10, 6, 'sp4_h_r_30')
// (10, 7, 'sp12_h_r_1')
// (10, 7, 'sp12_v_t_22')
// (10, 7, 'sp4_h_l_43')
// (10, 7, 'sp4_h_r_3')
// (10, 8, 'sp12_v_b_22')
// (10, 9, 'sp12_v_b_21')
// (10, 10, 'sp12_v_b_18')
// (10, 10, 'sp4_h_r_29')
// (10, 11, 'sp12_v_b_17')
// (10, 12, 'sp12_v_b_14')
// (10, 13, 'sp12_v_b_13')
// (10, 14, 'sp12_v_b_10')
// (10, 14, 'sp4_h_r_33')
// (10, 15, 'sp12_h_r_1')
// (10, 15, 'sp12_v_b_9')
// (10, 15, 'sp12_v_t_22')
// (10, 16, 'sp12_v_b_22')
// (10, 16, 'sp12_v_b_6')
// (10, 16, 'sp4_h_l_38')
// (10, 16, 'sp4_h_r_0')
// (10, 17, 'local_g2_5')
// (10, 17, 'lutff_7/in_0')
// (10, 17, 'sp12_v_b_21')
// (10, 17, 'sp12_v_b_5')
// (10, 18, 'local_g3_2')
// (10, 18, 'lutff_4/in_1')
// (10, 18, 'sp12_v_b_18')
// (10, 18, 'sp12_v_b_2')
// (10, 19, 'sp12_v_b_1')
// (10, 19, 'sp12_v_b_17')
// (10, 20, 'local_g3_6')
// (10, 20, 'lutff_1/in_2')
// (10, 20, 'lutff_5/in_0')
// (10, 20, 'sp12_v_b_14')
// (10, 21, 'sp12_v_b_13')
// (10, 22, 'sp12_v_b_10')
// (10, 23, 'sp12_v_b_9')
// (10, 24, 'sp12_v_b_6')
// (10, 25, 'sp12_v_b_5')
// (10, 26, 'sp12_v_b_2')
// (10, 27, 'sp12_v_b_1')
// (11, 2, 'local_g0_6')
// (11, 2, 'lutff_1/in_1')
// (11, 2, 'sp4_h_r_21')
// (11, 2, 'sp4_h_r_22')
// (11, 3, 'local_g0_1')
// (11, 3, 'lutff_7/in_2')
// (11, 3, 'sp4_h_r_17')
// (11, 6, 'local_g0_6')
// (11, 6, 'lutff_3/in_1')
// (11, 6, 'sp4_h_r_14')
// (11, 6, 'sp4_h_r_26')
// (11, 6, 'sp4_h_r_43')
// (11, 7, 'sp12_h_r_2')
// (11, 7, 'sp4_h_r_14')
// (11, 7, 'sp4_h_r_2')
// (11, 7, 'sp4_r_v_b_42')
// (11, 8, 'sp4_r_v_b_31')
// (11, 9, 'sp4_r_v_b_18')
// (11, 10, 'sp4_h_r_40')
// (11, 10, 'sp4_r_v_b_7')
// (11, 11, 'sp4_r_v_b_44')
// (11, 12, 'sp4_r_v_b_33')
// (11, 13, 'sp4_r_v_b_20')
// (11, 14, 'sp4_h_r_44')
// (11, 14, 'sp4_r_v_b_9')
// (11, 15, 'sp12_h_r_2')
// (11, 16, 'sp4_h_r_13')
// (12, 2, 'sp4_h_r_32')
// (12, 2, 'sp4_h_r_35')
// (12, 3, 'sp4_h_r_28')
// (12, 6, 'sp4_h_l_43')
// (12, 6, 'sp4_h_r_1')
// (12, 6, 'sp4_h_r_27')
// (12, 6, 'sp4_h_r_39')
// (12, 6, 'sp4_h_r_6')
// (12, 6, 'sp4_v_t_42')
// (12, 7, 'local_g1_7')
// (12, 7, 'lutff_3/in_3')
// (12, 7, 'sp12_h_r_5')
// (12, 7, 'sp4_h_r_15')
// (12, 7, 'sp4_h_r_27')
// (12, 7, 'sp4_v_b_42')
// (12, 8, 'local_g2_7')
// (12, 8, 'lutff_6/in_1')
// (12, 8, 'sp4_v_b_31')
// (12, 9, 'sp4_v_b_18')
// (12, 10, 'sp4_h_l_40')
// (12, 10, 'sp4_h_r_9')
// (12, 10, 'sp4_v_b_7')
// (12, 10, 'sp4_v_t_44')
// (12, 11, 'sp4_v_b_44')
// (12, 12, 'sp4_v_b_33')
// (12, 13, 'sp4_v_b_20')
// (12, 14, 'sp4_h_l_44')
// (12, 14, 'sp4_v_b_9')
// (12, 15, 'sp12_h_r_5')
// (12, 16, 'sp4_h_r_24')
// (13, 2, 'sp4_h_r_45')
// (13, 2, 'sp4_h_r_46')
// (13, 3, 'sp4_h_r_41')
// (13, 3, 'sp4_r_v_b_37')
// (13, 4, 'sp4_r_v_b_24')
// (13, 5, 'sp4_r_v_b_13')
// (13, 6, 'sp4_h_l_39')
// (13, 6, 'sp4_h_r_11')
// (13, 6, 'sp4_h_r_12')
// (13, 6, 'sp4_h_r_19')
// (13, 6, 'sp4_h_r_38')
// (13, 6, 'sp4_r_v_b_0')
// (13, 7, 'sp12_h_r_6')
// (13, 7, 'sp4_h_r_26')
// (13, 7, 'sp4_h_r_38')
// (13, 10, 'sp4_h_r_20')
// (13, 15, 'sp12_h_r_6')
// (13, 16, 'sp4_h_r_37')
// (14, 2, 'sp4_h_l_45')
// (14, 2, 'sp4_h_l_46')
// (14, 2, 'sp4_h_r_8')
// (14, 2, 'sp4_v_t_37')
// (14, 3, 'local_g0_4')
// (14, 3, 'lutff_3/in_3')
// (14, 3, 'sp4_h_l_41')
// (14, 3, 'sp4_h_r_4')
// (14, 3, 'sp4_v_b_37')
// (14, 4, 'sp4_v_b_24')
// (14, 5, 'local_g1_5')
// (14, 5, 'lutff_0/in_2')
// (14, 5, 'sp4_v_b_13')
// (14, 6, 'sp4_h_l_38')
// (14, 6, 'sp4_h_r_22')
// (14, 6, 'sp4_h_r_25')
// (14, 6, 'sp4_h_r_30')
// (14, 6, 'sp4_h_r_7')
// (14, 6, 'sp4_v_b_0')
// (14, 7, 'sp12_h_r_9')
// (14, 7, 'sp4_h_l_38')
// (14, 7, 'sp4_h_r_0')
// (14, 7, 'sp4_h_r_39')
// (14, 10, 'sp4_h_r_33')
// (14, 15, 'sp12_h_r_9')
// (14, 16, 'sp4_h_l_37')
// (14, 16, 'sp4_h_r_9')
// (15, 2, 'sp4_h_r_21')
// (15, 3, 'sp4_h_r_17')
// (15, 3, 'sp4_r_v_b_47')
// (15, 4, 'local_g0_1')
// (15, 4, 'lutff_2/in_1')
// (15, 4, 'sp4_r_v_b_34')
// (15, 5, 'local_g3_7')
// (15, 5, 'lutff_3/in_1')
// (15, 5, 'sp4_r_v_b_23')
// (15, 6, 'sp4_h_r_18')
// (15, 6, 'sp4_h_r_35')
// (15, 6, 'sp4_h_r_36')
// (15, 6, 'sp4_h_r_43')
// (15, 6, 'sp4_r_v_b_10')
// (15, 7, 'sp12_h_r_10')
// (15, 7, 'sp4_h_l_39')
// (15, 7, 'sp4_h_r_13')
// (15, 7, 'sp4_h_r_6')
// (15, 7, 'sp4_r_v_b_41')
// (15, 8, 'sp4_r_v_b_28')
// (15, 9, 'sp4_r_v_b_17')
// (15, 10, 'sp4_h_r_44')
// (15, 10, 'sp4_r_v_b_4')
// (15, 15, 'sp12_h_r_10')
// (15, 16, 'sp4_h_r_20')
// (16, 2, 'local_g2_0')
// (16, 2, 'lutff_5/in_1')
// (16, 2, 'sp4_h_r_32')
// (16, 2, 'sp4_v_t_47')
// (16, 3, 'sp4_h_r_28')
// (16, 3, 'sp4_v_b_47')
// (16, 4, 'sp4_v_b_34')
// (16, 5, 'sp4_v_b_23')
// (16, 6, 'sp4_h_l_36')
// (16, 6, 'sp4_h_l_43')
// (16, 6, 'sp4_h_r_10')
// (16, 6, 'sp4_h_r_31')
// (16, 6, 'sp4_h_r_46')
// (16, 6, 'sp4_v_b_10')
// (16, 6, 'sp4_v_t_41')
// (16, 7, 'sp12_h_r_13')
// (16, 7, 'sp4_h_r_19')
// (16, 7, 'sp4_h_r_24')
// (16, 7, 'sp4_v_b_41')
// (16, 8, 'sp4_v_b_28')
// (16, 9, 'sp4_v_b_17')
// (16, 10, 'sp4_h_l_44')
// (16, 10, 'sp4_v_b_4')
// (16, 15, 'sp12_h_r_13')
// (16, 16, 'sp4_h_r_33')
// (17, 2, 'sp4_h_r_45')
// (17, 3, 'sp4_h_r_41')
// (17, 6, 'sp4_h_l_46')
// (17, 6, 'sp4_h_r_23')
// (17, 6, 'sp4_h_r_3')
// (17, 6, 'sp4_h_r_42')
// (17, 7, 'sp12_h_r_14')
// (17, 7, 'sp4_h_r_30')
// (17, 7, 'sp4_h_r_37')
// (17, 15, 'sp12_h_r_14')
// (17, 16, 'sp4_h_r_44')
// (18, 2, 'sp4_h_l_45')
// (18, 2, 'sp4_h_r_8')
// (18, 3, 'sp4_h_l_41')
// (18, 3, 'sp4_h_r_1')
// (18, 6, 'sp4_h_l_42')
// (18, 6, 'sp4_h_r_14')
// (18, 6, 'sp4_h_r_34')
// (18, 6, 'sp4_h_r_7')
// (18, 7, 'sp12_h_r_17')
// (18, 7, 'sp4_h_l_37')
// (18, 7, 'sp4_h_r_0')
// (18, 7, 'sp4_h_r_43')
// (18, 15, 'sp12_h_r_17')
// (18, 16, 'sp4_h_l_44')
// (18, 16, 'sp4_h_r_6')
// (19, 2, 'sp4_h_r_21')
// (19, 3, 'sp4_h_r_12')
// (19, 6, 'sp4_h_r_18')
// (19, 6, 'sp4_h_r_27')
// (19, 6, 'sp4_h_r_47')
// (19, 7, 'sp12_h_r_18')
// (19, 7, 'sp4_h_l_43')
// (19, 7, 'sp4_h_r_13')
// (19, 7, 'sp4_h_r_6')
// (19, 15, 'sp12_h_r_18')
// (19, 16, 'sp4_h_r_19')
// (20, 2, 'sp4_h_r_32')
// (20, 3, 'sp4_h_r_25')
// (20, 6, 'sp4_h_l_47')
// (20, 6, 'sp4_h_r_10')
// (20, 6, 'sp4_h_r_31')
// (20, 6, 'sp4_h_r_38')
// (20, 7, 'sp12_h_r_21')
// (20, 7, 'sp4_h_r_19')
// (20, 7, 'sp4_h_r_24')
// (20, 15, 'sp12_h_r_21')
// (20, 16, 'sp4_h_r_30')
// (21, 2, 'sp4_h_r_45')
// (21, 3, 'sp4_h_r_36')
// (21, 3, 'sp4_r_v_b_39')
// (21, 4, 'sp4_r_v_b_26')
// (21, 4, 'sp4_r_v_b_42')
// (21, 5, 'neigh_op_tnr_1')
// (21, 5, 'sp4_r_v_b_15')
// (21, 5, 'sp4_r_v_b_31')
// (21, 6, 'neigh_op_rgt_1')
// (21, 6, 'sp4_h_l_38')
// (21, 6, 'sp4_h_r_23')
// (21, 6, 'sp4_h_r_42')
// (21, 6, 'sp4_h_r_7')
// (21, 6, 'sp4_r_v_b_18')
// (21, 6, 'sp4_r_v_b_2')
// (21, 7, 'neigh_op_bnr_1')
// (21, 7, 'sp12_h_r_22')
// (21, 7, 'sp4_h_r_30')
// (21, 7, 'sp4_h_r_37')
// (21, 7, 'sp4_r_v_b_7')
// (21, 13, 'sp4_r_v_b_36')
// (21, 14, 'sp4_r_v_b_25')
// (21, 15, 'sp12_h_r_22')
// (21, 15, 'sp4_r_v_b_12')
// (21, 16, 'sp4_h_r_43')
// (21, 16, 'sp4_r_v_b_1')
// (22, 0, 'span12_vert_13')
// (22, 1, 'sp12_v_b_13')
// (22, 2, 'sp12_v_b_10')
// (22, 2, 'sp4_h_l_45')
// (22, 2, 'sp4_v_t_39')
// (22, 3, 'sp12_v_b_9')
// (22, 3, 'sp12_v_t_22')
// (22, 3, 'sp4_h_l_36')
// (22, 3, 'sp4_v_b_39')
// (22, 3, 'sp4_v_t_42')
// (22, 4, 'sp12_v_b_22')
// (22, 4, 'sp12_v_b_6')
// (22, 4, 'sp4_r_v_b_43')
// (22, 4, 'sp4_v_b_26')
// (22, 4, 'sp4_v_b_42')
// (22, 5, 'neigh_op_top_1')
// (22, 5, 'sp12_v_b_21')
// (22, 5, 'sp12_v_b_5')
// (22, 5, 'sp4_r_v_b_30')
// (22, 5, 'sp4_v_b_15')
// (22, 5, 'sp4_v_b_31')
// (22, 6, 'lutff_1/out')
// (22, 6, 'sp12_v_b_18')
// (22, 6, 'sp12_v_b_2')
// (22, 6, 'sp4_h_l_42')
// (22, 6, 'sp4_h_r_18')
// (22, 6, 'sp4_h_r_34')
// (22, 6, 'sp4_r_v_b_19')
// (22, 6, 'sp4_v_b_18')
// (22, 6, 'sp4_v_b_2')
// (22, 7, 'neigh_op_bot_1')
// (22, 7, 'sp12_h_l_22')
// (22, 7, 'sp12_v_b_1')
// (22, 7, 'sp12_v_b_17')
// (22, 7, 'sp4_h_l_37')
// (22, 7, 'sp4_h_r_43')
// (22, 7, 'sp4_r_v_b_6')
// (22, 7, 'sp4_v_b_7')
// (22, 8, 'sp12_v_b_14')
// (22, 9, 'sp12_v_b_13')
// (22, 10, 'sp12_v_b_10')
// (22, 11, 'sp12_v_b_9')
// (22, 12, 'sp12_v_b_6')
// (22, 12, 'sp4_v_t_36')
// (22, 13, 'sp12_v_b_5')
// (22, 13, 'sp4_v_b_36')
// (22, 14, 'sp12_v_b_2')
// (22, 14, 'sp4_v_b_25')
// (22, 15, 'sp12_h_l_22')
// (22, 15, 'sp12_v_b_1')
// (22, 15, 'sp4_v_b_12')
// (22, 16, 'sp4_h_l_43')
// (22, 16, 'sp4_v_b_1')
// (23, 3, 'sp4_v_t_43')
// (23, 4, 'sp4_v_b_43')
// (23, 5, 'neigh_op_tnl_1')
// (23, 5, 'sp4_v_b_30')
// (23, 6, 'neigh_op_lft_1')
// (23, 6, 'sp4_h_r_31')
// (23, 6, 'sp4_h_r_47')
// (23, 6, 'sp4_v_b_19')
// (23, 7, 'neigh_op_bnl_1')
// (23, 7, 'sp4_h_l_43')
// (23, 7, 'sp4_v_b_6')
// (24, 6, 'sp4_h_l_47')
// (24, 6, 'sp4_h_r_42')
// (25, 6, 'sp4_h_l_42')

reg n355 = 0;
// (2, 2, 'neigh_op_tnr_0')
// (2, 3, 'neigh_op_rgt_0')
// (2, 3, 'sp4_h_r_5')
// (2, 4, 'neigh_op_bnr_0')
// (3, 2, 'neigh_op_top_0')
// (3, 3, 'local_g1_0')
// (3, 3, 'lutff_0/out')
// (3, 3, 'lutff_3/in_0')
// (3, 3, 'sp4_h_r_16')
// (3, 4, 'neigh_op_bot_0')
// (4, 2, 'neigh_op_tnl_0')
// (4, 3, 'neigh_op_lft_0')
// (4, 3, 'sp4_h_r_29')
// (4, 4, 'neigh_op_bnl_0')
// (5, 1, 'sp4_r_v_b_29')
// (5, 2, 'local_g3_0')
// (5, 2, 'lutff_0/in_3')
// (5, 2, 'sp4_r_v_b_16')
// (5, 3, 'local_g1_5')
// (5, 3, 'lutff_7/in_1')
// (5, 3, 'sp4_h_r_40')
// (5, 3, 'sp4_r_v_b_5')
// (6, 0, 'span4_vert_29')
// (6, 1, 'sp4_v_b_29')
// (6, 2, 'sp4_v_b_16')
// (6, 3, 'sp4_h_l_40')
// (6, 3, 'sp4_v_b_5')

reg n356 = 0;
// (2, 2, 'neigh_op_tnr_1')
// (2, 3, 'neigh_op_rgt_1')
// (2, 4, 'neigh_op_bnr_1')
// (3, 2, 'neigh_op_top_1')
// (3, 3, 'lutff_1/out')
// (3, 3, 'sp4_h_r_2')
// (3, 4, 'local_g0_1')
// (3, 4, 'lutff_7/in_0')
// (3, 4, 'neigh_op_bot_1')
// (4, 2, 'local_g2_1')
// (4, 2, 'lutff_4/in_3')
// (4, 2, 'neigh_op_tnl_1')
// (4, 3, 'neigh_op_lft_1')
// (4, 3, 'sp4_h_r_15')
// (4, 4, 'neigh_op_bnl_1')
// (5, 3, 'sp4_h_r_26')
// (6, 3, 'sp4_h_r_39')
// (6, 4, 'sp4_r_v_b_39')
// (6, 5, 'sp4_r_v_b_26')
// (6, 6, 'sp4_r_v_b_15')
// (6, 7, 'sp4_r_v_b_2')
// (7, 3, 'sp4_h_l_39')
// (7, 3, 'sp4_v_t_39')
// (7, 4, 'local_g2_7')
// (7, 4, 'lutff_1/in_2')
// (7, 4, 'sp4_v_b_39')
// (7, 5, 'sp4_v_b_26')
// (7, 6, 'sp4_v_b_15')
// (7, 7, 'sp4_v_b_2')

reg n357 = 0;
// (2, 2, 'neigh_op_tnr_2')
// (2, 3, 'neigh_op_rgt_2')
// (2, 4, 'neigh_op_bnr_2')
// (3, 1, 'sp4_r_v_b_45')
// (3, 2, 'neigh_op_top_2')
// (3, 2, 'sp4_r_v_b_32')
// (3, 3, 'lutff_2/out')
// (3, 3, 'sp4_h_r_4')
// (3, 3, 'sp4_r_v_b_21')
// (3, 4, 'neigh_op_bot_2')
// (3, 4, 'sp4_r_v_b_8')
// (4, 0, 'span4_vert_45')
// (4, 1, 'sp4_v_b_45')
// (4, 2, 'neigh_op_tnl_2')
// (4, 2, 'sp4_v_b_32')
// (4, 3, 'neigh_op_lft_2')
// (4, 3, 'sp4_h_r_17')
// (4, 3, 'sp4_v_b_21')
// (4, 4, 'neigh_op_bnl_2')
// (4, 4, 'sp4_h_r_8')
// (4, 4, 'sp4_v_b_8')
// (5, 3, 'local_g2_4')
// (5, 3, 'lutff_5/in_1')
// (5, 3, 'sp4_h_r_28')
// (5, 4, 'local_g0_5')
// (5, 4, 'lutff_4/in_3')
// (5, 4, 'sp4_h_r_21')
// (6, 3, 'sp4_h_r_41')
// (6, 4, 'sp4_h_r_32')
// (7, 3, 'sp4_h_l_41')
// (7, 4, 'local_g3_5')
// (7, 4, 'lutff_6/in_2')
// (7, 4, 'sp4_h_r_45')
// (8, 4, 'sp4_h_l_45')

wire n358;
// (2, 2, 'neigh_op_tnr_3')
// (2, 3, 'neigh_op_rgt_3')
// (2, 4, 'neigh_op_bnr_3')
// (3, 2, 'neigh_op_top_3')
// (3, 3, 'lutff_3/out')
// (3, 3, 'sp4_h_r_6')
// (3, 4, 'neigh_op_bot_3')
// (4, 2, 'neigh_op_tnl_3')
// (4, 3, 'neigh_op_lft_3')
// (4, 3, 'sp4_h_r_19')
// (4, 4, 'neigh_op_bnl_3')
// (5, 3, 'sp4_h_r_30')
// (6, 3, 'sp4_h_r_43')
// (6, 4, 'sp4_r_v_b_46')
// (6, 5, 'sp4_r_v_b_35')
// (6, 6, 'sp4_r_v_b_22')
// (6, 7, 'sp4_r_v_b_11')
// (7, 3, 'sp4_h_l_43')
// (7, 3, 'sp4_v_t_46')
// (7, 4, 'sp4_v_b_46')
// (7, 5, 'local_g2_3')
// (7, 5, 'lutff_1/in_2')
// (7, 5, 'sp4_v_b_35')
// (7, 6, 'sp4_v_b_22')
// (7, 7, 'sp4_v_b_11')

reg n359 = 0;
// (2, 2, 'neigh_op_tnr_4')
// (2, 2, 'sp4_r_v_b_37')
// (2, 3, 'neigh_op_rgt_4')
// (2, 3, 'sp4_r_v_b_24')
// (2, 4, 'neigh_op_bnr_4')
// (2, 4, 'sp4_r_v_b_13')
// (2, 5, 'sp4_r_v_b_0')
// (3, 1, 'sp4_h_r_5')
// (3, 1, 'sp4_v_t_37')
// (3, 2, 'neigh_op_top_4')
// (3, 2, 'sp4_v_b_37')
// (3, 3, 'lutff_4/out')
// (3, 3, 'sp4_h_r_8')
// (3, 3, 'sp4_v_b_24')
// (3, 4, 'neigh_op_bot_4')
// (3, 4, 'sp4_v_b_13')
// (3, 5, 'sp4_v_b_0')
// (4, 1, 'sp4_h_r_16')
// (4, 2, 'neigh_op_tnl_4')
// (4, 3, 'neigh_op_lft_4')
// (4, 3, 'sp4_h_r_21')
// (4, 4, 'neigh_op_bnl_4')
// (5, 1, 'local_g3_5')
// (5, 1, 'lutff_3/in_1')
// (5, 1, 'sp4_h_r_29')
// (5, 3, 'local_g3_0')
// (5, 3, 'lutff_4/in_3')
// (5, 3, 'lutff_7/in_0')
// (5, 3, 'sp4_h_r_32')
// (6, 1, 'sp4_h_r_40')
// (6, 3, 'sp4_h_r_45')
// (7, 1, 'sp4_h_l_40')
// (7, 3, 'sp4_h_l_45')

wire n360;
// (2, 2, 'neigh_op_tnr_5')
// (2, 3, 'neigh_op_rgt_5')
// (2, 4, 'neigh_op_bnr_5')
// (2, 4, 'sp4_r_v_b_41')
// (2, 5, 'sp4_r_v_b_28')
// (2, 6, 'sp4_r_v_b_17')
// (2, 7, 'sp4_r_v_b_4')
// (2, 8, 'sp4_r_v_b_41')
// (2, 9, 'sp4_r_v_b_28')
// (2, 10, 'sp4_r_v_b_17')
// (2, 11, 'local_g1_4')
// (2, 11, 'lutff_2/in_1')
// (2, 11, 'sp4_r_v_b_4')
// (3, 2, 'neigh_op_top_5')
// (3, 3, 'lutff_5/out')
// (3, 3, 'sp4_h_r_10')
// (3, 3, 'sp4_v_t_41')
// (3, 4, 'neigh_op_bot_5')
// (3, 4, 'sp4_v_b_41')
// (3, 5, 'sp4_v_b_28')
// (3, 6, 'sp4_v_b_17')
// (3, 7, 'sp4_v_b_4')
// (3, 7, 'sp4_v_t_41')
// (3, 8, 'sp4_v_b_41')
// (3, 9, 'sp4_v_b_28')
// (3, 10, 'sp4_v_b_17')
// (3, 11, 'sp4_v_b_4')
// (4, 2, 'neigh_op_tnl_5')
// (4, 3, 'neigh_op_lft_5')
// (4, 3, 'sp4_h_r_23')
// (4, 4, 'neigh_op_bnl_5')
// (5, 3, 'sp4_h_r_34')
// (6, 3, 'sp4_h_r_47')
// (7, 3, 'sp4_h_l_47')

wire n361;
// (2, 2, 'sp4_h_r_7')
// (3, 2, 'sp4_h_r_18')
// (4, 2, 'local_g3_7')
// (4, 2, 'lutff_6/in_2')
// (4, 2, 'sp4_h_r_31')
// (5, 2, 'sp4_h_r_42')
// (6, 2, 'sp4_h_l_42')
// (6, 2, 'sp4_h_r_4')
// (7, 1, 'neigh_op_tnr_6')
// (7, 2, 'neigh_op_rgt_6')
// (7, 2, 'sp4_h_r_17')
// (7, 3, 'neigh_op_bnr_6')
// (8, 1, 'neigh_op_top_6')
// (8, 2, 'lutff_6/out')
// (8, 2, 'sp4_h_r_28')
// (8, 3, 'neigh_op_bot_6')
// (9, 1, 'neigh_op_tnl_6')
// (9, 2, 'neigh_op_lft_6')
// (9, 2, 'sp4_h_r_41')
// (9, 3, 'neigh_op_bnl_6')
// (10, 2, 'sp4_h_l_41')

wire n362;
// (2, 2, 'sp4_r_v_b_43')
// (2, 3, 'sp4_r_v_b_30')
// (2, 4, 'sp4_r_v_b_19')
// (2, 5, 'sp4_r_v_b_6')
// (3, 1, 'sp4_v_t_43')
// (3, 2, 'sp4_v_b_43')
// (3, 3, 'local_g2_6')
// (3, 3, 'lutff_3/in_3')
// (3, 3, 'sp4_v_b_30')
// (3, 4, 'sp4_v_b_19')
// (3, 5, 'local_g0_6')
// (3, 5, 'lutff_0/in_0')
// (3, 5, 'sp4_h_r_6')
// (3, 5, 'sp4_v_b_6')
// (4, 2, 'sp4_r_v_b_42')
// (4, 3, 'sp4_r_v_b_31')
// (4, 4, 'sp4_r_v_b_18')
// (4, 5, 'sp4_h_r_19')
// (4, 5, 'sp4_r_v_b_7')
// (4, 6, 'sp4_r_v_b_42')
// (4, 7, 'sp4_r_v_b_31')
// (4, 8, 'sp4_r_v_b_18')
// (4, 9, 'sp4_r_v_b_7')
// (4, 10, 'sp4_r_v_b_47')
// (4, 11, 'sp4_r_v_b_34')
// (4, 12, 'sp4_r_v_b_23')
// (4, 13, 'sp4_r_v_b_10')
// (5, 1, 'local_g1_0')
// (5, 1, 'lutff_3/in_0')
// (5, 1, 'sp4_h_r_8')
// (5, 1, 'sp4_v_t_42')
// (5, 2, 'sp4_v_b_42')
// (5, 3, 'sp4_v_b_31')
// (5, 4, 'local_g1_2')
// (5, 4, 'lutff_2/in_1')
// (5, 4, 'sp4_v_b_18')
// (5, 5, 'sp4_h_r_30')
// (5, 5, 'sp4_h_r_7')
// (5, 5, 'sp4_v_b_7')
// (5, 5, 'sp4_v_t_42')
// (5, 6, 'sp4_v_b_42')
// (5, 7, 'sp4_v_b_31')
// (5, 8, 'sp4_v_b_18')
// (5, 9, 'sp4_v_b_7')
// (5, 9, 'sp4_v_t_47')
// (5, 10, 'sp4_v_b_47')
// (5, 11, 'sp4_v_b_34')
// (5, 12, 'sp4_v_b_23')
// (5, 13, 'local_g0_2')
// (5, 13, 'lutff_5/in_1')
// (5, 13, 'sp4_v_b_10')
// (6, 1, 'sp4_h_r_21')
// (6, 2, 'sp4_r_v_b_38')
// (6, 3, 'sp4_r_v_b_27')
// (6, 4, 'sp4_r_v_b_14')
// (6, 5, 'sp4_h_r_18')
// (6, 5, 'sp4_h_r_43')
// (6, 5, 'sp4_r_v_b_3')
// (6, 6, 'sp4_r_v_b_47')
// (6, 7, 'sp4_r_v_b_34')
// (6, 8, 'sp4_r_v_b_23')
// (6, 9, 'sp4_r_v_b_10')
// (6, 10, 'sp4_r_v_b_36')
// (6, 11, 'sp4_h_r_7')
// (6, 11, 'sp4_r_v_b_25')
// (6, 12, 'sp4_r_v_b_12')
// (6, 13, 'sp4_r_v_b_1')
// (7, 1, 'sp4_h_r_32')
// (7, 1, 'sp4_v_t_38')
// (7, 2, 'sp4_v_b_38')
// (7, 3, 'sp4_v_b_27')
// (7, 4, 'local_g0_6')
// (7, 4, 'lutff_1/in_1')
// (7, 4, 'lutff_2/in_0')
// (7, 4, 'lutff_3/in_1')
// (7, 4, 'lutff_6/in_0')
// (7, 4, 'sp4_v_b_14')
// (7, 5, 'local_g0_2')
// (7, 5, 'lutff_0/in_2')
// (7, 5, 'lutff_1/in_3')
// (7, 5, 'lutff_5/in_1')
// (7, 5, 'sp4_h_l_43')
// (7, 5, 'sp4_h_r_10')
// (7, 5, 'sp4_h_r_31')
// (7, 5, 'sp4_v_b_3')
// (7, 5, 'sp4_v_t_47')
// (7, 6, 'sp4_v_b_47')
// (7, 7, 'sp4_v_b_34')
// (7, 8, 'sp4_v_b_23')
// (7, 9, 'sp4_v_b_10')
// (7, 9, 'sp4_v_t_36')
// (7, 10, 'sp4_v_b_36')
// (7, 11, 'local_g1_2')
// (7, 11, 'lutff_0/in_1')
// (7, 11, 'sp4_h_r_18')
// (7, 11, 'sp4_v_b_25')
// (7, 12, 'sp4_v_b_12')
// (7, 13, 'local_g0_1')
// (7, 13, 'lutff_1/in_2')
// (7, 13, 'lutff_7/in_0')
// (7, 13, 'sp4_v_b_1')
// (8, 1, 'sp4_h_r_45')
// (8, 2, 'sp4_r_v_b_39')
// (8, 3, 'sp4_r_v_b_26')
// (8, 4, 'neigh_op_tnr_1')
// (8, 4, 'sp4_r_v_b_15')
// (8, 4, 'sp4_r_v_b_47')
// (8, 5, 'neigh_op_rgt_1')
// (8, 5, 'sp4_h_r_23')
// (8, 5, 'sp4_h_r_42')
// (8, 5, 'sp4_r_v_b_2')
// (8, 5, 'sp4_r_v_b_34')
// (8, 6, 'neigh_op_bnr_1')
// (8, 6, 'sp4_r_v_b_23')
// (8, 7, 'sp4_r_v_b_10')
// (8, 8, 'sp4_r_v_b_43')
// (8, 9, 'sp4_r_v_b_30')
// (8, 10, 'local_g3_3')
// (8, 10, 'lutff_4/in_0')
// (8, 10, 'sp4_r_v_b_19')
// (8, 11, 'local_g1_6')
// (8, 11, 'lutff_2/in_3')
// (8, 11, 'lutff_3/in_0')
// (8, 11, 'sp4_h_r_31')
// (8, 11, 'sp4_r_v_b_6')
// (9, 1, 'sp4_h_l_45')
// (9, 1, 'sp4_v_t_39')
// (9, 2, 'sp12_v_t_22')
// (9, 2, 'sp4_v_b_39')
// (9, 3, 'sp12_v_b_22')
// (9, 3, 'sp4_v_b_26')
// (9, 3, 'sp4_v_t_47')
// (9, 4, 'neigh_op_top_1')
// (9, 4, 'sp12_v_b_21')
// (9, 4, 'sp4_r_v_b_46')
// (9, 4, 'sp4_v_b_15')
// (9, 4, 'sp4_v_b_47')
// (9, 5, 'local_g3_1')
// (9, 5, 'lutff_1/out')
// (9, 5, 'lutff_7/in_3')
// (9, 5, 'sp12_v_b_18')
// (9, 5, 'sp4_h_l_42')
// (9, 5, 'sp4_h_r_34')
// (9, 5, 'sp4_r_v_b_35')
// (9, 5, 'sp4_v_b_2')
// (9, 5, 'sp4_v_b_34')
// (9, 6, 'neigh_op_bot_1')
// (9, 6, 'sp12_v_b_17')
// (9, 6, 'sp4_r_v_b_22')
// (9, 6, 'sp4_v_b_23')
// (9, 7, 'sp12_v_b_14')
// (9, 7, 'sp4_r_v_b_11')
// (9, 7, 'sp4_v_b_10')
// (9, 7, 'sp4_v_t_43')
// (9, 8, 'sp12_v_b_13')
// (9, 8, 'sp4_r_v_b_39')
// (9, 8, 'sp4_v_b_43')
// (9, 9, 'sp12_v_b_10')
// (9, 9, 'sp4_r_v_b_26')
// (9, 9, 'sp4_v_b_30')
// (9, 10, 'local_g1_3')
// (9, 10, 'lutff_1/in_3')
// (9, 10, 'lutff_3/in_3')
// (9, 10, 'sp12_v_b_9')
// (9, 10, 'sp4_r_v_b_15')
// (9, 10, 'sp4_v_b_19')
// (9, 11, 'sp12_v_b_6')
// (9, 11, 'sp4_h_r_42')
// (9, 11, 'sp4_r_v_b_2')
// (9, 11, 'sp4_v_b_6')
// (9, 12, 'local_g2_5')
// (9, 12, 'lutff_7/in_2')
// (9, 12, 'sp12_v_b_5')
// (9, 13, 'local_g2_2')
// (9, 13, 'lutff_0/in_2')
// (9, 13, 'lutff_6/in_2')
// (9, 13, 'lutff_7/in_3')
// (9, 13, 'sp12_v_b_2')
// (9, 14, 'sp12_v_b_1')
// (10, 3, 'sp4_v_t_46')
// (10, 4, 'neigh_op_tnl_1')
// (10, 4, 'sp4_v_b_46')
// (10, 5, 'neigh_op_lft_1')
// (10, 5, 'sp4_h_r_47')
// (10, 5, 'sp4_v_b_35')
// (10, 6, 'neigh_op_bnl_1')
// (10, 6, 'sp4_v_b_22')
// (10, 7, 'sp4_v_b_11')
// (10, 7, 'sp4_v_t_39')
// (10, 8, 'sp4_v_b_39')
// (10, 9, 'sp4_v_b_26')
// (10, 10, 'sp4_v_b_15')
// (10, 11, 'sp4_h_l_42')
// (10, 11, 'sp4_v_b_2')
// (11, 5, 'sp4_h_l_47')

wire n363;
// (2, 2, 'sp4_r_v_b_46')
// (2, 3, 'sp4_r_v_b_35')
// (2, 4, 'sp4_r_v_b_22')
// (2, 5, 'sp4_r_v_b_11')
// (2, 6, 'sp4_r_v_b_45')
// (2, 7, 'local_g2_0')
// (2, 7, 'lutff_7/in_3')
// (2, 7, 'sp4_r_v_b_32')
// (2, 8, 'sp4_r_v_b_21')
// (2, 9, 'sp4_r_v_b_8')
// (2, 10, 'sp4_r_v_b_45')
// (2, 11, 'sp4_r_v_b_32')
// (2, 12, 'sp4_r_v_b_21')
// (2, 13, 'sp4_r_v_b_8')
// (2, 14, 'sp4_r_v_b_45')
// (2, 15, 'sp4_r_v_b_32')
// (2, 16, 'neigh_op_tnr_4')
// (2, 16, 'sp4_r_v_b_21')
// (2, 17, 'local_g2_4')
// (2, 17, 'lutff_7/in_3')
// (2, 17, 'neigh_op_rgt_4')
// (2, 17, 'sp4_r_v_b_8')
// (2, 18, 'neigh_op_bnr_4')
// (3, 1, 'sp4_v_t_46')
// (3, 2, 'sp4_v_b_46')
// (3, 3, 'local_g2_3')
// (3, 3, 'lutff_5/in_0')
// (3, 3, 'sp4_v_b_35')
// (3, 4, 'sp4_v_b_22')
// (3, 5, 'sp4_v_b_11')
// (3, 5, 'sp4_v_t_45')
// (3, 6, 'sp4_v_b_45')
// (3, 7, 'local_g3_0')
// (3, 7, 'lutff_1/in_0')
// (3, 7, 'sp4_v_b_32')
// (3, 8, 'sp4_v_b_21')
// (3, 9, 'sp4_v_b_8')
// (3, 9, 'sp4_v_t_45')
// (3, 10, 'sp4_v_b_45')
// (3, 11, 'sp4_v_b_32')
// (3, 12, 'sp4_v_b_21')
// (3, 13, 'sp4_v_b_8')
// (3, 13, 'sp4_v_t_45')
// (3, 14, 'sp4_v_b_45')
// (3, 15, 'sp4_v_b_32')
// (3, 16, 'neigh_op_top_4')
// (3, 16, 'sp4_v_b_21')
// (3, 17, 'lutff_4/out')
// (3, 17, 'sp4_v_b_8')
// (3, 18, 'neigh_op_bot_4')
// (4, 16, 'neigh_op_tnl_4')
// (4, 17, 'neigh_op_lft_4')
// (4, 18, 'neigh_op_bnl_4')

wire n364;
// (2, 3, 'neigh_op_tnr_1')
// (2, 4, 'neigh_op_rgt_1')
// (2, 5, 'neigh_op_bnr_1')
// (3, 3, 'neigh_op_top_1')
// (3, 4, 'lutff_1/out')
// (3, 5, 'local_g1_1')
// (3, 5, 'lutff_3/in_3')
// (3, 5, 'neigh_op_bot_1')
// (4, 3, 'neigh_op_tnl_1')
// (4, 4, 'neigh_op_lft_1')
// (4, 5, 'neigh_op_bnl_1')

reg n365 = 0;
// (2, 3, 'neigh_op_tnr_2')
// (2, 4, 'neigh_op_rgt_2')
// (2, 4, 'sp4_h_r_9')
// (2, 5, 'neigh_op_bnr_2')
// (3, 3, 'neigh_op_top_2')
// (3, 4, 'lutff_2/out')
// (3, 4, 'sp4_h_r_20')
// (3, 5, 'local_g0_2')
// (3, 5, 'lutff_6/in_0')
// (3, 5, 'neigh_op_bot_2')
// (4, 3, 'neigh_op_tnl_2')
// (4, 4, 'neigh_op_lft_2')
// (4, 4, 'sp4_h_r_33')
// (4, 5, 'local_g3_2')
// (4, 5, 'lutff_3/in_0')
// (4, 5, 'neigh_op_bnl_2')
// (5, 4, 'sp4_h_r_44')
// (5, 5, 'sp4_r_v_b_44')
// (5, 6, 'local_g2_1')
// (5, 6, 'lutff_3/in_0')
// (5, 6, 'sp4_r_v_b_33')
// (5, 7, 'sp4_r_v_b_20')
// (5, 8, 'sp4_r_v_b_9')
// (6, 4, 'sp4_h_l_44')
// (6, 4, 'sp4_v_t_44')
// (6, 5, 'sp4_v_b_44')
// (6, 6, 'sp4_v_b_33')
// (6, 7, 'sp4_v_b_20')
// (6, 8, 'sp4_v_b_9')

wire n366;
// (2, 3, 'neigh_op_tnr_3')
// (2, 4, 'neigh_op_rgt_3')
// (2, 5, 'neigh_op_bnr_3')
// (3, 3, 'local_g1_3')
// (3, 3, 'lutff_5/in_3')
// (3, 3, 'neigh_op_top_3')
// (3, 4, 'lutff_3/out')
// (3, 5, 'neigh_op_bot_3')
// (4, 3, 'neigh_op_tnl_3')
// (4, 4, 'neigh_op_lft_3')
// (4, 5, 'neigh_op_bnl_3')

wire n367;
// (2, 3, 'neigh_op_tnr_4')
// (2, 4, 'local_g2_4')
// (2, 4, 'lutff_5/in_1')
// (2, 4, 'neigh_op_rgt_4')
// (2, 5, 'neigh_op_bnr_4')
// (3, 3, 'neigh_op_top_4')
// (3, 4, 'lutff_4/out')
// (3, 5, 'neigh_op_bot_4')
// (4, 3, 'neigh_op_tnl_4')
// (4, 4, 'neigh_op_lft_4')
// (4, 5, 'neigh_op_bnl_4')

wire n368;
// (2, 3, 'neigh_op_tnr_5')
// (2, 4, 'neigh_op_rgt_5')
// (2, 5, 'neigh_op_bnr_5')
// (3, 3, 'neigh_op_top_5')
// (3, 4, 'local_g2_5')
// (3, 4, 'lutff_4/in_3')
// (3, 4, 'lutff_5/out')
// (3, 5, 'neigh_op_bot_5')
// (4, 3, 'neigh_op_tnl_5')
// (4, 4, 'neigh_op_lft_5')
// (4, 5, 'neigh_op_bnl_5')

wire n369;
// (2, 3, 'neigh_op_tnr_6')
// (2, 4, 'neigh_op_rgt_6')
// (2, 5, 'neigh_op_bnr_6')
// (3, 3, 'neigh_op_top_6')
// (3, 4, 'local_g2_6')
// (3, 4, 'lutff_1/in_1')
// (3, 4, 'lutff_6/out')
// (3, 5, 'neigh_op_bot_6')
// (4, 3, 'neigh_op_tnl_6')
// (4, 4, 'neigh_op_lft_6')
// (4, 5, 'neigh_op_bnl_6')

wire n370;
// (2, 3, 'neigh_op_tnr_7')
// (2, 4, 'neigh_op_rgt_7')
// (2, 5, 'neigh_op_bnr_7')
// (3, 3, 'neigh_op_top_7')
// (3, 4, 'lutff_7/out')
// (3, 5, 'neigh_op_bot_7')
// (4, 3, 'neigh_op_tnl_7')
// (4, 4, 'local_g0_7')
// (4, 4, 'lutff_7/in_0')
// (4, 4, 'neigh_op_lft_7')
// (4, 5, 'neigh_op_bnl_7')

reg n371 = 0;
// (2, 3, 'sp4_r_v_b_47')
// (2, 4, 'sp4_r_v_b_34')
// (2, 5, 'local_g3_7')
// (2, 5, 'lutff_2/in_0')
// (2, 5, 'sp4_r_v_b_23')
// (2, 6, 'sp4_r_v_b_10')
// (3, 1, 'sp4_r_v_b_40')
// (3, 2, 'local_g0_5')
// (3, 2, 'lutff_0/in_3')
// (3, 2, 'sp4_r_v_b_29')
// (3, 2, 'sp4_v_t_47')
// (3, 3, 'sp4_r_v_b_16')
// (3, 3, 'sp4_v_b_47')
// (3, 4, 'local_g1_5')
// (3, 4, 'lutff_6/in_0')
// (3, 4, 'sp4_r_v_b_5')
// (3, 4, 'sp4_v_b_34')
// (3, 5, 'sp4_r_v_b_40')
// (3, 5, 'sp4_v_b_23')
// (3, 6, 'local_g1_0')
// (3, 6, 'lutff_5/in_2')
// (3, 6, 'sp4_h_r_0')
// (3, 6, 'sp4_h_r_5')
// (3, 6, 'sp4_r_v_b_29')
// (3, 6, 'sp4_v_b_10')
// (3, 7, 'sp4_r_v_b_16')
// (3, 8, 'sp4_r_v_b_5')
// (4, 0, 'span4_vert_40')
// (4, 1, 'local_g3_0')
// (4, 1, 'lutff_5/in_2')
// (4, 1, 'sp4_v_b_40')
// (4, 2, 'sp4_v_b_29')
// (4, 3, 'sp4_v_b_16')
// (4, 4, 'sp4_h_r_5')
// (4, 4, 'sp4_v_b_5')
// (4, 4, 'sp4_v_t_40')
// (4, 5, 'local_g3_0')
// (4, 5, 'lutff_0/in_3')
// (4, 5, 'sp4_r_v_b_37')
// (4, 5, 'sp4_v_b_40')
// (4, 6, 'local_g1_0')
// (4, 6, 'lutff_2/in_3')
// (4, 6, 'sp4_h_r_13')
// (4, 6, 'sp4_h_r_16')
// (4, 6, 'sp4_r_v_b_24')
// (4, 6, 'sp4_v_b_29')
// (4, 7, 'local_g0_0')
// (4, 7, 'lutff_1/in_1')
// (4, 7, 'sp4_r_v_b_13')
// (4, 7, 'sp4_v_b_16')
// (4, 8, 'sp4_r_v_b_0')
// (4, 8, 'sp4_v_b_5')
// (5, 4, 'sp4_h_r_0')
// (5, 4, 'sp4_h_r_16')
// (5, 4, 'sp4_v_t_37')
// (5, 5, 'sp4_v_b_37')
// (5, 6, 'sp4_h_r_24')
// (5, 6, 'sp4_h_r_29')
// (5, 6, 'sp4_v_b_24')
// (5, 7, 'sp4_v_b_13')
// (5, 8, 'local_g0_0')
// (5, 8, 'lutff_0/in_0')
// (5, 8, 'sp4_v_b_0')
// (6, 3, 'neigh_op_tnr_4')
// (6, 3, 'sp4_r_v_b_37')
// (6, 4, 'neigh_op_rgt_4')
// (6, 4, 'sp4_h_r_13')
// (6, 4, 'sp4_h_r_29')
// (6, 4, 'sp4_r_v_b_24')
// (6, 5, 'neigh_op_bnr_4')
// (6, 5, 'sp4_r_v_b_13')
// (6, 6, 'sp4_h_r_37')
// (6, 6, 'sp4_h_r_40')
// (6, 6, 'sp4_r_v_b_0')
// (7, 2, 'sp4_v_t_37')
// (7, 3, 'local_g1_4')
// (7, 3, 'lutff_4/in_3')
// (7, 3, 'neigh_op_top_4')
// (7, 3, 'sp4_v_b_37')
// (7, 4, 'lutff_4/out')
// (7, 4, 'sp4_h_r_24')
// (7, 4, 'sp4_h_r_40')
// (7, 4, 'sp4_v_b_24')
// (7, 5, 'neigh_op_bot_4')
// (7, 5, 'sp4_v_b_13')
// (7, 6, 'sp4_h_l_37')
// (7, 6, 'sp4_h_l_40')
// (7, 6, 'sp4_v_b_0')
// (8, 3, 'neigh_op_tnl_4')
// (8, 4, 'neigh_op_lft_4')
// (8, 4, 'sp4_h_l_40')
// (8, 4, 'sp4_h_r_37')
// (8, 5, 'neigh_op_bnl_4')
// (9, 4, 'sp4_h_l_37')

wire n372;
// (2, 4, 'local_g0_2')
// (2, 4, 'lutff_5/in_3')
// (2, 4, 'sp4_h_r_2')
// (2, 7, 'local_g0_1')
// (2, 7, 'lutff_3/in_0')
// (2, 7, 'sp4_h_r_1')
// (3, 1, 'sp4_r_v_b_33')
// (3, 2, 'local_g3_4')
// (3, 2, 'lutff_6/in_3')
// (3, 2, 'sp4_r_v_b_20')
// (3, 3, 'sp4_r_v_b_9')
// (3, 4, 'sp4_h_r_15')
// (3, 4, 'sp4_r_v_b_44')
// (3, 5, 'sp4_r_v_b_33')
// (3, 6, 'sp4_r_v_b_20')
// (3, 7, 'sp4_h_r_12')
// (3, 7, 'sp4_r_v_b_9')
// (4, 0, 'span4_vert_33')
// (4, 1, 'sp4_v_b_33')
// (4, 2, 'sp4_v_b_20')
// (4, 3, 'sp4_v_b_9')
// (4, 3, 'sp4_v_t_44')
// (4, 4, 'sp4_h_r_26')
// (4, 4, 'sp4_r_v_b_41')
// (4, 4, 'sp4_v_b_44')
// (4, 5, 'local_g0_4')
// (4, 5, 'lutff_0/in_0')
// (4, 5, 'sp4_r_v_b_28')
// (4, 5, 'sp4_v_b_33')
// (4, 6, 'local_g2_2')
// (4, 6, 'lutff_2/in_0')
// (4, 6, 'lutff_3/in_3')
// (4, 6, 'neigh_op_tnr_2')
// (4, 6, 'sp4_r_v_b_17')
// (4, 6, 'sp4_v_b_20')
// (4, 7, 'local_g3_1')
// (4, 7, 'lutff_6/in_0')
// (4, 7, 'neigh_op_rgt_2')
// (4, 7, 'sp4_h_r_25')
// (4, 7, 'sp4_h_r_9')
// (4, 7, 'sp4_r_v_b_4')
// (4, 7, 'sp4_v_b_9')
// (4, 8, 'neigh_op_bnr_2')
// (5, 3, 'sp4_v_t_41')
// (5, 4, 'sp4_h_r_39')
// (5, 4, 'sp4_v_b_41')
// (5, 5, 'sp4_r_v_b_45')
// (5, 5, 'sp4_v_b_28')
// (5, 6, 'neigh_op_top_2')
// (5, 6, 'sp4_r_v_b_32')
// (5, 6, 'sp4_v_b_17')
// (5, 7, 'lutff_2/out')
// (5, 7, 'sp4_h_r_20')
// (5, 7, 'sp4_h_r_36')
// (5, 7, 'sp4_r_v_b_21')
// (5, 7, 'sp4_v_b_4')
// (5, 8, 'neigh_op_bot_2')
// (5, 8, 'sp4_r_v_b_8')
// (6, 4, 'sp4_h_l_39')
// (6, 4, 'sp4_v_t_45')
// (6, 5, 'sp4_v_b_45')
// (6, 6, 'neigh_op_tnl_2')
// (6, 6, 'sp4_v_b_32')
// (6, 7, 'neigh_op_lft_2')
// (6, 7, 'sp4_h_l_36')
// (6, 7, 'sp4_h_r_33')
// (6, 7, 'sp4_v_b_21')
// (6, 8, 'neigh_op_bnl_2')
// (6, 8, 'sp4_v_b_8')
// (7, 7, 'sp4_h_r_44')
// (8, 7, 'sp4_h_l_44')

wire n373;
// (2, 4, 'neigh_op_tnr_0')
// (2, 5, 'neigh_op_rgt_0')
// (2, 5, 'sp4_h_r_5')
// (2, 6, 'neigh_op_bnr_0')
// (3, 4, 'neigh_op_top_0')
// (3, 5, 'lutff_0/out')
// (3, 5, 'sp4_h_r_16')
// (3, 6, 'neigh_op_bot_0')
// (4, 4, 'neigh_op_tnl_0')
// (4, 5, 'neigh_op_lft_0')
// (4, 5, 'sp4_h_r_29')
// (4, 6, 'neigh_op_bnl_0')
// (5, 5, 'sp4_h_r_40')
// (6, 5, 'sp4_h_l_40')
// (6, 5, 'sp4_h_r_5')
// (7, 5, 'local_g1_0')
// (7, 5, 'lutff_5/in_2')
// (7, 5, 'sp4_h_r_16')
// (8, 5, 'sp4_h_r_29')
// (9, 5, 'sp4_h_r_40')
// (10, 5, 'sp4_h_l_40')

wire n374;
// (2, 4, 'neigh_op_tnr_1')
// (2, 5, 'neigh_op_rgt_1')
// (2, 6, 'local_g1_1')
// (2, 6, 'lutff_6/in_0')
// (2, 6, 'neigh_op_bnr_1')
// (3, 3, 'sp4_r_v_b_43')
// (3, 4, 'neigh_op_top_1')
// (3, 4, 'sp4_r_v_b_30')
// (3, 5, 'lutff_1/out')
// (3, 5, 'sp4_r_v_b_19')
// (3, 6, 'neigh_op_bot_1')
// (3, 6, 'sp4_r_v_b_6')
// (4, 2, 'sp4_v_t_43')
// (4, 3, 'sp4_v_b_43')
// (4, 4, 'neigh_op_tnl_1')
// (4, 4, 'sp4_v_b_30')
// (4, 5, 'neigh_op_lft_1')
// (4, 5, 'sp4_v_b_19')
// (4, 6, 'local_g0_6')
// (4, 6, 'lutff_2/in_2')
// (4, 6, 'neigh_op_bnl_1')
// (4, 6, 'sp4_v_b_6')

wire n375;
// (2, 4, 'neigh_op_tnr_2')
// (2, 5, 'local_g2_2')
// (2, 5, 'lutff_4/in_0')
// (2, 5, 'neigh_op_rgt_2')
// (2, 6, 'neigh_op_bnr_2')
// (3, 4, 'neigh_op_top_2')
// (3, 5, 'lutff_2/out')
// (3, 6, 'neigh_op_bot_2')
// (4, 4, 'neigh_op_tnl_2')
// (4, 5, 'neigh_op_lft_2')
// (4, 6, 'neigh_op_bnl_2')

wire n376;
// (2, 4, 'neigh_op_tnr_3')
// (2, 5, 'neigh_op_rgt_3')
// (2, 6, 'neigh_op_bnr_3')
// (3, 4, 'local_g0_3')
// (3, 4, 'lutff_3/in_2')
// (3, 4, 'neigh_op_top_3')
// (3, 5, 'lutff_3/out')
// (3, 6, 'neigh_op_bot_3')
// (4, 4, 'neigh_op_tnl_3')
// (4, 5, 'neigh_op_lft_3')
// (4, 6, 'neigh_op_bnl_3')

wire n377;
// (2, 4, 'neigh_op_tnr_4')
// (2, 5, 'neigh_op_rgt_4')
// (2, 6, 'neigh_op_bnr_4')
// (3, 4, 'neigh_op_top_4')
// (3, 5, 'local_g0_4')
// (3, 5, 'lutff_4/out')
// (3, 5, 'lutff_5/in_1')
// (3, 6, 'neigh_op_bot_4')
// (4, 4, 'neigh_op_tnl_4')
// (4, 5, 'neigh_op_lft_4')
// (4, 6, 'neigh_op_bnl_4')

wire n378;
// (2, 4, 'neigh_op_tnr_5')
// (2, 5, 'neigh_op_rgt_5')
// (2, 6, 'neigh_op_bnr_5')
// (3, 4, 'neigh_op_top_5')
// (3, 5, 'lutff_5/out')
// (3, 6, 'neigh_op_bot_5')
// (4, 4, 'neigh_op_tnl_5')
// (4, 5, 'local_g1_5')
// (4, 5, 'lutff_4/in_0')
// (4, 5, 'neigh_op_lft_5')
// (4, 6, 'neigh_op_bnl_5')

wire n379;
// (2, 4, 'neigh_op_tnr_6')
// (2, 5, 'neigh_op_rgt_6')
// (2, 6, 'neigh_op_bnr_6')
// (3, 4, 'neigh_op_top_6')
// (3, 5, 'lutff_6/out')
// (3, 6, 'neigh_op_bot_6')
// (4, 4, 'local_g2_6')
// (4, 4, 'lutff_0/in_0')
// (4, 4, 'neigh_op_tnl_6')
// (4, 5, 'neigh_op_lft_6')
// (4, 6, 'neigh_op_bnl_6')

reg n380 = 0;
// (2, 4, 'sp4_h_r_10')
// (3, 4, 'local_g1_7')
// (3, 4, 'lutff_7/in_1')
// (3, 4, 'sp4_h_r_23')
// (3, 4, 'sp4_r_v_b_46')
// (3, 5, 'local_g0_0')
// (3, 5, 'lutff_0/in_2')
// (3, 5, 'sp4_r_v_b_35')
// (3, 6, 'sp4_r_v_b_22')
// (3, 7, 'sp4_r_v_b_11')
// (4, 2, 'neigh_op_tnr_3')
// (4, 3, 'neigh_op_rgt_3')
// (4, 3, 'sp4_h_r_11')
// (4, 3, 'sp4_v_t_46')
// (4, 4, 'neigh_op_bnr_3')
// (4, 4, 'sp4_h_r_34')
// (4, 4, 'sp4_v_b_46')
// (4, 5, 'sp4_v_b_35')
// (4, 6, 'sp4_v_b_22')
// (4, 7, 'sp4_v_b_11')
// (5, 1, 'sp4_r_v_b_47')
// (5, 2, 'neigh_op_top_3')
// (5, 2, 'sp4_r_v_b_34')
// (5, 3, 'local_g3_3')
// (5, 3, 'lutff_3/out')
// (5, 3, 'lutff_4/in_0')
// (5, 3, 'sp4_h_r_22')
// (5, 3, 'sp4_r_v_b_23')
// (5, 4, 'neigh_op_bot_3')
// (5, 4, 'sp4_h_r_47')
// (5, 4, 'sp4_r_v_b_10')
// (6, 0, 'span4_vert_47')
// (6, 1, 'sp4_v_b_47')
// (6, 2, 'neigh_op_tnl_3')
// (6, 2, 'sp4_v_b_34')
// (6, 3, 'neigh_op_lft_3')
// (6, 3, 'sp4_h_r_35')
// (6, 3, 'sp4_v_b_23')
// (6, 4, 'neigh_op_bnl_3')
// (6, 4, 'sp4_h_l_47')
// (6, 4, 'sp4_v_b_10')
// (7, 3, 'sp4_h_r_46')
// (8, 3, 'sp4_h_l_46')

reg n381 = 0;
// (2, 4, 'sp4_h_r_4')
// (3, 2, 'sp4_r_v_b_36')
// (3, 3, 'neigh_op_tnr_6')
// (3, 3, 'sp4_r_v_b_25')
// (3, 4, 'neigh_op_rgt_6')
// (3, 4, 'sp4_h_r_17')
// (3, 4, 'sp4_r_v_b_12')
// (3, 5, 'neigh_op_bnr_6')
// (3, 5, 'sp4_r_v_b_1')
// (4, 1, 'sp4_v_t_36')
// (4, 2, 'local_g2_4')
// (4, 2, 'lutff_4/in_0')
// (4, 2, 'sp4_v_b_36')
// (4, 3, 'neigh_op_top_6')
// (4, 3, 'sp4_v_b_25')
// (4, 4, 'lutff_6/out')
// (4, 4, 'sp4_h_r_28')
// (4, 4, 'sp4_v_b_12')
// (4, 5, 'neigh_op_bot_6')
// (4, 5, 'sp4_v_b_1')
// (5, 3, 'neigh_op_tnl_6')
// (5, 4, 'local_g1_6')
// (5, 4, 'lutff_6/in_1')
// (5, 4, 'neigh_op_lft_6')
// (5, 4, 'sp4_h_r_41')
// (5, 5, 'neigh_op_bnl_6')
// (6, 4, 'sp4_h_l_41')
// (6, 4, 'sp4_h_r_7')
// (7, 4, 'local_g1_2')
// (7, 4, 'lutff_2/in_1')
// (7, 4, 'sp4_h_r_18')
// (8, 4, 'sp4_h_r_31')
// (9, 4, 'sp4_h_r_42')
// (10, 4, 'sp4_h_l_42')

reg n382 = 0;
// (2, 5, 'local_g2_3')
// (2, 5, 'lutff_7/in_2')
// (2, 5, 'neigh_op_tnr_3')
// (2, 6, 'neigh_op_rgt_3')
// (2, 6, 'sp4_h_r_11')
// (2, 7, 'neigh_op_bnr_3')
// (3, 5, 'neigh_op_top_3')
// (3, 6, 'lutff_3/out')
// (3, 6, 'sp4_h_r_22')
// (3, 6, 'sp4_r_v_b_39')
// (3, 7, 'neigh_op_bot_3')
// (3, 7, 'sp4_r_v_b_26')
// (3, 8, 'sp4_r_v_b_15')
// (3, 9, 'sp4_r_v_b_2')
// (4, 5, 'neigh_op_tnl_3')
// (4, 5, 'sp4_v_t_39')
// (4, 6, 'neigh_op_lft_3')
// (4, 6, 'sp4_h_r_35')
// (4, 6, 'sp4_v_b_39')
// (4, 7, 'neigh_op_bnl_3')
// (4, 7, 'sp4_v_b_26')
// (4, 8, 'sp4_v_b_15')
// (4, 9, 'local_g0_2')
// (4, 9, 'lutff_5/in_1')
// (4, 9, 'sp4_v_b_2')
// (5, 3, 'sp4_r_v_b_40')
// (5, 4, 'sp4_r_v_b_29')
// (5, 5, 'local_g3_0')
// (5, 5, 'lutff_5/in_2')
// (5, 5, 'sp4_r_v_b_16')
// (5, 6, 'sp4_h_r_46')
// (5, 6, 'sp4_r_v_b_5')
// (6, 2, 'sp4_v_t_40')
// (6, 3, 'sp4_v_b_40')
// (6, 4, 'sp4_v_b_29')
// (6, 5, 'sp4_v_b_16')
// (6, 6, 'sp4_h_l_46')
// (6, 6, 'sp4_v_b_5')

wire n383;
// (2, 5, 'local_g3_6')
// (2, 5, 'lutff_0/in_1')
// (2, 5, 'neigh_op_tnr_6')
// (2, 6, 'neigh_op_rgt_6')
// (2, 7, 'neigh_op_bnr_6')
// (3, 4, 'sp4_r_v_b_37')
// (3, 5, 'neigh_op_top_6')
// (3, 5, 'sp4_r_v_b_24')
// (3, 6, 'lutff_6/out')
// (3, 6, 'sp4_r_v_b_13')
// (3, 7, 'neigh_op_bot_6')
// (3, 7, 'sp4_r_v_b_0')
// (4, 3, 'sp4_h_r_0')
// (4, 3, 'sp4_v_t_37')
// (4, 4, 'sp4_v_b_37')
// (4, 5, 'neigh_op_tnl_6')
// (4, 5, 'sp4_v_b_24')
// (4, 6, 'neigh_op_lft_6')
// (4, 6, 'sp4_v_b_13')
// (4, 7, 'neigh_op_bnl_6')
// (4, 7, 'sp4_v_b_0')
// (5, 3, 'local_g0_5')
// (5, 3, 'lutff_2/in_3')
// (5, 3, 'sp4_h_r_13')
// (6, 3, 'sp4_h_r_24')
// (7, 3, 'sp4_h_r_37')
// (8, 3, 'sp4_h_l_37')

wire n384;
// (2, 5, 'neigh_op_tnr_0')
// (2, 6, 'neigh_op_rgt_0')
// (2, 7, 'neigh_op_bnr_0')
// (3, 5, 'local_g1_0')
// (3, 5, 'lutff_3/in_0')
// (3, 5, 'neigh_op_top_0')
// (3, 6, 'lutff_0/out')
// (3, 7, 'neigh_op_bot_0')
// (4, 5, 'neigh_op_tnl_0')
// (4, 6, 'neigh_op_lft_0')
// (4, 7, 'neigh_op_bnl_0')

wire n385;
// (2, 5, 'neigh_op_tnr_1')
// (2, 6, 'neigh_op_rgt_1')
// (2, 7, 'neigh_op_bnr_1')
// (3, 5, 'neigh_op_top_1')
// (3, 6, 'lutff_1/out')
// (3, 7, 'neigh_op_bot_1')
// (4, 5, 'neigh_op_tnl_1')
// (4, 6, 'local_g0_1')
// (4, 6, 'lutff_3/in_0')
// (4, 6, 'neigh_op_lft_1')
// (4, 7, 'neigh_op_bnl_1')

wire n386;
// (2, 5, 'neigh_op_tnr_2')
// (2, 6, 'neigh_op_rgt_2')
// (2, 7, 'neigh_op_bnr_2')
// (3, 5, 'neigh_op_top_2')
// (3, 6, 'lutff_2/out')
// (3, 7, 'neigh_op_bot_2')
// (4, 5, 'neigh_op_tnl_2')
// (4, 6, 'local_g1_2')
// (4, 6, 'lutff_7/in_2')
// (4, 6, 'neigh_op_lft_2')
// (4, 7, 'neigh_op_bnl_2')

wire n387;
// (2, 5, 'neigh_op_tnr_5')
// (2, 6, 'neigh_op_rgt_5')
// (2, 7, 'neigh_op_bnr_5')
// (3, 5, 'neigh_op_top_5')
// (3, 6, 'local_g3_5')
// (3, 6, 'lutff_0/in_2')
// (3, 6, 'lutff_5/out')
// (3, 7, 'neigh_op_bot_5')
// (4, 5, 'neigh_op_tnl_5')
// (4, 6, 'neigh_op_lft_5')
// (4, 7, 'neigh_op_bnl_5')

wire n388;
// (2, 5, 'neigh_op_tnr_7')
// (2, 6, 'local_g2_7')
// (2, 6, 'lutff_7/in_0')
// (2, 6, 'neigh_op_rgt_7')
// (2, 7, 'neigh_op_bnr_7')
// (3, 5, 'neigh_op_top_7')
// (3, 6, 'lutff_7/out')
// (3, 7, 'neigh_op_bot_7')
// (4, 5, 'local_g2_7')
// (4, 5, 'lutff_0/in_1')
// (4, 5, 'neigh_op_tnl_7')
// (4, 6, 'neigh_op_lft_7')
// (4, 7, 'neigh_op_bnl_7')

reg n389 = 0;
// (2, 5, 'sp4_h_r_4')
// (3, 5, 'local_g0_1')
// (3, 5, 'lutff_0/in_1')
// (3, 5, 'sp4_h_r_17')
// (4, 1, 'local_g3_4')
// (4, 1, 'lutff_3/in_0')
// (4, 1, 'neigh_op_tnr_4')
// (4, 2, 'neigh_op_rgt_4')
// (4, 3, 'local_g0_4')
// (4, 3, 'lutff_7/in_3')
// (4, 3, 'neigh_op_bnr_4')
// (4, 5, 'sp4_h_r_28')
// (5, 1, 'neigh_op_top_4')
// (5, 2, 'lutff_4/out')
// (5, 2, 'sp4_r_v_b_41')
// (5, 3, 'neigh_op_bot_4')
// (5, 3, 'sp4_r_v_b_28')
// (5, 4, 'sp4_r_v_b_17')
// (5, 5, 'sp4_h_r_41')
// (5, 5, 'sp4_r_v_b_4')
// (6, 1, 'neigh_op_tnl_4')
// (6, 1, 'sp4_v_t_41')
// (6, 2, 'neigh_op_lft_4')
// (6, 2, 'sp4_v_b_41')
// (6, 3, 'neigh_op_bnl_4')
// (6, 3, 'sp4_v_b_28')
// (6, 4, 'sp4_v_b_17')
// (6, 5, 'sp4_h_l_41')
// (6, 5, 'sp4_v_b_4')

reg n390 = 0;
// (2, 5, 'sp4_h_r_6')
// (3, 4, 'neigh_op_tnr_7')
// (3, 5, 'local_g3_7')
// (3, 5, 'lutff_6/in_2')
// (3, 5, 'neigh_op_rgt_7')
// (3, 5, 'sp4_h_r_19')
// (3, 6, 'neigh_op_bnr_7')
// (4, 4, 'neigh_op_top_7')
// (4, 5, 'local_g1_7')
// (4, 5, 'lutff_3/in_1')
// (4, 5, 'lutff_7/out')
// (4, 5, 'sp4_h_r_30')
// (4, 6, 'neigh_op_bot_7')
// (5, 4, 'neigh_op_tnl_7')
// (5, 5, 'neigh_op_lft_7')
// (5, 5, 'sp4_h_r_43')
// (5, 6, 'neigh_op_bnl_7')
// (6, 5, 'sp4_h_l_43')
// (6, 5, 'sp4_h_r_6')
// (7, 5, 'local_g0_3')
// (7, 5, 'lutff_6/in_3')
// (7, 5, 'sp4_h_r_19')
// (8, 5, 'sp4_h_r_30')
// (9, 5, 'sp4_h_r_43')
// (10, 5, 'sp4_h_l_43')

wire n391;
// (2, 5, 'sp4_r_v_b_46')
// (2, 6, 'sp4_r_v_b_35')
// (2, 7, 'local_g3_6')
// (2, 7, 'lutff_0/in_3')
// (2, 7, 'lutff_7/in_2')
// (2, 7, 'sp4_r_v_b_22')
// (2, 8, 'sp4_r_v_b_11')
// (2, 9, 'sp4_r_v_b_38')
// (2, 10, 'neigh_op_tnr_7')
// (2, 10, 'sp4_r_v_b_27')
// (2, 11, 'neigh_op_rgt_7')
// (2, 11, 'sp4_r_v_b_14')
// (2, 12, 'neigh_op_bnr_7')
// (2, 12, 'sp4_r_v_b_3')
// (3, 4, 'sp4_v_t_46')
// (3, 5, 'sp4_v_b_46')
// (3, 6, 'sp4_v_b_35')
// (3, 7, 'sp4_v_b_22')
// (3, 8, 'sp4_v_b_11')
// (3, 8, 'sp4_v_t_38')
// (3, 9, 'sp4_v_b_38')
// (3, 10, 'neigh_op_top_7')
// (3, 10, 'sp4_v_b_27')
// (3, 11, 'lutff_7/out')
// (3, 11, 'sp4_v_b_14')
// (3, 12, 'local_g0_7')
// (3, 12, 'lutff_6/in_1')
// (3, 12, 'neigh_op_bot_7')
// (3, 12, 'sp4_v_b_3')
// (4, 10, 'neigh_op_tnl_7')
// (4, 11, 'local_g1_7')
// (4, 11, 'lutff_2/in_2')
// (4, 11, 'neigh_op_lft_7')
// (4, 12, 'neigh_op_bnl_7')

wire n392;
// (2, 6, 'lutff_1/cout')
// (2, 6, 'lutff_2/in_3')

wire n393;
// (2, 6, 'lutff_2/cout')
// (2, 6, 'lutff_3/in_3')

wire n394;
// (2, 6, 'lutff_3/cout')
// (2, 6, 'lutff_4/in_3')

wire n395;
// (2, 6, 'lutff_4/cout')
// (2, 6, 'lutff_5/in_3')

reg n396 = 0;
// (2, 6, 'neigh_op_tnr_0')
// (2, 7, 'neigh_op_rgt_0')
// (2, 8, 'neigh_op_bnr_0')
// (3, 4, 'sp4_r_v_b_36')
// (3, 5, 'sp4_r_v_b_25')
// (3, 6, 'neigh_op_top_0')
// (3, 6, 'sp4_r_v_b_12')
// (3, 7, 'lutff_0/out')
// (3, 7, 'sp4_r_v_b_1')
// (3, 8, 'neigh_op_bot_0')
// (4, 3, 'sp4_v_t_36')
// (4, 4, 'sp4_v_b_36')
// (4, 5, 'local_g2_1')
// (4, 5, 'lutff_5/in_0')
// (4, 5, 'sp4_v_b_25')
// (4, 6, 'neigh_op_tnl_0')
// (4, 6, 'sp4_v_b_12')
// (4, 7, 'neigh_op_lft_0')
// (4, 7, 'sp4_v_b_1')
// (4, 8, 'local_g3_0')
// (4, 8, 'lutff_2/in_1')
// (4, 8, 'lutff_4/in_1')
// (4, 8, 'neigh_op_bnl_0')

wire n397;
// (2, 6, 'neigh_op_tnr_1')
// (2, 7, 'local_g3_1')
// (2, 7, 'lutff_0/in_2')
// (2, 7, 'lutff_2/in_0')
// (2, 7, 'neigh_op_rgt_1')
// (2, 8, 'neigh_op_bnr_1')
// (3, 6, 'neigh_op_top_1')
// (3, 7, 'lutff_1/out')
// (3, 8, 'neigh_op_bot_1')
// (4, 6, 'neigh_op_tnl_1')
// (4, 7, 'neigh_op_lft_1')
// (4, 8, 'neigh_op_bnl_1')

reg n398 = 0;
// (2, 6, 'neigh_op_tnr_2')
// (2, 7, 'neigh_op_rgt_2')
// (2, 7, 'sp4_h_r_9')
// (2, 8, 'neigh_op_bnr_2')
// (3, 6, 'local_g1_2')
// (3, 6, 'lutff_7/in_0')
// (3, 6, 'neigh_op_top_2')
// (3, 7, 'lutff_2/out')
// (3, 7, 'sp4_h_r_20')
// (3, 7, 'sp4_r_v_b_37')
// (3, 8, 'neigh_op_bot_2')
// (3, 8, 'sp4_r_v_b_24')
// (3, 9, 'sp4_r_v_b_13')
// (3, 10, 'sp4_r_v_b_0')
// (4, 6, 'neigh_op_tnl_2')
// (4, 6, 'sp4_v_t_37')
// (4, 7, 'neigh_op_lft_2')
// (4, 7, 'sp4_h_r_33')
// (4, 7, 'sp4_v_b_37')
// (4, 8, 'local_g2_2')
// (4, 8, 'lutff_0/in_2')
// (4, 8, 'lutff_1/in_3')
// (4, 8, 'lutff_5/in_3')
// (4, 8, 'neigh_op_bnl_2')
// (4, 8, 'sp4_v_b_24')
// (4, 9, 'local_g1_5')
// (4, 9, 'lutff_1/in_3')
// (4, 9, 'sp4_v_b_13')
// (4, 10, 'sp4_v_b_0')
// (5, 4, 'sp4_r_v_b_38')
// (5, 5, 'sp4_r_v_b_27')
// (5, 6, 'local_g2_6')
// (5, 6, 'lutff_7/in_1')
// (5, 6, 'sp4_r_v_b_14')
// (5, 7, 'sp4_h_r_44')
// (5, 7, 'sp4_r_v_b_3')
// (6, 3, 'sp4_v_t_38')
// (6, 4, 'sp4_v_b_38')
// (6, 5, 'sp4_v_b_27')
// (6, 6, 'sp4_v_b_14')
// (6, 7, 'sp4_h_l_44')
// (6, 7, 'sp4_v_b_3')

wire n399;
// (2, 6, 'neigh_op_tnr_4')
// (2, 7, 'neigh_op_rgt_4')
// (2, 8, 'neigh_op_bnr_4')
// (3, 6, 'neigh_op_top_4')
// (3, 7, 'lutff_4/out')
// (3, 8, 'neigh_op_bot_4')
// (4, 6, 'local_g2_4')
// (4, 6, 'lutff_5/in_1')
// (4, 6, 'neigh_op_tnl_4')
// (4, 7, 'neigh_op_lft_4')
// (4, 8, 'neigh_op_bnl_4')

reg n400 = 0;
// (2, 6, 'neigh_op_tnr_5')
// (2, 7, 'neigh_op_rgt_5')
// (2, 8, 'neigh_op_bnr_5')
// (3, 6, 'neigh_op_top_5')
// (3, 7, 'lutff_5/out')
// (3, 7, 'sp4_r_v_b_43')
// (3, 8, 'neigh_op_bot_5')
// (3, 8, 'sp4_r_v_b_30')
// (3, 9, 'sp4_r_v_b_19')
// (3, 10, 'sp4_r_v_b_6')
// (4, 6, 'neigh_op_tnl_5')
// (4, 6, 'sp4_v_t_43')
// (4, 7, 'local_g0_5')
// (4, 7, 'lutff_3/in_2')
// (4, 7, 'neigh_op_lft_5')
// (4, 7, 'sp4_v_b_43')
// (4, 8, 'neigh_op_bnl_5')
// (4, 8, 'sp4_v_b_30')
// (4, 9, 'local_g0_3')
// (4, 9, 'lutff_2/in_1')
// (4, 9, 'sp4_v_b_19')
// (4, 10, 'sp4_v_b_6')

reg n401 = 0;
// (2, 6, 'neigh_op_tnr_7')
// (2, 7, 'neigh_op_rgt_7')
// (2, 8, 'neigh_op_bnr_7')
// (3, 5, 'sp4_r_v_b_39')
// (3, 6, 'neigh_op_top_7')
// (3, 6, 'sp4_r_v_b_26')
// (3, 7, 'lutff_7/out')
// (3, 7, 'sp4_r_v_b_15')
// (3, 7, 'sp4_r_v_b_47')
// (3, 8, 'neigh_op_bot_7')
// (3, 8, 'sp4_r_v_b_2')
// (3, 8, 'sp4_r_v_b_34')
// (3, 9, 'sp4_r_v_b_23')
// (3, 10, 'sp4_r_v_b_10')
// (4, 4, 'sp4_v_t_39')
// (4, 5, 'local_g3_7')
// (4, 5, 'lutff_5/in_3')
// (4, 5, 'sp4_v_b_39')
// (4, 6, 'neigh_op_tnl_7')
// (4, 6, 'sp4_v_b_26')
// (4, 6, 'sp4_v_t_47')
// (4, 7, 'neigh_op_lft_7')
// (4, 7, 'sp4_v_b_15')
// (4, 7, 'sp4_v_b_47')
// (4, 8, 'local_g3_7')
// (4, 8, 'lutff_1/in_1')
// (4, 8, 'neigh_op_bnl_7')
// (4, 8, 'sp4_v_b_2')
// (4, 8, 'sp4_v_b_34')
// (4, 9, 'local_g0_7')
// (4, 9, 'lutff_4/in_1')
// (4, 9, 'sp4_v_b_23')
// (4, 10, 'sp4_v_b_10')

wire n402;
// (2, 6, 'sp4_h_r_5')
// (3, 6, 'sp4_h_r_16')
// (4, 5, 'neigh_op_tnr_4')
// (4, 6, 'local_g2_5')
// (4, 6, 'lutff_3/in_2')
// (4, 6, 'lutff_4/in_3')
// (4, 6, 'neigh_op_rgt_4')
// (4, 6, 'sp4_h_r_29')
// (4, 7, 'local_g1_4')
// (4, 7, 'lutff_6/in_3')
// (4, 7, 'neigh_op_bnr_4')
// (5, 5, 'neigh_op_top_4')
// (5, 6, 'lutff_4/out')
// (5, 6, 'sp4_h_r_40')
// (5, 7, 'neigh_op_bot_4')
// (6, 5, 'neigh_op_tnl_4')
// (6, 6, 'neigh_op_lft_4')
// (6, 6, 'sp4_h_l_40')
// (6, 7, 'neigh_op_bnl_4')

wire n403;
// (2, 7, 'neigh_op_tnr_1')
// (2, 8, 'neigh_op_rgt_1')
// (2, 9, 'neigh_op_bnr_1')
// (3, 7, 'neigh_op_top_1')
// (3, 8, 'local_g3_1')
// (3, 8, 'lutff_1/out')
// (3, 8, 'lutff_5/in_1')
// (3, 9, 'neigh_op_bot_1')
// (4, 7, 'neigh_op_tnl_1')
// (4, 8, 'neigh_op_lft_1')
// (4, 9, 'neigh_op_bnl_1')

wire n404;
// (2, 7, 'neigh_op_tnr_2')
// (2, 8, 'neigh_op_rgt_2')
// (2, 9, 'neigh_op_bnr_2')
// (3, 7, 'neigh_op_top_2')
// (3, 8, 'local_g0_2')
// (3, 8, 'lutff_2/out')
// (3, 8, 'lutff_7/in_3')
// (3, 9, 'neigh_op_bot_2')
// (4, 7, 'neigh_op_tnl_2')
// (4, 8, 'neigh_op_lft_2')
// (4, 9, 'neigh_op_bnl_2')

reg n405 = 0;
// (2, 7, 'neigh_op_tnr_3')
// (2, 8, 'neigh_op_rgt_3')
// (2, 9, 'neigh_op_bnr_3')
// (3, 7, 'neigh_op_top_3')
// (3, 8, 'lutff_3/out')
// (3, 9, 'local_g1_3')
// (3, 9, 'lutff_3/in_1')
// (3, 9, 'neigh_op_bot_3')
// (4, 7, 'neigh_op_tnl_3')
// (4, 8, 'neigh_op_lft_3')
// (4, 9, 'neigh_op_bnl_3')

reg n406 = 0;
// (2, 7, 'neigh_op_tnr_4')
// (2, 8, 'neigh_op_rgt_4')
// (2, 9, 'neigh_op_bnr_4')
// (3, 7, 'neigh_op_top_4')
// (3, 8, 'lutff_4/out')
// (3, 9, 'local_g1_4')
// (3, 9, 'lutff_0/in_1')
// (3, 9, 'neigh_op_bot_4')
// (4, 7, 'neigh_op_tnl_4')
// (4, 8, 'neigh_op_lft_4')
// (4, 9, 'local_g2_4')
// (4, 9, 'lutff_7/in_1')
// (4, 9, 'neigh_op_bnl_4')

reg n407 = 0;
// (2, 7, 'neigh_op_tnr_5')
// (2, 8, 'neigh_op_rgt_5')
// (2, 9, 'neigh_op_bnr_5')
// (3, 7, 'neigh_op_top_5')
// (3, 8, 'lutff_5/out')
// (3, 9, 'local_g1_5')
// (3, 9, 'lutff_1/in_1')
// (3, 9, 'neigh_op_bot_5')
// (4, 7, 'neigh_op_tnl_5')
// (4, 8, 'neigh_op_lft_5')
// (4, 9, 'neigh_op_bnl_5')

wire n408;
// (2, 7, 'neigh_op_tnr_6')
// (2, 8, 'neigh_op_rgt_6')
// (2, 9, 'neigh_op_bnr_6')
// (3, 7, 'neigh_op_top_6')
// (3, 8, 'lutff_6/out')
// (3, 9, 'local_g0_6')
// (3, 9, 'lutff_6/in_2')
// (3, 9, 'neigh_op_bot_6')
// (4, 7, 'neigh_op_tnl_6')
// (4, 8, 'neigh_op_lft_6')
// (4, 9, 'neigh_op_bnl_6')

reg n409 = 0;
// (2, 7, 'neigh_op_tnr_7')
// (2, 8, 'neigh_op_rgt_7')
// (2, 9, 'neigh_op_bnr_7')
// (3, 7, 'neigh_op_top_7')
// (3, 8, 'lutff_7/out')
// (3, 9, 'local_g1_7')
// (3, 9, 'lutff_2/in_2')
// (3, 9, 'neigh_op_bot_7')
// (4, 7, 'neigh_op_tnl_7')
// (4, 8, 'neigh_op_lft_7')
// (4, 9, 'neigh_op_bnl_7')

reg n410 = 0;
// (2, 7, 'sp4_h_r_3')
// (3, 4, 'sp4_r_v_b_41')
// (3, 5, 'sp4_r_v_b_28')
// (3, 6, 'local_g3_1')
// (3, 6, 'lutff_1/in_1')
// (3, 6, 'sp4_r_v_b_17')
// (3, 7, 'local_g1_6')
// (3, 7, 'lutff_4/in_3')
// (3, 7, 'sp4_h_r_14')
// (3, 7, 'sp4_r_v_b_4')
// (4, 3, 'sp4_v_t_41')
// (4, 4, 'sp4_v_b_41')
// (4, 5, 'sp4_v_b_28')
// (4, 6, 'neigh_op_tnr_3')
// (4, 6, 'sp4_v_b_17')
// (4, 7, 'neigh_op_rgt_3')
// (4, 7, 'sp4_h_r_11')
// (4, 7, 'sp4_h_r_27')
// (4, 7, 'sp4_v_b_4')
// (4, 8, 'neigh_op_bnr_3')
// (5, 6, 'local_g0_3')
// (5, 6, 'lutff_1/in_2')
// (5, 6, 'neigh_op_top_3')
// (5, 7, 'lutff_3/out')
// (5, 7, 'sp4_h_r_22')
// (5, 7, 'sp4_h_r_38')
// (5, 7, 'sp4_r_v_b_39')
// (5, 8, 'neigh_op_bot_3')
// (5, 8, 'sp4_r_v_b_26')
// (5, 9, 'local_g2_7')
// (5, 9, 'lutff_3/in_2')
// (5, 9, 'sp4_r_v_b_15')
// (5, 10, 'sp4_r_v_b_2')
// (6, 6, 'neigh_op_tnl_3')
// (6, 6, 'sp4_v_t_39')
// (6, 7, 'neigh_op_lft_3')
// (6, 7, 'sp4_h_l_38')
// (6, 7, 'sp4_h_r_35')
// (6, 7, 'sp4_v_b_39')
// (6, 8, 'neigh_op_bnl_3')
// (6, 8, 'sp4_v_b_26')
// (6, 9, 'sp4_v_b_15')
// (6, 10, 'sp4_v_b_2')
// (7, 7, 'sp4_h_r_46')
// (8, 7, 'sp4_h_l_46')

wire n411;
// (2, 8, 'lutff_1/cout')
// (2, 8, 'lutff_2/in_3')

wire n412;
// (2, 8, 'lutff_2/cout')
// (2, 8, 'lutff_3/in_3')

wire n413;
// (2, 8, 'lutff_3/cout')
// (2, 8, 'lutff_4/in_3')

wire n414;
// (2, 8, 'neigh_op_tnr_1')
// (2, 9, 'neigh_op_rgt_1')
// (2, 10, 'neigh_op_bnr_1')
// (3, 8, 'neigh_op_top_1')
// (3, 9, 'local_g2_1')
// (3, 9, 'lutff_1/out')
// (3, 9, 'lutff_6/in_3')
// (3, 10, 'neigh_op_bot_1')
// (4, 8, 'neigh_op_tnl_1')
// (4, 9, 'neigh_op_lft_1')
// (4, 10, 'neigh_op_bnl_1')

wire n415;
// (2, 8, 'neigh_op_tnr_2')
// (2, 9, 'neigh_op_rgt_2')
// (2, 10, 'neigh_op_bnr_2')
// (3, 8, 'neigh_op_top_2')
// (3, 9, 'local_g1_2')
// (3, 9, 'lutff_2/out')
// (3, 9, 'lutff_5/in_2')
// (3, 10, 'neigh_op_bot_2')
// (4, 8, 'neigh_op_tnl_2')
// (4, 9, 'neigh_op_lft_2')
// (4, 10, 'neigh_op_bnl_2')

wire n416;
// (2, 8, 'neigh_op_tnr_3')
// (2, 9, 'neigh_op_rgt_3')
// (2, 10, 'neigh_op_bnr_3')
// (3, 8, 'local_g0_3')
// (3, 8, 'lutff_6/in_3')
// (3, 8, 'neigh_op_top_3')
// (3, 9, 'lutff_3/out')
// (3, 10, 'neigh_op_bot_3')
// (4, 8, 'neigh_op_tnl_3')
// (4, 9, 'neigh_op_lft_3')
// (4, 10, 'neigh_op_bnl_3')

wire n417;
// (2, 8, 'neigh_op_tnr_4')
// (2, 9, 'neigh_op_rgt_4')
// (2, 10, 'neigh_op_bnr_4')
// (3, 8, 'local_g1_4')
// (3, 8, 'lutff_6/in_1')
// (3, 8, 'neigh_op_top_4')
// (3, 9, 'lutff_4/out')
// (3, 10, 'neigh_op_bot_4')
// (4, 8, 'neigh_op_tnl_4')
// (4, 9, 'neigh_op_lft_4')
// (4, 10, 'neigh_op_bnl_4')

wire n418;
// (2, 8, 'neigh_op_tnr_5')
// (2, 9, 'neigh_op_rgt_5')
// (2, 10, 'neigh_op_bnr_5')
// (3, 8, 'neigh_op_top_5')
// (3, 9, 'local_g3_5')
// (3, 9, 'lutff_5/out')
// (3, 9, 'lutff_6/in_0')
// (3, 10, 'neigh_op_bot_5')
// (4, 8, 'neigh_op_tnl_5')
// (4, 9, 'neigh_op_lft_5')
// (4, 10, 'neigh_op_bnl_5')

reg n419 = 0;
// (2, 8, 'neigh_op_tnr_7')
// (2, 9, 'neigh_op_rgt_7')
// (2, 10, 'neigh_op_bnr_7')
// (3, 8, 'neigh_op_top_7')
// (3, 9, 'local_g0_7')
// (3, 9, 'lutff_7/in_0')
// (3, 9, 'lutff_7/out')
// (3, 10, 'local_g1_7')
// (3, 10, 'lutff_4/in_0')
// (3, 10, 'neigh_op_bot_7')
// (4, 8, 'neigh_op_tnl_7')
// (4, 9, 'neigh_op_lft_7')
// (4, 10, 'neigh_op_bnl_7')

wire n420;
// (2, 9, 'lutff_1/cout')
// (2, 9, 'lutff_2/in_3')

wire n421;
// (2, 9, 'lutff_2/cout')
// (2, 9, 'lutff_3/in_3')

reg n422 = 0;
// (2, 9, 'sp4_r_v_b_42')
// (2, 10, 'sp4_r_v_b_31')
// (2, 11, 'sp4_r_v_b_18')
// (2, 12, 'local_g1_7')
// (2, 12, 'lutff_7/in_1')
// (2, 12, 'sp4_r_v_b_7')
// (2, 13, 'sp4_r_v_b_42')
// (2, 14, 'sp4_r_v_b_31')
// (2, 15, 'local_g3_2')
// (2, 15, 'lutff_7/in_2')
// (2, 15, 'sp4_r_v_b_18')
// (2, 16, 'sp4_r_v_b_7')
// (3, 8, 'sp4_v_t_42')
// (3, 9, 'sp4_v_b_42')
// (3, 10, 'sp4_v_b_31')
// (3, 11, 'sp4_v_b_18')
// (3, 12, 'sp4_h_r_7')
// (3, 12, 'sp4_v_b_7')
// (3, 12, 'sp4_v_t_42')
// (3, 13, 'sp4_v_b_42')
// (3, 14, 'sp4_v_b_31')
// (3, 15, 'sp4_v_b_18')
// (3, 16, 'sp4_v_b_7')
// (4, 12, 'sp4_h_r_18')
// (4, 14, 'sp4_r_v_b_43')
// (4, 15, 'sp4_r_v_b_30')
// (4, 16, 'sp4_r_v_b_19')
// (4, 17, 'sp4_r_v_b_6')
// (5, 12, 'sp4_h_r_31')
// (5, 13, 'sp4_h_r_0')
// (5, 13, 'sp4_v_t_43')
// (5, 14, 'sp4_v_b_43')
// (5, 15, 'sp4_v_b_30')
// (5, 16, 'local_g1_3')
// (5, 16, 'lutff_4/in_0')
// (5, 16, 'sp4_v_b_19')
// (5, 17, 'sp4_v_b_6')
// (6, 12, 'sp4_h_r_42')
// (6, 13, 'sp4_h_r_13')
// (7, 12, 'sp4_h_l_42')
// (7, 12, 'sp4_h_r_11')
// (7, 13, 'sp4_h_r_24')
// (8, 12, 'sp4_h_r_22')
// (8, 13, 'sp4_h_r_37')
// (9, 12, 'sp4_h_r_35')
// (9, 13, 'sp4_h_l_37')
// (9, 13, 'sp4_h_r_0')
// (10, 12, 'neigh_op_tnr_4')
// (10, 12, 'sp4_h_r_46')
// (10, 13, 'neigh_op_rgt_4')
// (10, 13, 'sp4_h_r_13')
// (10, 13, 'sp4_r_v_b_40')
// (10, 14, 'neigh_op_bnr_4')
// (10, 14, 'sp4_r_v_b_29')
// (10, 15, 'sp4_r_v_b_16')
// (10, 16, 'sp4_r_v_b_5')
// (11, 12, 'neigh_op_top_4')
// (11, 12, 'sp4_h_l_46')
// (11, 12, 'sp4_v_t_40')
// (11, 13, 'lutff_4/out')
// (11, 13, 'sp4_h_r_24')
// (11, 13, 'sp4_v_b_40')
// (11, 14, 'neigh_op_bot_4')
// (11, 14, 'sp4_v_b_29')
// (11, 15, 'sp4_v_b_16')
// (11, 16, 'local_g0_5')
// (11, 16, 'lutff_4/in_1')
// (11, 16, 'sp4_v_b_5')
// (12, 12, 'neigh_op_tnl_4')
// (12, 13, 'neigh_op_lft_4')
// (12, 13, 'sp4_h_r_37')
// (12, 14, 'neigh_op_bnl_4')
// (13, 13, 'sp4_h_l_37')

wire n423;
// (2, 10, 'local_g3_6')
// (2, 10, 'lutff_5/in_2')
// (2, 10, 'neigh_op_tnr_6')
// (2, 11, 'local_g3_6')
// (2, 11, 'lutff_7/in_0')
// (2, 11, 'neigh_op_rgt_6')
// (2, 11, 'sp4_h_r_1')
// (2, 12, 'local_g0_6')
// (2, 12, 'lutff_5/in_3')
// (2, 12, 'neigh_op_bnr_6')
// (3, 10, 'neigh_op_top_6')
// (3, 10, 'sp4_r_v_b_40')
// (3, 11, 'lutff_6/out')
// (3, 11, 'sp4_h_r_12')
// (3, 11, 'sp4_r_v_b_29')
// (3, 12, 'neigh_op_bot_6')
// (3, 12, 'sp4_r_v_b_16')
// (3, 13, 'sp4_r_v_b_5')
// (4, 9, 'sp4_h_r_5')
// (4, 9, 'sp4_v_t_40')
// (4, 10, 'neigh_op_tnl_6')
// (4, 10, 'sp4_v_b_40')
// (4, 11, 'neigh_op_lft_6')
// (4, 11, 'sp4_h_r_25')
// (4, 11, 'sp4_v_b_29')
// (4, 12, 'neigh_op_bnl_6')
// (4, 12, 'sp4_v_b_16')
// (4, 13, 'sp4_v_b_5')
// (5, 9, 'sp4_h_r_16')
// (5, 11, 'sp4_h_r_36')
// (6, 9, 'sp4_h_r_29')
// (6, 11, 'sp4_h_l_36')
// (6, 11, 'sp4_h_r_4')
// (7, 9, 'sp4_h_r_40')
// (7, 11, 'sp4_h_r_17')
// (8, 9, 'sp4_h_l_40')
// (8, 9, 'sp4_h_r_8')
// (8, 11, 'sp4_h_r_28')
// (9, 9, 'sp4_h_r_21')
// (9, 11, 'local_g3_1')
// (9, 11, 'lutff_6/in_2')
// (9, 11, 'sp4_h_r_41')
// (10, 9, 'sp4_h_r_32')
// (10, 11, 'sp4_h_l_41')
// (10, 11, 'sp4_h_r_7')
// (11, 9, 'sp4_h_r_45')
// (11, 11, 'sp4_h_r_18')
// (12, 9, 'local_g0_3')
// (12, 9, 'lutff_6/in_3')
// (12, 9, 'sp4_h_l_45')
// (12, 9, 'sp4_h_r_11')
// (12, 11, 'sp4_h_r_31')
// (13, 9, 'sp4_h_r_22')
// (13, 11, 'sp4_h_r_42')
// (14, 9, 'sp4_h_r_35')
// (14, 11, 'local_g0_7')
// (14, 11, 'lutff_6/in_3')
// (14, 11, 'sp4_h_l_42')
// (14, 11, 'sp4_h_r_7')
// (15, 9, 'sp4_h_r_46')
// (15, 11, 'sp4_h_r_18')
// (16, 9, 'sp4_h_l_46')
// (16, 11, 'sp4_h_r_31')
// (17, 11, 'sp4_h_r_42')
// (18, 11, 'sp4_h_l_42')

wire n424;
// (2, 10, 'neigh_op_tnr_1')
// (2, 10, 'sp4_r_v_b_47')
// (2, 11, 'neigh_op_rgt_1')
// (2, 11, 'sp4_r_v_b_34')
// (2, 12, 'neigh_op_bnr_1')
// (2, 12, 'sp4_r_v_b_23')
// (2, 13, 'sp4_r_v_b_10')
// (3, 9, 'sp4_v_t_47')
// (3, 10, 'neigh_op_top_1')
// (3, 10, 'sp4_r_v_b_46')
// (3, 10, 'sp4_v_b_47')
// (3, 11, 'lutff_1/out')
// (3, 11, 'sp4_r_v_b_35')
// (3, 11, 'sp4_v_b_34')
// (3, 12, 'neigh_op_bot_1')
// (3, 12, 'sp4_r_v_b_22')
// (3, 12, 'sp4_v_b_23')
// (3, 13, 'local_g1_2')
// (3, 13, 'lutff_2/in_1')
// (3, 13, 'sp4_r_v_b_11')
// (3, 13, 'sp4_v_b_10')
// (4, 9, 'sp4_v_t_46')
// (4, 10, 'neigh_op_tnl_1')
// (4, 10, 'sp4_v_b_46')
// (4, 11, 'neigh_op_lft_1')
// (4, 11, 'sp4_v_b_35')
// (4, 12, 'neigh_op_bnl_1')
// (4, 12, 'sp4_v_b_22')
// (4, 13, 'local_g0_3')
// (4, 13, 'lutff_1/in_2')
// (4, 13, 'sp4_v_b_11')

reg n425 = 0;
// (2, 10, 'neigh_op_tnr_2')
// (2, 11, 'neigh_op_rgt_2')
// (2, 12, 'neigh_op_bnr_2')
// (3, 10, 'neigh_op_top_2')
// (3, 11, 'lutff_2/out')
// (3, 12, 'local_g1_2')
// (3, 12, 'lutff_3/in_0')
// (3, 12, 'neigh_op_bot_2')
// (4, 10, 'neigh_op_tnl_2')
// (4, 11, 'neigh_op_lft_2')
// (4, 12, 'neigh_op_bnl_2')

reg n426 = 0;
// (2, 10, 'sp4_r_v_b_37')
// (2, 11, 'sp4_r_v_b_24')
// (2, 12, 'local_g2_5')
// (2, 12, 'lutff_7/in_0')
// (2, 12, 'sp4_r_v_b_13')
// (2, 13, 'sp4_r_v_b_0')
// (3, 9, 'sp4_v_t_37')
// (3, 10, 'sp4_v_b_37')
// (3, 11, 'sp4_v_b_24')
// (3, 12, 'sp4_v_b_13')
// (3, 13, 'sp4_h_r_0')
// (3, 13, 'sp4_v_b_0')
// (4, 13, 'sp4_h_r_13')
// (5, 13, 'sp4_h_r_24')
// (6, 13, 'sp4_h_r_37')
// (7, 13, 'sp4_h_l_37')
// (7, 13, 'sp4_h_r_0')
// (8, 13, 'sp4_h_r_13')
// (9, 13, 'sp4_h_r_24')
// (10, 13, 'sp4_h_r_37')
// (10, 14, 'sp4_r_v_b_43')
// (10, 15, 'sp4_r_v_b_30')
// (10, 16, 'sp4_r_v_b_19')
// (10, 17, 'sp4_r_v_b_6')
// (10, 18, 'sp4_r_v_b_43')
// (10, 19, 'sp4_r_v_b_30')
// (10, 20, 'neigh_op_tnr_3')
// (10, 20, 'sp4_r_v_b_19')
// (10, 21, 'neigh_op_rgt_3')
// (10, 21, 'sp4_r_v_b_6')
// (10, 22, 'neigh_op_bnr_3')
// (11, 13, 'sp4_h_l_37')
// (11, 13, 'sp4_v_t_43')
// (11, 14, 'sp4_v_b_43')
// (11, 15, 'sp4_v_b_30')
// (11, 16, 'sp4_v_b_19')
// (11, 17, 'sp4_v_b_6')
// (11, 17, 'sp4_v_t_43')
// (11, 18, 'sp4_v_b_43')
// (11, 19, 'local_g2_6')
// (11, 19, 'lutff_5/in_3')
// (11, 19, 'sp4_v_b_30')
// (11, 20, 'neigh_op_top_3')
// (11, 20, 'sp4_v_b_19')
// (11, 21, 'local_g3_3')
// (11, 21, 'lutff_3/in_3')
// (11, 21, 'lutff_3/out')
// (11, 21, 'sp4_v_b_6')
// (11, 22, 'neigh_op_bot_3')
// (12, 20, 'neigh_op_tnl_3')
// (12, 21, 'neigh_op_lft_3')
// (12, 22, 'neigh_op_bnl_3')

wire n427;
// (2, 11, 'local_g2_4')
// (2, 11, 'lutff_2/in_2')
// (2, 11, 'neigh_op_tnr_4')
// (2, 12, 'neigh_op_rgt_4')
// (2, 13, 'neigh_op_bnr_4')
// (3, 11, 'neigh_op_top_4')
// (3, 12, 'lutff_4/out')
// (3, 13, 'neigh_op_bot_4')
// (4, 11, 'neigh_op_tnl_4')
// (4, 12, 'neigh_op_lft_4')
// (4, 13, 'neigh_op_bnl_4')

wire n428;
// (2, 11, 'local_g2_5')
// (2, 11, 'lutff_2/in_3')
// (2, 11, 'neigh_op_tnr_5')
// (2, 12, 'neigh_op_rgt_5')
// (2, 13, 'neigh_op_bnr_5')
// (3, 11, 'neigh_op_top_5')
// (3, 12, 'lutff_5/out')
// (3, 13, 'neigh_op_bot_5')
// (4, 11, 'neigh_op_tnl_5')
// (4, 12, 'neigh_op_lft_5')
// (4, 13, 'neigh_op_bnl_5')

wire n429;
// (2, 11, 'local_g2_6')
// (2, 11, 'lutff_2/in_0')
// (2, 11, 'neigh_op_tnr_6')
// (2, 12, 'neigh_op_rgt_6')
// (2, 13, 'neigh_op_bnr_6')
// (3, 11, 'neigh_op_top_6')
// (3, 12, 'lutff_6/out')
// (3, 13, 'neigh_op_bot_6')
// (4, 11, 'neigh_op_tnl_6')
// (4, 12, 'neigh_op_lft_6')
// (4, 13, 'neigh_op_bnl_6')

wire n430;
// (2, 11, 'neigh_op_tnr_0')
// (2, 12, 'neigh_op_rgt_0')
// (2, 13, 'neigh_op_bnr_0')
// (3, 11, 'neigh_op_top_0')
// (3, 12, 'lutff_0/out')
// (3, 13, 'local_g0_0')
// (3, 13, 'lutff_1/in_1')
// (3, 13, 'neigh_op_bot_0')
// (4, 11, 'neigh_op_tnl_0')
// (4, 12, 'neigh_op_lft_0')
// (4, 13, 'local_g2_0')
// (4, 13, 'lutff_0/in_2')
// (4, 13, 'neigh_op_bnl_0')

wire n431;
// (2, 11, 'neigh_op_tnr_1')
// (2, 12, 'neigh_op_rgt_1')
// (2, 13, 'local_g1_1')
// (2, 13, 'lutff_2/in_2')
// (2, 13, 'neigh_op_bnr_1')
// (3, 11, 'neigh_op_top_1')
// (3, 12, 'lutff_1/out')
// (3, 13, 'neigh_op_bot_1')
// (4, 11, 'neigh_op_tnl_1')
// (4, 12, 'neigh_op_lft_1')
// (4, 13, 'neigh_op_bnl_1')

wire n432;
// (2, 11, 'neigh_op_tnr_2')
// (2, 12, 'neigh_op_rgt_2')
// (2, 13, 'local_g0_2')
// (2, 13, 'lutff_global/cen')
// (2, 13, 'neigh_op_bnr_2')
// (3, 11, 'neigh_op_top_2')
// (3, 12, 'lutff_2/out')
// (3, 13, 'neigh_op_bot_2')
// (4, 11, 'neigh_op_tnl_2')
// (4, 12, 'local_g0_2')
// (4, 12, 'lutff_global/cen')
// (4, 12, 'neigh_op_lft_2')
// (4, 13, 'neigh_op_bnl_2')

wire n433;
// (2, 12, 'neigh_op_tnr_7')
// (2, 13, 'neigh_op_rgt_7')
// (2, 14, 'neigh_op_bnr_7')
// (3, 12, 'neigh_op_top_7')
// (3, 13, 'local_g2_7')
// (3, 13, 'lutff_3/in_2')
// (3, 13, 'lutff_7/out')
// (3, 14, 'local_g1_7')
// (3, 14, 'lutff_0/in_2')
// (3, 14, 'neigh_op_bot_7')
// (4, 12, 'neigh_op_tnl_7')
// (4, 13, 'local_g1_7')
// (4, 13, 'lutff_2/in_2')
// (4, 13, 'neigh_op_lft_7')
// (4, 14, 'neigh_op_bnl_7')

wire n434;
// (2, 12, 'sp4_r_v_b_36')
// (2, 13, 'sp4_r_v_b_25')
// (2, 14, 'neigh_op_tnr_4')
// (2, 14, 'sp4_r_v_b_12')
// (2, 15, 'neigh_op_rgt_4')
// (2, 15, 'sp4_r_v_b_1')
// (2, 16, 'neigh_op_bnr_4')
// (3, 11, 'sp4_v_t_36')
// (3, 12, 'local_g2_4')
// (3, 12, 'lutff_1/in_1')
// (3, 12, 'sp4_r_v_b_44')
// (3, 12, 'sp4_v_b_36')
// (3, 13, 'sp4_r_v_b_33')
// (3, 13, 'sp4_v_b_25')
// (3, 14, 'neigh_op_top_4')
// (3, 14, 'sp4_r_v_b_20')
// (3, 14, 'sp4_v_b_12')
// (3, 15, 'lutff_4/out')
// (3, 15, 'sp4_h_r_8')
// (3, 15, 'sp4_r_v_b_9')
// (3, 15, 'sp4_v_b_1')
// (3, 16, 'neigh_op_bot_4')
// (4, 11, 'sp4_v_t_44')
// (4, 12, 'sp4_v_b_44')
// (4, 13, 'local_g2_1')
// (4, 13, 'lutff_6/in_1')
// (4, 13, 'sp4_v_b_33')
// (4, 14, 'neigh_op_tnl_4')
// (4, 14, 'sp4_v_b_20')
// (4, 15, 'neigh_op_lft_4')
// (4, 15, 'sp4_h_r_21')
// (4, 15, 'sp4_v_b_9')
// (4, 16, 'local_g3_4')
// (4, 16, 'lutff_5/in_0')
// (4, 16, 'lutff_6/in_1')
// (4, 16, 'neigh_op_bnl_4')
// (5, 15, 'sp4_h_r_32')
// (6, 15, 'sp4_h_r_45')
// (7, 15, 'sp4_h_l_45')

wire n435;
// (2, 13, 'local_g2_4')
// (2, 13, 'lutff_6/in_0')
// (2, 13, 'sp4_r_v_b_36')
// (2, 14, 'neigh_op_tnr_6')
// (2, 14, 'sp4_r_v_b_25')
// (2, 15, 'neigh_op_rgt_6')
// (2, 15, 'sp4_r_v_b_12')
// (2, 16, 'neigh_op_bnr_6')
// (2, 16, 'sp4_r_v_b_1')
// (3, 12, 'sp4_v_t_36')
// (3, 13, 'sp4_v_b_36')
// (3, 14, 'neigh_op_top_6')
// (3, 14, 'sp4_v_b_25')
// (3, 15, 'local_g0_6')
// (3, 15, 'lutff_3/in_3')
// (3, 15, 'lutff_6/out')
// (3, 15, 'sp4_v_b_12')
// (3, 16, 'neigh_op_bot_6')
// (3, 16, 'sp4_v_b_1')
// (4, 14, 'neigh_op_tnl_6')
// (4, 15, 'neigh_op_lft_6')
// (4, 16, 'neigh_op_bnl_6')

wire n436;
// (2, 13, 'neigh_op_tnr_3')
// (2, 14, 'neigh_op_rgt_3')
// (2, 15, 'neigh_op_bnr_3')
// (3, 13, 'neigh_op_top_3')
// (3, 14, 'lutff_3/out')
// (3, 15, 'neigh_op_bot_3')
// (4, 13, 'neigh_op_tnl_3')
// (4, 14, 'local_g1_3')
// (4, 14, 'lutff_3/in_1')
// (4, 14, 'neigh_op_lft_3')
// (4, 15, 'neigh_op_bnl_3')

reg n437 = 0;
// (2, 14, 'local_g2_5')
// (2, 14, 'lutff_3/in_0')
// (2, 14, 'sp4_r_v_b_37')
// (2, 15, 'sp4_r_v_b_24')
// (2, 16, 'sp4_r_v_b_13')
// (2, 17, 'sp4_r_v_b_0')
// (2, 18, 'sp4_r_v_b_41')
// (2, 19, 'sp4_r_v_b_28')
// (2, 20, 'neigh_op_tnr_2')
// (2, 20, 'sp4_r_v_b_17')
// (2, 21, 'neigh_op_rgt_2')
// (2, 21, 'sp4_h_r_9')
// (2, 21, 'sp4_r_v_b_4')
// (2, 22, 'neigh_op_bnr_2')
// (3, 13, 'sp4_v_t_37')
// (3, 14, 'sp4_v_b_37')
// (3, 15, 'sp4_v_b_24')
// (3, 16, 'sp4_v_b_13')
// (3, 17, 'sp4_v_b_0')
// (3, 17, 'sp4_v_t_41')
// (3, 18, 'sp4_v_b_41')
// (3, 19, 'sp4_r_v_b_45')
// (3, 19, 'sp4_v_b_28')
// (3, 20, 'neigh_op_top_2')
// (3, 20, 'sp4_r_v_b_32')
// (3, 20, 'sp4_v_b_17')
// (3, 21, 'local_g3_2')
// (3, 21, 'lutff_2/out')
// (3, 21, 'lutff_3/in_0')
// (3, 21, 'sp4_h_r_20')
// (3, 21, 'sp4_h_r_4')
// (3, 21, 'sp4_r_v_b_21')
// (3, 21, 'sp4_v_b_4')
// (3, 22, 'neigh_op_bot_2')
// (3, 22, 'sp4_r_v_b_8')
// (4, 18, 'sp4_v_t_45')
// (4, 19, 'sp4_v_b_45')
// (4, 20, 'neigh_op_tnl_2')
// (4, 20, 'sp4_v_b_32')
// (4, 21, 'neigh_op_lft_2')
// (4, 21, 'sp4_h_r_17')
// (4, 21, 'sp4_h_r_33')
// (4, 21, 'sp4_v_b_21')
// (4, 22, 'neigh_op_bnl_2')
// (4, 22, 'sp4_h_r_2')
// (4, 22, 'sp4_v_b_8')
// (5, 21, 'sp4_h_r_28')
// (5, 21, 'sp4_h_r_44')
// (5, 22, 'sp4_h_r_15')
// (6, 21, 'sp4_h_l_44')
// (6, 21, 'sp4_h_r_41')
// (6, 21, 'sp4_h_r_9')
// (6, 22, 'sp4_h_r_26')
// (7, 21, 'local_g1_7')
// (7, 21, 'lutff_2/in_2')
// (7, 21, 'sp4_h_l_41')
// (7, 21, 'sp4_h_r_20')
// (7, 21, 'sp4_h_r_4')
// (7, 21, 'sp4_h_r_7')
// (7, 22, 'sp4_h_r_39')
// (8, 21, 'local_g0_1')
// (8, 21, 'local_g3_1')
// (8, 21, 'lutff_0/in_1')
// (8, 21, 'lutff_2/in_2')
// (8, 21, 'sp4_h_r_17')
// (8, 21, 'sp4_h_r_18')
// (8, 21, 'sp4_h_r_33')
// (8, 22, 'local_g0_5')
// (8, 22, 'lutff_0/in_1')
// (8, 22, 'lutff_3/in_2')
// (8, 22, 'lutff_7/in_0')
// (8, 22, 'sp4_h_l_39')
// (8, 22, 'sp4_h_r_10')
// (8, 22, 'sp4_h_r_5')
// (9, 21, 'local_g2_4')
// (9, 21, 'local_g3_4')
// (9, 21, 'lutff_2/in_0')
// (9, 21, 'lutff_3/in_0')
// (9, 21, 'lutff_6/in_2')
// (9, 21, 'sp4_h_r_28')
// (9, 21, 'sp4_h_r_31')
// (9, 21, 'sp4_h_r_44')
// (9, 22, 'local_g0_0')
// (9, 22, 'local_g1_7')
// (9, 22, 'lutff_6/in_2')
// (9, 22, 'lutff_7/in_3')
// (9, 22, 'sp4_h_r_16')
// (9, 22, 'sp4_h_r_23')
// (10, 21, 'sp4_h_l_44')
// (10, 21, 'sp4_h_r_41')
// (10, 21, 'sp4_h_r_42')
// (10, 22, 'sp4_h_r_29')
// (10, 22, 'sp4_h_r_34')
// (11, 21, 'sp4_h_l_41')
// (11, 21, 'sp4_h_l_42')
// (11, 22, 'sp4_h_r_40')
// (11, 22, 'sp4_h_r_47')
// (12, 22, 'sp4_h_l_40')
// (12, 22, 'sp4_h_l_47')

reg n438 = 0;
// (2, 14, 'neigh_op_tnr_0')
// (2, 15, 'neigh_op_rgt_0')
// (2, 16, 'neigh_op_bnr_0')
// (3, 14, 'neigh_op_top_0')
// (3, 15, 'local_g2_0')
// (3, 15, 'lutff_0/in_2')
// (3, 15, 'lutff_0/out')
// (3, 15, 'lutff_2/in_2')
// (3, 16, 'neigh_op_bot_0')
// (4, 14, 'neigh_op_tnl_0')
// (4, 15, 'neigh_op_lft_0')
// (4, 16, 'neigh_op_bnl_0')

wire n439;
// (2, 14, 'neigh_op_tnr_1')
// (2, 15, 'neigh_op_rgt_1')
// (2, 15, 'sp4_h_r_7')
// (2, 16, 'neigh_op_bnr_1')
// (3, 14, 'neigh_op_top_1')
// (3, 15, 'lutff_1/out')
// (3, 15, 'sp4_h_r_18')
// (3, 16, 'neigh_op_bot_1')
// (4, 14, 'local_g2_1')
// (4, 14, 'lutff_5/in_2')
// (4, 14, 'neigh_op_tnl_1')
// (4, 15, 'neigh_op_lft_1')
// (4, 15, 'sp4_h_r_31')
// (4, 16, 'neigh_op_bnl_1')
// (5, 12, 'sp4_r_v_b_36')
// (5, 13, 'sp4_r_v_b_25')
// (5, 14, 'local_g2_4')
// (5, 14, 'lutff_0/in_2')
// (5, 14, 'sp4_r_v_b_12')
// (5, 15, 'sp4_h_r_42')
// (5, 15, 'sp4_r_v_b_1')
// (6, 11, 'sp4_v_t_36')
// (6, 12, 'sp4_v_b_36')
// (6, 13, 'sp4_v_b_25')
// (6, 14, 'sp4_v_b_12')
// (6, 15, 'sp4_h_l_42')
// (6, 15, 'sp4_v_b_1')

wire n440;
// (2, 14, 'neigh_op_tnr_2')
// (2, 15, 'neigh_op_rgt_2')
// (2, 16, 'neigh_op_bnr_2')
// (3, 12, 'sp4_r_v_b_40')
// (3, 13, 'sp4_r_v_b_29')
// (3, 14, 'neigh_op_top_2')
// (3, 14, 'sp4_r_v_b_16')
// (3, 15, 'lutff_2/out')
// (3, 15, 'sp4_r_v_b_5')
// (3, 16, 'neigh_op_bot_2')
// (4, 11, 'sp4_v_t_40')
// (4, 12, 'sp4_v_b_40')
// (4, 13, 'local_g3_5')
// (4, 13, 'lutff_7/in_3')
// (4, 13, 'sp4_v_b_29')
// (4, 14, 'neigh_op_tnl_2')
// (4, 14, 'sp4_v_b_16')
// (4, 15, 'neigh_op_lft_2')
// (4, 15, 'sp4_v_b_5')
// (4, 16, 'neigh_op_bnl_2')

wire n441;
// (2, 14, 'neigh_op_tnr_3')
// (2, 15, 'neigh_op_rgt_3')
// (2, 16, 'neigh_op_bnr_3')
// (3, 14, 'neigh_op_top_3')
// (3, 15, 'lutff_3/out')
// (3, 15, 'sp4_h_r_6')
// (3, 16, 'neigh_op_bot_3')
// (4, 14, 'neigh_op_tnl_3')
// (4, 15, 'neigh_op_lft_3')
// (4, 15, 'sp4_h_r_19')
// (4, 16, 'neigh_op_bnl_3')
// (5, 15, 'local_g3_6')
// (5, 15, 'lutff_4/in_3')
// (5, 15, 'sp4_h_r_30')
// (6, 15, 'sp4_h_r_43')
// (7, 15, 'sp4_h_l_43')

reg n442 = 0;
// (2, 14, 'neigh_op_tnr_5')
// (2, 15, 'neigh_op_rgt_5')
// (2, 16, 'neigh_op_bnr_5')
// (3, 14, 'neigh_op_top_5')
// (3, 15, 'local_g3_5')
// (3, 15, 'lutff_2/in_0')
// (3, 15, 'lutff_5/in_3')
// (3, 15, 'lutff_5/out')
// (3, 16, 'neigh_op_bot_5')
// (4, 14, 'neigh_op_tnl_5')
// (4, 15, 'neigh_op_lft_5')
// (4, 16, 'neigh_op_bnl_5')

wire n443;
// (2, 14, 'neigh_op_tnr_7')
// (2, 15, 'local_g3_7')
// (2, 15, 'lutff_6/in_0')
// (2, 15, 'neigh_op_rgt_7')
// (2, 16, 'neigh_op_bnr_7')
// (3, 14, 'neigh_op_top_7')
// (3, 15, 'lutff_7/out')
// (3, 15, 'sp4_r_v_b_47')
// (3, 16, 'neigh_op_bot_7')
// (3, 16, 'sp4_r_v_b_34')
// (3, 17, 'sp4_r_v_b_23')
// (3, 18, 'local_g2_2')
// (3, 18, 'lutff_7/in_1')
// (3, 18, 'sp4_r_v_b_10')
// (4, 14, 'local_g3_7')
// (4, 14, 'lutff_2/in_0')
// (4, 14, 'neigh_op_tnl_7')
// (4, 14, 'sp4_v_t_47')
// (4, 15, 'local_g0_7')
// (4, 15, 'lutff_3/in_0')
// (4, 15, 'neigh_op_lft_7')
// (4, 15, 'sp4_v_b_47')
// (4, 16, 'neigh_op_bnl_7')
// (4, 16, 'sp4_v_b_34')
// (4, 17, 'sp4_v_b_23')
// (4, 18, 'sp4_v_b_10')

wire n444;
// (2, 14, 'sp4_h_r_6')
// (3, 13, 'local_g0_2')
// (3, 13, 'lutff_4/in_2')
// (3, 13, 'sp4_h_r_10')
// (3, 14, 'local_g0_3')
// (3, 14, 'lutff_1/in_2')
// (3, 14, 'sp4_h_r_19')
// (4, 12, 'neigh_op_tnr_1')
// (4, 13, 'local_g3_1')
// (4, 13, 'lutff_3/in_1')
// (4, 13, 'neigh_op_rgt_1')
// (4, 13, 'sp4_h_r_23')
// (4, 14, 'neigh_op_bnr_1')
// (4, 14, 'sp4_h_r_30')
// (5, 11, 'sp4_r_v_b_43')
// (5, 12, 'neigh_op_top_1')
// (5, 12, 'sp4_r_v_b_30')
// (5, 13, 'lutff_1/out')
// (5, 13, 'sp4_h_r_34')
// (5, 13, 'sp4_r_v_b_19')
// (5, 14, 'neigh_op_bot_1')
// (5, 14, 'sp4_h_r_43')
// (5, 14, 'sp4_r_v_b_6')
// (6, 10, 'sp4_v_t_43')
// (6, 11, 'sp4_v_b_43')
// (6, 12, 'neigh_op_tnl_1')
// (6, 12, 'sp4_v_b_30')
// (6, 13, 'neigh_op_lft_1')
// (6, 13, 'sp4_h_r_47')
// (6, 13, 'sp4_v_b_19')
// (6, 14, 'neigh_op_bnl_1')
// (6, 14, 'sp4_h_l_43')
// (6, 14, 'sp4_v_b_6')
// (7, 13, 'sp4_h_l_47')

reg n445 = 0;
// (2, 15, 'neigh_op_tnr_0')
// (2, 16, 'neigh_op_rgt_0')
// (2, 17, 'neigh_op_bnr_0')
// (3, 13, 'sp4_r_v_b_36')
// (3, 14, 'sp4_r_v_b_25')
// (3, 15, 'neigh_op_top_0')
// (3, 15, 'sp4_r_v_b_12')
// (3, 16, 'local_g1_0')
// (3, 16, 'lutff_0/in_3')
// (3, 16, 'lutff_0/out')
// (3, 16, 'sp4_r_v_b_1')
// (3, 17, 'neigh_op_bot_0')
// (4, 12, 'sp4_v_t_36')
// (4, 13, 'local_g3_4')
// (4, 13, 'lutff_7/in_0')
// (4, 13, 'sp4_v_b_36')
// (4, 14, 'sp4_v_b_25')
// (4, 15, 'neigh_op_tnl_0')
// (4, 15, 'sp4_v_b_12')
// (4, 16, 'neigh_op_lft_0')
// (4, 16, 'sp4_v_b_1')
// (4, 17, 'neigh_op_bnl_0')

reg n446 = 0;
// (2, 15, 'neigh_op_tnr_1')
// (2, 16, 'neigh_op_rgt_1')
// (2, 17, 'neigh_op_bnr_1')
// (3, 11, 'sp4_r_v_b_42')
// (3, 12, 'sp4_r_v_b_31')
// (3, 13, 'sp4_r_v_b_18')
// (3, 14, 'sp4_r_v_b_7')
// (3, 15, 'local_g1_1')
// (3, 15, 'lutff_4/in_2')
// (3, 15, 'lutff_6/in_2')
// (3, 15, 'neigh_op_top_1')
// (3, 15, 'sp4_r_v_b_46')
// (3, 16, 'local_g0_1')
// (3, 16, 'lutff_1/in_0')
// (3, 16, 'lutff_1/out')
// (3, 16, 'sp4_r_v_b_35')
// (3, 17, 'neigh_op_bot_1')
// (3, 17, 'sp4_r_v_b_22')
// (3, 18, 'sp4_r_v_b_11')
// (4, 10, 'sp4_v_t_42')
// (4, 11, 'local_g2_2')
// (4, 11, 'lutff_7/in_3')
// (4, 11, 'sp4_v_b_42')
// (4, 12, 'sp4_v_b_31')
// (4, 13, 'sp4_v_b_18')
// (4, 14, 'sp4_v_b_7')
// (4, 14, 'sp4_v_t_46')
// (4, 15, 'local_g2_1')
// (4, 15, 'lutff_0/in_3')
// (4, 15, 'neigh_op_tnl_1')
// (4, 15, 'sp4_v_b_46')
// (4, 16, 'neigh_op_lft_1')
// (4, 16, 'sp4_v_b_35')
// (4, 17, 'local_g3_1')
// (4, 17, 'lutff_3/in_3')
// (4, 17, 'neigh_op_bnl_1')
// (4, 17, 'sp4_v_b_22')
// (4, 18, 'sp4_v_b_11')

wire n447;
// (2, 15, 'neigh_op_tnr_2')
// (2, 16, 'neigh_op_rgt_2')
// (2, 17, 'neigh_op_bnr_2')
// (3, 15, 'local_g0_2')
// (3, 15, 'lutff_7/in_3')
// (3, 15, 'neigh_op_top_2')
// (3, 16, 'lutff_2/out')
// (3, 17, 'neigh_op_bot_2')
// (4, 15, 'neigh_op_tnl_2')
// (4, 16, 'neigh_op_lft_2')
// (4, 17, 'neigh_op_bnl_2')

wire n448;
// (2, 15, 'neigh_op_tnr_4')
// (2, 16, 'neigh_op_rgt_4')
// (2, 17, 'neigh_op_bnr_4')
// (3, 15, 'neigh_op_top_4')
// (3, 16, 'lutff_4/out')
// (3, 16, 'sp4_h_r_8')
// (3, 17, 'neigh_op_bot_4')
// (4, 15, 'neigh_op_tnl_4')
// (4, 16, 'local_g1_4')
// (4, 16, 'lutff_7/in_2')
// (4, 16, 'neigh_op_lft_4')
// (4, 16, 'sp4_h_r_21')
// (4, 17, 'local_g2_4')
// (4, 17, 'lutff_0/in_2')
// (4, 17, 'lutff_5/in_1')
// (4, 17, 'lutff_6/in_0')
// (4, 17, 'lutff_7/in_3')
// (4, 17, 'neigh_op_bnl_4')
// (5, 16, 'sp4_h_r_32')
// (6, 16, 'sp4_h_r_45')
// (6, 17, 'sp4_r_v_b_45')
// (6, 18, 'sp4_r_v_b_32')
// (6, 19, 'sp4_r_v_b_21')
// (6, 20, 'sp4_r_v_b_8')
// (7, 16, 'sp4_h_l_45')
// (7, 16, 'sp4_v_t_45')
// (7, 17, 'local_g3_5')
// (7, 17, 'lutff_1/in_3')
// (7, 17, 'lutff_2/in_0')
// (7, 17, 'lutff_4/in_2')
// (7, 17, 'lutff_5/in_3')
// (7, 17, 'sp4_v_b_45')
// (7, 18, 'sp4_v_b_32')
// (7, 19, 'sp4_v_b_21')
// (7, 20, 'sp4_v_b_8')

wire n449;
// (2, 15, 'neigh_op_tnr_7')
// (2, 16, 'neigh_op_rgt_7')
// (2, 16, 'sp4_h_r_3')
// (2, 17, 'neigh_op_bnr_7')
// (3, 11, 'sp4_r_v_b_47')
// (3, 12, 'sp4_r_v_b_34')
// (3, 13, 'sp4_r_v_b_23')
// (3, 14, 'sp4_r_v_b_10')
// (3, 15, 'neigh_op_top_7')
// (3, 15, 'sp4_r_v_b_42')
// (3, 16, 'local_g2_7')
// (3, 16, 'lutff_0/in_1')
// (3, 16, 'lutff_7/out')
// (3, 16, 'sp4_h_r_14')
// (3, 16, 'sp4_r_v_b_31')
// (3, 17, 'neigh_op_bot_7')
// (3, 17, 'sp4_r_v_b_18')
// (3, 18, 'sp4_r_v_b_7')
// (4, 10, 'sp4_v_t_47')
// (4, 11, 'sp4_v_b_47')
// (4, 12, 'sp4_v_b_34')
// (4, 13, 'sp4_v_b_23')
// (4, 14, 'local_g1_2')
// (4, 14, 'lutff_2/in_1')
// (4, 14, 'sp4_v_b_10')
// (4, 14, 'sp4_v_t_42')
// (4, 15, 'neigh_op_tnl_7')
// (4, 15, 'sp4_v_b_42')
// (4, 16, 'neigh_op_lft_7')
// (4, 16, 'sp4_h_r_27')
// (4, 16, 'sp4_v_b_31')
// (4, 17, 'neigh_op_bnl_7')
// (4, 17, 'sp4_v_b_18')
// (4, 18, 'sp4_v_b_7')
// (5, 13, 'sp4_r_v_b_38')
// (5, 14, 'sp4_r_v_b_27')
// (5, 15, 'local_g2_6')
// (5, 15, 'lutff_7/in_3')
// (5, 15, 'sp4_r_v_b_14')
// (5, 16, 'local_g2_6')
// (5, 16, 'lutff_2/in_0')
// (5, 16, 'sp4_h_r_38')
// (5, 16, 'sp4_r_v_b_3')
// (6, 12, 'sp4_v_t_38')
// (6, 13, 'sp4_v_b_38')
// (6, 14, 'sp4_v_b_27')
// (6, 15, 'sp4_v_b_14')
// (6, 16, 'sp4_h_l_38')
// (6, 16, 'sp4_v_b_3')

reg n450 = 0;
// (2, 15, 'sp4_h_r_4')
// (3, 14, 'neigh_op_tnr_6')
// (3, 15, 'neigh_op_rgt_6')
// (3, 15, 'sp4_h_r_17')
// (3, 16, 'neigh_op_bnr_6')
// (4, 14, 'neigh_op_top_6')
// (4, 15, 'lutff_6/out')
// (4, 15, 'sp4_h_r_28')
// (4, 16, 'neigh_op_bot_6')
// (5, 12, 'local_g3_7')
// (5, 12, 'lutff_0/in_2')
// (5, 12, 'sp4_r_v_b_47')
// (5, 13, 'sp4_r_v_b_34')
// (5, 14, 'neigh_op_tnl_6')
// (5, 14, 'sp4_r_v_b_23')
// (5, 15, 'neigh_op_lft_6')
// (5, 15, 'sp4_h_r_41')
// (5, 15, 'sp4_r_v_b_10')
// (5, 16, 'neigh_op_bnl_6')
// (6, 11, 'sp4_v_t_47')
// (6, 12, 'sp4_v_b_47')
// (6, 13, 'sp4_v_b_34')
// (6, 14, 'sp4_v_b_23')
// (6, 15, 'sp4_h_l_41')
// (6, 15, 'sp4_v_b_10')

wire n451;
// (2, 15, 'sp4_h_r_9')
// (3, 15, 'sp12_h_r_0')
// (3, 15, 'sp4_h_r_20')
// (4, 14, 'neigh_op_tnr_6')
// (4, 15, 'local_g1_3')
// (4, 15, 'lutff_global/cen')
// (4, 15, 'neigh_op_rgt_6')
// (4, 15, 'sp12_h_r_3')
// (4, 15, 'sp4_h_r_33')
// (4, 16, 'neigh_op_bnr_6')
// (5, 12, 'sp4_r_v_b_38')
// (5, 13, 'sp4_r_v_b_27')
// (5, 14, 'neigh_op_top_6')
// (5, 14, 'sp4_r_v_b_14')
// (5, 15, 'local_g1_3')
// (5, 15, 'lutff_6/out')
// (5, 15, 'lutff_global/cen')
// (5, 15, 'sp12_h_r_4')
// (5, 15, 'sp4_h_r_44')
// (5, 15, 'sp4_r_v_b_3')
// (5, 16, 'neigh_op_bot_6')
// (6, 11, 'sp4_v_t_38')
// (6, 12, 'sp4_v_b_38')
// (6, 13, 'sp4_v_b_27')
// (6, 14, 'neigh_op_tnl_6')
// (6, 14, 'sp4_v_b_14')
// (6, 15, 'neigh_op_lft_6')
// (6, 15, 'sp12_h_r_7')
// (6, 15, 'sp4_h_l_44')
// (6, 15, 'sp4_v_b_3')
// (6, 16, 'neigh_op_bnl_6')
// (7, 15, 'sp12_h_r_8')
// (8, 15, 'sp12_h_r_11')
// (9, 15, 'sp12_h_r_12')
// (10, 15, 'sp12_h_r_15')
// (11, 15, 'sp12_h_r_16')
// (12, 15, 'sp12_h_r_19')
// (13, 15, 'sp12_h_r_20')
// (14, 15, 'sp12_h_r_23')
// (15, 15, 'sp12_h_l_23')

reg n452 = 0;
// (2, 16, 'local_g0_4')
// (2, 16, 'local_g1_4')
// (2, 16, 'lutff_0/in_1')
// (2, 16, 'lutff_4/in_1')
// (2, 16, 'lutff_5/in_3')
// (2, 16, 'lutff_7/in_0')
// (2, 16, 'sp4_h_r_4')
// (3, 15, 'local_g2_6')
// (3, 15, 'lutff_6/in_0')
// (3, 15, 'neigh_op_tnr_6')
// (3, 16, 'neigh_op_rgt_6')
// (3, 16, 'sp4_h_r_17')
// (3, 17, 'neigh_op_bnr_6')
// (4, 10, 'sp4_r_v_b_45')
// (4, 11, 'local_g0_3')
// (4, 11, 'lutff_7/in_0')
// (4, 11, 'sp4_r_v_b_32')
// (4, 12, 'sp4_r_v_b_21')
// (4, 13, 'sp4_r_v_b_8')
// (4, 14, 'sp4_r_v_b_37')
// (4, 15, 'neigh_op_top_6')
// (4, 15, 'sp4_r_v_b_24')
// (4, 16, 'local_g0_6')
// (4, 16, 'lutff_6/in_2')
// (4, 16, 'lutff_6/out')
// (4, 16, 'sp4_h_r_28')
// (4, 16, 'sp4_r_v_b_13')
// (4, 17, 'neigh_op_bot_6')
// (4, 17, 'sp4_r_v_b_0')
// (5, 9, 'sp4_v_t_45')
// (5, 10, 'sp4_v_b_45')
// (5, 11, 'sp4_v_b_32')
// (5, 12, 'sp4_v_b_21')
// (5, 13, 'sp4_v_b_8')
// (5, 13, 'sp4_v_t_37')
// (5, 14, 'sp4_v_b_37')
// (5, 15, 'neigh_op_tnl_6')
// (5, 15, 'sp4_v_b_24')
// (5, 16, 'neigh_op_lft_6')
// (5, 16, 'sp4_h_r_41')
// (5, 16, 'sp4_v_b_13')
// (5, 17, 'neigh_op_bnl_6')
// (5, 17, 'sp4_v_b_0')
// (6, 16, 'sp4_h_l_41')

wire n453;
// (2, 16, 'neigh_op_tnr_3')
// (2, 17, 'neigh_op_rgt_3')
// (2, 18, 'neigh_op_bnr_3')
// (3, 14, 'sp4_r_v_b_42')
// (3, 15, 'local_g0_7')
// (3, 15, 'lutff_7/in_2')
// (3, 15, 'sp4_r_v_b_31')
// (3, 16, 'neigh_op_top_3')
// (3, 16, 'sp4_r_v_b_18')
// (3, 17, 'lutff_3/out')
// (3, 17, 'sp4_r_v_b_7')
// (3, 18, 'neigh_op_bot_3')
// (4, 13, 'sp4_v_t_42')
// (4, 14, 'sp4_v_b_42')
// (4, 15, 'sp4_v_b_31')
// (4, 16, 'neigh_op_tnl_3')
// (4, 16, 'sp4_v_b_18')
// (4, 17, 'neigh_op_lft_3')
// (4, 17, 'sp4_v_b_7')
// (4, 18, 'neigh_op_bnl_3')

wire n454;
// (2, 16, 'neigh_op_tnr_6')
// (2, 17, 'neigh_op_rgt_6')
// (2, 18, 'neigh_op_bnr_6')
// (3, 16, 'neigh_op_top_6')
// (3, 17, 'lutff_6/out')
// (3, 18, 'neigh_op_bot_6')
// (4, 16, 'neigh_op_tnl_6')
// (4, 17, 'local_g0_6')
// (4, 17, 'lutff_0/in_0')
// (4, 17, 'neigh_op_lft_6')
// (4, 18, 'neigh_op_bnl_6')

reg n455 = 0;
// (2, 16, 'sp4_h_r_8')
// (3, 13, 'sp4_r_v_b_37')
// (3, 14, 'sp4_r_v_b_24')
// (3, 15, 'neigh_op_tnr_0')
// (3, 15, 'sp4_r_v_b_13')
// (3, 16, 'neigh_op_rgt_0')
// (3, 16, 'sp4_h_r_21')
// (3, 16, 'sp4_r_v_b_0')
// (3, 17, 'neigh_op_bnr_0')
// (4, 10, 'sp4_r_v_b_41')
// (4, 11, 'sp4_r_v_b_28')
// (4, 12, 'sp4_r_v_b_17')
// (4, 12, 'sp4_v_t_37')
// (4, 13, 'sp4_r_v_b_4')
// (4, 13, 'sp4_v_b_37')
// (4, 14, 'local_g3_1')
// (4, 14, 'lutff_3/in_3')
// (4, 14, 'sp4_r_v_b_41')
// (4, 14, 'sp4_v_b_24')
// (4, 15, 'local_g1_5')
// (4, 15, 'lutff_1/in_1')
// (4, 15, 'neigh_op_top_0')
// (4, 15, 'sp4_r_v_b_28')
// (4, 15, 'sp4_v_b_13')
// (4, 16, 'local_g3_0')
// (4, 16, 'lutff_0/in_3')
// (4, 16, 'lutff_0/out')
// (4, 16, 'lutff_4/in_3')
// (4, 16, 'sp4_h_r_32')
// (4, 16, 'sp4_r_v_b_17')
// (4, 16, 'sp4_v_b_0')
// (4, 17, 'neigh_op_bot_0')
// (4, 17, 'sp4_r_v_b_4')
// (5, 9, 'sp4_v_t_41')
// (5, 10, 'sp4_v_b_41')
// (5, 11, 'sp4_v_b_28')
// (5, 12, 'local_g1_1')
// (5, 12, 'lutff_6/in_2')
// (5, 12, 'sp4_v_b_17')
// (5, 13, 'local_g1_4')
// (5, 13, 'lutff_0/in_1')
// (5, 13, 'sp4_h_r_4')
// (5, 13, 'sp4_v_b_4')
// (5, 13, 'sp4_v_t_41')
// (5, 14, 'sp4_v_b_41')
// (5, 15, 'neigh_op_tnl_0')
// (5, 15, 'sp4_v_b_28')
// (5, 16, 'local_g3_5')
// (5, 16, 'lutff_5/in_3')
// (5, 16, 'neigh_op_lft_0')
// (5, 16, 'sp4_h_r_45')
// (5, 16, 'sp4_v_b_17')
// (5, 17, 'neigh_op_bnl_0')
// (5, 17, 'sp4_v_b_4')
// (6, 13, 'sp4_h_r_17')
// (6, 16, 'sp4_h_l_45')
// (7, 13, 'sp4_h_r_28')
// (8, 13, 'sp4_h_r_41')
// (9, 13, 'sp4_h_l_41')

reg n456 = 0;
// (2, 17, 'local_g0_0')
// (2, 17, 'lutff_1/in_1')
// (2, 17, 'sp4_h_r_8')
// (3, 16, 'neigh_op_tnr_0')
// (3, 17, 'local_g2_0')
// (3, 17, 'lutff_6/in_2')
// (3, 17, 'neigh_op_rgt_0')
// (3, 17, 'sp4_h_r_21')
// (3, 18, 'neigh_op_bnr_0')
// (4, 16, 'neigh_op_top_0')
// (4, 17, 'local_g1_0')
// (4, 17, 'lutff_0/out')
// (4, 17, 'lutff_1/in_2')
// (4, 17, 'sp4_h_r_32')
// (4, 18, 'neigh_op_bot_0')
// (5, 16, 'neigh_op_tnl_0')
// (5, 17, 'neigh_op_lft_0')
// (5, 17, 'sp4_h_r_45')
// (5, 18, 'neigh_op_bnl_0')
// (6, 17, 'sp4_h_l_45')

wire n457;
// (2, 17, 'local_g3_4')
// (2, 17, 'lutff_3/in_0')
// (2, 17, 'neigh_op_tnr_4')
// (2, 18, 'neigh_op_rgt_4')
// (2, 19, 'neigh_op_bnr_4')
// (3, 17, 'local_g0_4')
// (3, 17, 'lutff_3/in_1')
// (3, 17, 'neigh_op_top_4')
// (3, 18, 'lutff_4/out')
// (3, 19, 'neigh_op_bot_4')
// (4, 17, 'neigh_op_tnl_4')
// (4, 18, 'neigh_op_lft_4')
// (4, 19, 'neigh_op_bnl_4')

wire n458;
// (2, 17, 'lutff_1/cout')
// (2, 17, 'lutff_2/in_3')

wire n459;
// (2, 17, 'neigh_op_tnr_1')
// (2, 18, 'local_g2_1')
// (2, 18, 'lutff_3/in_0')
// (2, 18, 'neigh_op_rgt_1')
// (2, 19, 'neigh_op_bnr_1')
// (3, 17, 'neigh_op_top_1')
// (3, 18, 'lutff_1/out')
// (3, 19, 'neigh_op_bot_1')
// (4, 17, 'neigh_op_tnl_1')
// (4, 18, 'neigh_op_lft_1')
// (4, 19, 'neigh_op_bnl_1')

wire n460;
// (2, 17, 'neigh_op_tnr_2')
// (2, 18, 'neigh_op_rgt_2')
// (2, 19, 'neigh_op_bnr_2')
// (3, 17, 'neigh_op_top_2')
// (3, 18, 'local_g1_2')
// (3, 18, 'lutff_2/out')
// (3, 18, 'lutff_3/in_0')
// (3, 19, 'neigh_op_bot_2')
// (4, 17, 'neigh_op_tnl_2')
// (4, 18, 'neigh_op_lft_2')
// (4, 19, 'neigh_op_bnl_2')

reg n461 = 0;
// (2, 17, 'neigh_op_tnr_3')
// (2, 18, 'neigh_op_rgt_3')
// (2, 19, 'neigh_op_bnr_3')
// (3, 17, 'neigh_op_top_3')
// (3, 18, 'local_g2_3')
// (3, 18, 'lutff_2/in_1')
// (3, 18, 'lutff_3/out')
// (3, 18, 'lutff_6/in_3')
// (3, 19, 'neigh_op_bot_3')
// (4, 17, 'neigh_op_tnl_3')
// (4, 18, 'neigh_op_lft_3')
// (4, 19, 'neigh_op_bnl_3')

wire n462;
// (2, 17, 'neigh_op_tnr_5')
// (2, 18, 'neigh_op_rgt_5')
// (2, 19, 'neigh_op_bnr_5')
// (3, 17, 'neigh_op_top_5')
// (3, 18, 'lutff_5/out')
// (3, 19, 'local_g0_5')
// (3, 19, 'lutff_6/in_1')
// (3, 19, 'neigh_op_bot_5')
// (4, 17, 'local_g3_5')
// (4, 17, 'lutff_2/in_2')
// (4, 17, 'neigh_op_tnl_5')
// (4, 18, 'neigh_op_lft_5')
// (4, 19, 'neigh_op_bnl_5')

wire n463;
// (2, 17, 'neigh_op_tnr_6')
// (2, 18, 'neigh_op_rgt_6')
// (2, 19, 'neigh_op_bnr_6')
// (3, 17, 'neigh_op_top_6')
// (3, 18, 'local_g0_6')
// (3, 18, 'lutff_5/in_3')
// (3, 18, 'lutff_6/out')
// (3, 19, 'neigh_op_bot_6')
// (4, 17, 'neigh_op_tnl_6')
// (4, 18, 'neigh_op_lft_6')
// (4, 19, 'neigh_op_bnl_6')

wire n464;
// (2, 17, 'neigh_op_tnr_7')
// (2, 18, 'neigh_op_rgt_7')
// (2, 19, 'neigh_op_bnr_7')
// (3, 17, 'neigh_op_top_7')
// (3, 18, 'local_g2_7')
// (3, 18, 'lutff_5/in_0')
// (3, 18, 'lutff_7/out')
// (3, 19, 'neigh_op_bot_7')
// (4, 17, 'neigh_op_tnl_7')
// (4, 18, 'neigh_op_lft_7')
// (4, 19, 'local_g2_7')
// (4, 19, 'lutff_6/in_1')
// (4, 19, 'neigh_op_bnl_7')

reg n465 = 0;
// (2, 17, 'sp4_h_r_7')
// (3, 17, 'local_g0_2')
// (3, 17, 'lutff_0/in_2')
// (3, 17, 'lutff_1/in_3')
// (3, 17, 'lutff_4/in_0')
// (3, 17, 'sp4_h_r_18')
// (4, 17, 'sp4_h_r_31')
// (5, 17, 'sp4_h_r_42')
// (6, 16, 'neigh_op_tnr_1')
// (6, 17, 'neigh_op_rgt_1')
// (6, 17, 'sp4_h_l_42')
// (6, 17, 'sp4_h_r_7')
// (6, 18, 'neigh_op_bnr_1')
// (7, 16, 'neigh_op_top_1')
// (7, 17, 'local_g0_1')
// (7, 17, 'lutff_1/in_2')
// (7, 17, 'lutff_1/out')
// (7, 17, 'sp4_h_r_18')
// (7, 18, 'neigh_op_bot_1')
// (8, 16, 'neigh_op_tnl_1')
// (8, 17, 'neigh_op_lft_1')
// (8, 17, 'sp4_h_r_31')
// (8, 18, 'neigh_op_bnl_1')
// (9, 17, 'sp4_h_r_42')
// (10, 17, 'sp4_h_l_42')

wire n466;
// (2, 17, 'sp4_r_v_b_45')
// (2, 18, 'sp4_r_v_b_32')
// (2, 19, 'neigh_op_tnr_4')
// (2, 19, 'sp4_r_v_b_21')
// (2, 20, 'neigh_op_rgt_4')
// (2, 20, 'sp4_r_v_b_8')
// (2, 21, 'neigh_op_bnr_4')
// (3, 16, 'sp4_v_t_45')
// (3, 17, 'local_g3_5')
// (3, 17, 'lutff_7/in_3')
// (3, 17, 'sp4_v_b_45')
// (3, 18, 'sp4_v_b_32')
// (3, 19, 'neigh_op_top_4')
// (3, 19, 'sp4_v_b_21')
// (3, 20, 'lutff_4/out')
// (3, 20, 'sp4_h_r_8')
// (3, 20, 'sp4_r_v_b_41')
// (3, 20, 'sp4_v_b_8')
// (3, 21, 'neigh_op_bot_4')
// (3, 21, 'sp4_r_v_b_28')
// (3, 22, 'sp4_r_v_b_17')
// (3, 23, 'sp4_r_v_b_4')
// (4, 19, 'neigh_op_tnl_4')
// (4, 19, 'sp4_h_r_4')
// (4, 19, 'sp4_v_t_41')
// (4, 20, 'neigh_op_lft_4')
// (4, 20, 'sp4_h_r_21')
// (4, 20, 'sp4_v_b_41')
// (4, 21, 'neigh_op_bnl_4')
// (4, 21, 'sp4_v_b_28')
// (4, 22, 'sp4_v_b_17')
// (4, 23, 'sp4_v_b_4')
// (5, 19, 'local_g1_1')
// (5, 19, 'lutff_4/in_2')
// (5, 19, 'sp4_h_r_17')
// (5, 20, 'sp4_h_r_32')
// (6, 19, 'sp4_h_r_28')
// (6, 20, 'sp4_h_r_45')
// (7, 19, 'sp4_h_r_41')
// (7, 20, 'sp4_h_l_45')
// (7, 20, 'sp4_h_r_4')
// (8, 19, 'sp4_h_l_41')
// (8, 20, 'local_g0_1')
// (8, 20, 'lutff_7/in_0')
// (8, 20, 'sp4_h_r_17')
// (9, 20, 'sp4_h_r_28')
// (10, 20, 'sp4_h_r_41')
// (10, 21, 'sp4_r_v_b_44')
// (10, 22, 'sp4_r_v_b_33')
// (10, 23, 'sp4_r_v_b_20')
// (10, 24, 'sp4_r_v_b_9')
// (10, 25, 'sp4_r_v_b_40')
// (10, 26, 'sp4_r_v_b_29')
// (10, 27, 'sp4_r_v_b_16')
// (10, 28, 'sp4_r_v_b_5')
// (10, 29, 'sp4_r_v_b_40')
// (10, 30, 'sp4_r_v_b_29')
// (11, 20, 'sp4_h_l_41')
// (11, 20, 'sp4_v_t_44')
// (11, 21, 'sp4_v_b_44')
// (11, 22, 'sp4_v_b_33')
// (11, 23, 'sp4_v_b_20')
// (11, 24, 'sp4_v_b_9')
// (11, 24, 'sp4_v_t_40')
// (11, 25, 'sp4_v_b_40')
// (11, 26, 'sp4_v_b_29')
// (11, 27, 'sp4_v_b_16')
// (11, 28, 'sp4_v_b_5')
// (11, 28, 'sp4_v_t_40')
// (11, 29, 'sp4_v_b_40')
// (11, 30, 'local_g3_5')
// (11, 30, 'lutff_0/in_2')
// (11, 30, 'sp4_v_b_29')
// (11, 31, 'span4_vert_16')

wire n467;
// (2, 18, 'neigh_op_tnr_1')
// (2, 19, 'neigh_op_rgt_1')
// (2, 20, 'neigh_op_bnr_1')
// (3, 18, 'neigh_op_top_1')
// (3, 19, 'lutff_1/out')
// (3, 20, 'neigh_op_bot_1')
// (4, 18, 'neigh_op_tnl_1')
// (4, 19, 'neigh_op_lft_1')
// (4, 20, 'local_g3_1')
// (4, 20, 'lutff_7/in_3')
// (4, 20, 'neigh_op_bnl_1')

wire n468;
// (2, 18, 'neigh_op_tnr_2')
// (2, 19, 'neigh_op_rgt_2')
// (2, 20, 'neigh_op_bnr_2')
// (3, 18, 'neigh_op_top_2')
// (3, 19, 'lutff_2/out')
// (3, 20, 'local_g0_2')
// (3, 20, 'lutff_2/in_2')
// (3, 20, 'neigh_op_bot_2')
// (4, 18, 'neigh_op_tnl_2')
// (4, 19, 'neigh_op_lft_2')
// (4, 20, 'neigh_op_bnl_2')

wire n469;
// (2, 18, 'neigh_op_tnr_3')
// (2, 19, 'neigh_op_rgt_3')
// (2, 20, 'neigh_op_bnr_3')
// (3, 18, 'neigh_op_top_3')
// (3, 19, 'lutff_3/out')
// (3, 19, 'sp4_r_v_b_39')
// (3, 20, 'local_g1_2')
// (3, 20, 'lutff_3/in_0')
// (3, 20, 'neigh_op_bot_3')
// (3, 20, 'sp4_r_v_b_26')
// (3, 21, 'sp4_r_v_b_15')
// (3, 22, 'sp4_r_v_b_2')
// (4, 18, 'neigh_op_tnl_3')
// (4, 18, 'sp4_v_t_39')
// (4, 19, 'neigh_op_lft_3')
// (4, 19, 'sp4_v_b_39')
// (4, 20, 'neigh_op_bnl_3')
// (4, 20, 'sp4_v_b_26')
// (4, 21, 'sp4_v_b_15')
// (4, 22, 'sp4_v_b_2')

wire n470;
// (2, 18, 'neigh_op_tnr_4')
// (2, 19, 'neigh_op_rgt_4')
// (2, 20, 'neigh_op_bnr_4')
// (3, 18, 'neigh_op_top_4')
// (3, 19, 'lutff_4/out')
// (3, 20, 'neigh_op_bot_4')
// (4, 18, 'neigh_op_tnl_4')
// (4, 19, 'neigh_op_lft_4')
// (4, 20, 'local_g2_4')
// (4, 20, 'lutff_4/in_2')
// (4, 20, 'neigh_op_bnl_4')

wire n471;
// (2, 18, 'neigh_op_tnr_5')
// (2, 19, 'neigh_op_rgt_5')
// (2, 20, 'neigh_op_bnr_5')
// (3, 18, 'neigh_op_top_5')
// (3, 19, 'lutff_5/out')
// (3, 20, 'local_g0_5')
// (3, 20, 'lutff_6/in_1')
// (3, 20, 'neigh_op_bot_5')
// (4, 18, 'neigh_op_tnl_5')
// (4, 19, 'neigh_op_lft_5')
// (4, 20, 'neigh_op_bnl_5')

wire n472;
// (2, 18, 'neigh_op_tnr_6')
// (2, 19, 'neigh_op_rgt_6')
// (2, 20, 'neigh_op_bnr_6')
// (3, 18, 'neigh_op_top_6')
// (3, 19, 'lutff_6/out')
// (3, 20, 'neigh_op_bot_6')
// (4, 18, 'neigh_op_tnl_6')
// (4, 19, 'local_g1_6')
// (4, 19, 'lutff_7/in_2')
// (4, 19, 'neigh_op_lft_6')
// (4, 20, 'neigh_op_bnl_6')

wire n473;
// (2, 18, 'neigh_op_tnr_7')
// (2, 19, 'neigh_op_rgt_7')
// (2, 20, 'neigh_op_bnr_7')
// (3, 18, 'local_g0_7')
// (3, 18, 'lutff_7/in_0')
// (3, 18, 'neigh_op_top_7')
// (3, 19, 'lutff_7/out')
// (3, 20, 'local_g1_7')
// (3, 20, 'lutff_1/in_1')
// (3, 20, 'neigh_op_bot_7')
// (4, 18, 'neigh_op_tnl_7')
// (4, 19, 'neigh_op_lft_7')
// (4, 20, 'neigh_op_bnl_7')

wire n474;
// (2, 18, 'sp4_h_r_6')
// (3, 18, 'sp4_h_r_19')
// (3, 19, 'sp4_h_r_2')
// (4, 18, 'neigh_op_tnr_5')
// (4, 18, 'sp4_h_r_30')
// (4, 19, 'neigh_op_rgt_5')
// (4, 19, 'sp4_h_r_15')
// (4, 20, 'neigh_op_bnr_5')
// (5, 18, 'local_g3_3')
// (5, 18, 'lutff_global/cen')
// (5, 18, 'neigh_op_top_5')
// (5, 18, 'sp4_h_r_43')
// (5, 19, 'local_g2_2')
// (5, 19, 'lutff_5/out')
// (5, 19, 'lutff_global/cen')
// (5, 19, 'sp4_h_r_26')
// (5, 19, 'sp4_r_v_b_43')
// (5, 20, 'neigh_op_bot_5')
// (5, 20, 'sp4_r_v_b_30')
// (5, 21, 'sp4_r_v_b_19')
// (5, 22, 'sp4_r_v_b_6')
// (6, 18, 'neigh_op_tnl_5')
// (6, 18, 'sp4_h_l_43')
// (6, 18, 'sp4_v_t_43')
// (6, 19, 'neigh_op_lft_5')
// (6, 19, 'sp4_h_r_39')
// (6, 19, 'sp4_v_b_43')
// (6, 20, 'neigh_op_bnl_5')
// (6, 20, 'sp4_v_b_30')
// (6, 21, 'sp4_v_b_19')
// (6, 22, 'sp4_v_b_6')
// (7, 19, 'sp4_h_l_39')

wire n475;
// (2, 18, 'sp4_r_v_b_42')
// (2, 19, 'local_g3_1')
// (2, 19, 'lutff_4/in_2')
// (2, 19, 'neigh_op_tnr_1')
// (2, 19, 'sp4_r_v_b_31')
// (2, 20, 'local_g3_1')
// (2, 20, 'lutff_0/in_2')
// (2, 20, 'lutff_2/in_2')
// (2, 20, 'neigh_op_rgt_1')
// (2, 20, 'sp4_r_v_b_18')
// (2, 21, 'neigh_op_bnr_1')
// (2, 21, 'sp4_r_v_b_7')
// (3, 17, 'sp4_h_r_0')
// (3, 17, 'sp4_v_t_42')
// (3, 18, 'sp4_v_b_42')
// (3, 19, 'neigh_op_top_1')
// (3, 19, 'sp4_v_b_31')
// (3, 20, 'lutff_1/out')
// (3, 20, 'sp4_v_b_18')
// (3, 21, 'neigh_op_bot_1')
// (3, 21, 'sp4_v_b_7')
// (4, 17, 'sp4_h_r_13')
// (4, 19, 'neigh_op_tnl_1')
// (4, 20, 'neigh_op_lft_1')
// (4, 21, 'neigh_op_bnl_1')
// (5, 17, 'local_g2_0')
// (5, 17, 'lutff_7/in_3')
// (5, 17, 'sp4_h_r_24')
// (6, 17, 'sp4_h_r_37')
// (7, 17, 'sp4_h_l_37')

wire n476;
// (2, 19, 'lutff_1/cout')
// (2, 19, 'lutff_2/in_3')

reg n477 = 0;
// (2, 19, 'neigh_op_tnr_0')
// (2, 20, 'neigh_op_rgt_0')
// (2, 20, 'sp4_h_r_5')
// (2, 21, 'neigh_op_bnr_0')
// (3, 18, 'sp4_r_v_b_41')
// (3, 19, 'local_g1_0')
// (3, 19, 'lutff_2/in_1')
// (3, 19, 'neigh_op_top_0')
// (3, 19, 'sp4_r_v_b_28')
// (3, 19, 'sp4_r_v_b_44')
// (3, 20, 'lutff_0/out')
// (3, 20, 'sp4_h_r_16')
// (3, 20, 'sp4_r_v_b_17')
// (3, 20, 'sp4_r_v_b_33')
// (3, 21, 'neigh_op_bot_0')
// (3, 21, 'sp4_r_v_b_20')
// (3, 21, 'sp4_r_v_b_4')
// (3, 22, 'sp4_r_v_b_9')
// (4, 17, 'sp4_h_r_9')
// (4, 17, 'sp4_v_t_41')
// (4, 18, 'sp4_h_r_2')
// (4, 18, 'sp4_v_b_41')
// (4, 18, 'sp4_v_t_44')
// (4, 19, 'local_g3_0')
// (4, 19, 'lutff_0/in_1')
// (4, 19, 'neigh_op_tnl_0')
// (4, 19, 'sp4_v_b_28')
// (4, 19, 'sp4_v_b_44')
// (4, 20, 'neigh_op_lft_0')
// (4, 20, 'sp4_h_r_29')
// (4, 20, 'sp4_v_b_17')
// (4, 20, 'sp4_v_b_33')
// (4, 21, 'local_g2_0')
// (4, 21, 'lutff_6/in_2')
// (4, 21, 'neigh_op_bnl_0')
// (4, 21, 'sp4_v_b_20')
// (4, 21, 'sp4_v_b_4')
// (4, 22, 'sp4_v_b_9')
// (5, 9, 'sp4_r_v_b_46')
// (5, 10, 'sp4_r_v_b_35')
// (5, 11, 'sp4_r_v_b_22')
// (5, 12, 'sp4_r_v_b_11')
// (5, 13, 'sp4_r_v_b_46')
// (5, 14, 'sp4_r_v_b_35')
// (5, 15, 'sp4_r_v_b_22')
// (5, 16, 'sp4_r_v_b_11')
// (5, 17, 'sp4_h_r_20')
// (5, 17, 'sp4_r_v_b_46')
// (5, 18, 'sp4_h_r_15')
// (5, 18, 'sp4_r_v_b_35')
// (5, 19, 'sp4_r_v_b_22')
// (5, 20, 'sp4_h_r_40')
// (5, 20, 'sp4_r_v_b_11')
// (6, 8, 'sp4_h_r_4')
// (6, 8, 'sp4_v_t_46')
// (6, 9, 'sp4_v_b_46')
// (6, 10, 'sp4_v_b_35')
// (6, 11, 'sp4_v_b_22')
// (6, 12, 'sp4_v_b_11')
// (6, 12, 'sp4_v_t_46')
// (6, 13, 'sp4_v_b_46')
// (6, 14, 'sp4_v_b_35')
// (6, 15, 'sp4_v_b_22')
// (6, 16, 'sp4_h_r_11')
// (6, 16, 'sp4_v_b_11')
// (6, 16, 'sp4_v_t_46')
// (6, 17, 'sp4_h_r_33')
// (6, 17, 'sp4_v_b_46')
// (6, 18, 'sp4_h_r_26')
// (6, 18, 'sp4_v_b_35')
// (6, 19, 'sp4_v_b_22')
// (6, 20, 'sp4_h_l_40')
// (6, 20, 'sp4_v_b_11')
// (7, 8, 'sp4_h_r_17')
// (7, 16, 'sp4_h_r_22')
// (7, 17, 'local_g2_4')
// (7, 17, 'lutff_6/in_0')
// (7, 17, 'sp4_h_r_44')
// (7, 18, 'sp4_h_r_39')
// (8, 8, 'sp4_h_r_28')
// (8, 16, 'sp4_h_r_35')
// (8, 17, 'sp4_h_l_44')
// (8, 18, 'local_g1_5')
// (8, 18, 'lutff_3/in_3')
// (8, 18, 'lutff_5/in_3')
// (8, 18, 'sp4_h_l_39')
// (8, 18, 'sp4_h_r_5')
// (9, 5, 'sp4_r_v_b_41')
// (9, 6, 'sp4_r_v_b_28')
// (9, 7, 'local_g3_1')
// (9, 7, 'lutff_7/in_3')
// (9, 7, 'sp4_r_v_b_17')
// (9, 8, 'sp4_h_r_41')
// (9, 8, 'sp4_r_v_b_4')
// (9, 13, 'sp4_r_v_b_46')
// (9, 14, 'sp4_r_v_b_35')
// (9, 15, 'local_g3_6')
// (9, 15, 'lutff_4/in_3')
// (9, 15, 'sp4_r_v_b_22')
// (9, 16, 'sp4_h_r_46')
// (9, 16, 'sp4_r_v_b_11')
// (9, 18, 'sp4_h_r_16')
// (10, 4, 'sp4_v_t_41')
// (10, 5, 'sp4_v_b_41')
// (10, 6, 'sp4_v_b_28')
// (10, 7, 'sp4_v_b_17')
// (10, 8, 'sp4_h_l_41')
// (10, 8, 'sp4_v_b_4')
// (10, 12, 'sp4_v_t_46')
// (10, 13, 'sp4_v_b_46')
// (10, 14, 'sp4_v_b_35')
// (10, 15, 'sp4_v_b_22')
// (10, 16, 'sp4_h_l_46')
// (10, 16, 'sp4_v_b_11')
// (10, 18, 'sp4_h_r_29')
// (11, 18, 'sp4_h_r_40')
// (12, 18, 'sp4_h_l_40')

wire n478;
// (2, 19, 'neigh_op_tnr_2')
// (2, 20, 'neigh_op_rgt_2')
// (2, 21, 'neigh_op_bnr_2')
// (3, 19, 'neigh_op_top_2')
// (3, 20, 'local_g2_2')
// (3, 20, 'lutff_0/in_2')
// (3, 20, 'lutff_2/out')
// (3, 21, 'neigh_op_bot_2')
// (4, 19, 'neigh_op_tnl_2')
// (4, 20, 'neigh_op_lft_2')
// (4, 21, 'neigh_op_bnl_2')

wire n479;
// (2, 19, 'neigh_op_tnr_3')
// (2, 20, 'neigh_op_rgt_3')
// (2, 21, 'neigh_op_bnr_3')
// (3, 19, 'neigh_op_top_3')
// (3, 20, 'local_g0_3')
// (3, 20, 'lutff_3/out')
// (3, 20, 'lutff_5/in_2')
// (3, 21, 'neigh_op_bot_3')
// (4, 19, 'neigh_op_tnl_3')
// (4, 20, 'neigh_op_lft_3')
// (4, 21, 'neigh_op_bnl_3')

wire n480;
// (2, 19, 'neigh_op_tnr_6')
// (2, 20, 'neigh_op_rgt_6')
// (2, 21, 'neigh_op_bnr_6')
// (3, 19, 'neigh_op_top_6')
// (3, 20, 'lutff_6/out')
// (3, 21, 'neigh_op_bot_6')
// (4, 19, 'neigh_op_tnl_6')
// (4, 20, 'local_g0_6')
// (4, 20, 'lutff_0/in_0')
// (4, 20, 'neigh_op_lft_6')
// (4, 21, 'neigh_op_bnl_6')

wire n481;
// (2, 19, 'sp4_r_v_b_37')
// (2, 20, 'sp4_r_v_b_24')
// (2, 21, 'sp4_r_v_b_13')
// (2, 22, 'sp4_r_v_b_0')
// (3, 18, 'sp4_v_t_37')
// (3, 19, 'sp4_v_b_37')
// (3, 20, 'local_g2_0')
// (3, 20, 'lutff_6/in_0')
// (3, 20, 'sp4_v_b_24')
// (3, 21, 'neigh_op_tnr_1')
// (3, 21, 'sp4_v_b_13')
// (3, 22, 'neigh_op_rgt_1')
// (3, 22, 'sp4_h_r_7')
// (3, 22, 'sp4_v_b_0')
// (3, 23, 'neigh_op_bnr_1')
// (4, 21, 'neigh_op_top_1')
// (4, 22, 'lutff_1/out')
// (4, 22, 'sp4_h_r_18')
// (4, 23, 'neigh_op_bot_1')
// (5, 21, 'neigh_op_tnl_1')
// (5, 22, 'neigh_op_lft_1')
// (5, 22, 'sp4_h_r_31')
// (5, 23, 'neigh_op_bnl_1')
// (6, 22, 'sp4_h_r_42')
// (7, 22, 'sp4_h_l_42')

reg n482 = 0;
// (2, 20, 'neigh_op_tnr_0')
// (2, 21, 'neigh_op_rgt_0')
// (2, 22, 'neigh_op_bnr_0')
// (3, 20, 'neigh_op_top_0')
// (3, 21, 'local_g2_0')
// (3, 21, 'lutff_0/in_2')
// (3, 21, 'lutff_0/out')
// (3, 21, 'lutff_1/in_1')
// (3, 22, 'neigh_op_bot_0')
// (4, 20, 'neigh_op_tnl_0')
// (4, 21, 'neigh_op_lft_0')
// (4, 22, 'neigh_op_bnl_0')

reg n483 = 0;
// (2, 20, 'neigh_op_tnr_3')
// (2, 21, 'neigh_op_rgt_3')
// (2, 21, 'sp4_h_r_11')
// (2, 22, 'neigh_op_bnr_3')
// (3, 13, 'sp4_r_v_b_45')
// (3, 14, 'sp4_r_v_b_32')
// (3, 15, 'sp4_r_v_b_21')
// (3, 16, 'sp4_r_v_b_8')
// (3, 17, 'sp4_r_v_b_40')
// (3, 18, 'sp4_r_v_b_29')
// (3, 19, 'sp4_r_v_b_16')
// (3, 20, 'neigh_op_top_3')
// (3, 20, 'sp4_r_v_b_5')
// (3, 21, 'local_g0_3')
// (3, 21, 'lutff_2/in_1')
// (3, 21, 'lutff_3/out')
// (3, 21, 'lutff_4/in_3')
// (3, 21, 'sp4_h_r_22')
// (3, 21, 'sp4_r_v_b_39')
// (3, 22, 'neigh_op_bot_3')
// (3, 22, 'sp4_r_v_b_26')
// (3, 23, 'sp4_r_v_b_15')
// (3, 24, 'sp4_r_v_b_2')
// (4, 12, 'sp4_h_r_1')
// (4, 12, 'sp4_v_t_45')
// (4, 13, 'sp4_v_b_45')
// (4, 14, 'sp4_v_b_32')
// (4, 15, 'sp4_v_b_21')
// (4, 16, 'sp4_v_b_8')
// (4, 16, 'sp4_v_t_40')
// (4, 17, 'sp4_v_b_40')
// (4, 18, 'sp4_v_b_29')
// (4, 19, 'sp4_v_b_16')
// (4, 20, 'neigh_op_tnl_3')
// (4, 20, 'sp4_v_b_5')
// (4, 20, 'sp4_v_t_39')
// (4, 21, 'neigh_op_lft_3')
// (4, 21, 'sp4_h_r_35')
// (4, 21, 'sp4_v_b_39')
// (4, 22, 'neigh_op_bnl_3')
// (4, 22, 'sp4_v_b_26')
// (4, 23, 'sp4_v_b_15')
// (4, 24, 'sp4_v_b_2')
// (5, 12, 'local_g0_4')
// (5, 12, 'lutff_2/in_0')
// (5, 12, 'sp4_h_r_12')
// (5, 21, 'sp4_h_r_46')
// (6, 12, 'sp4_h_r_25')
// (6, 21, 'sp4_h_l_46')
// (6, 21, 'sp4_h_r_11')
// (7, 12, 'sp4_h_r_36')
// (7, 21, 'sp4_h_r_22')
// (8, 12, 'sp4_h_l_36')
// (8, 21, 'sp4_h_r_35')
// (9, 10, 'sp4_r_v_b_46')
// (9, 11, 'sp4_r_v_b_35')
// (9, 12, 'sp4_r_v_b_22')
// (9, 13, 'sp4_r_v_b_11')
// (9, 14, 'sp4_r_v_b_45')
// (9, 15, 'sp4_r_v_b_32')
// (9, 16, 'sp4_r_v_b_21')
// (9, 17, 'sp4_r_v_b_8')
// (9, 18, 'sp4_r_v_b_40')
// (9, 19, 'sp4_r_v_b_29')
// (9, 20, 'sp4_r_v_b_16')
// (9, 21, 'sp4_h_r_46')
// (9, 21, 'sp4_r_v_b_5')
// (10, 9, 'sp4_v_t_46')
// (10, 10, 'sp4_v_b_46')
// (10, 11, 'local_g3_3')
// (10, 11, 'lutff_5/in_3')
// (10, 11, 'sp4_v_b_35')
// (10, 12, 'sp4_v_b_22')
// (10, 13, 'sp4_v_b_11')
// (10, 13, 'sp4_v_t_45')
// (10, 14, 'sp4_v_b_45')
// (10, 15, 'sp4_v_b_32')
// (10, 16, 'sp4_v_b_21')
// (10, 17, 'sp4_v_b_8')
// (10, 17, 'sp4_v_t_40')
// (10, 18, 'sp4_v_b_40')
// (10, 19, 'sp4_v_b_29')
// (10, 20, 'sp4_v_b_16')
// (10, 21, 'sp4_h_l_46')
// (10, 21, 'sp4_v_b_5')

wire n484;
// (2, 20, 'neigh_op_tnr_4')
// (2, 21, 'neigh_op_rgt_4')
// (2, 22, 'neigh_op_bnr_4')
// (3, 20, 'neigh_op_top_4')
// (3, 21, 'local_g2_4')
// (3, 21, 'lutff_3/in_1')
// (3, 21, 'lutff_4/out')
// (3, 22, 'neigh_op_bot_4')
// (4, 20, 'neigh_op_tnl_4')
// (4, 21, 'neigh_op_lft_4')
// (4, 22, 'neigh_op_bnl_4')

reg n485 = 0;
// (2, 20, 'neigh_op_tnr_5')
// (2, 21, 'neigh_op_rgt_5')
// (2, 22, 'neigh_op_bnr_5')
// (3, 20, 'neigh_op_top_5')
// (3, 21, 'local_g0_5')
// (3, 21, 'lutff_5/out')
// (3, 21, 'lutff_7/in_2')
// (3, 21, 'sp4_h_r_10')
// (3, 22, 'neigh_op_bot_5')
// (4, 20, 'neigh_op_tnl_5')
// (4, 21, 'neigh_op_lft_5')
// (4, 21, 'sp4_h_r_23')
// (4, 22, 'neigh_op_bnl_5')
// (5, 21, 'sp4_h_r_34')
// (6, 21, 'sp4_h_r_47')
// (7, 21, 'local_g0_1')
// (7, 21, 'lutff_5/in_2')
// (7, 21, 'sp4_h_l_47')
// (7, 21, 'sp4_h_r_1')
// (8, 21, 'sp4_h_r_12')
// (9, 21, 'sp4_h_r_25')
// (10, 21, 'sp4_h_r_36')
// (11, 21, 'sp4_h_l_36')

reg n486 = 0;
// (2, 20, 'neigh_op_tnr_6')
// (2, 21, 'neigh_op_rgt_6')
// (2, 22, 'neigh_op_bnr_6')
// (3, 20, 'local_g0_6')
// (3, 20, 'lutff_4/in_0')
// (3, 20, 'neigh_op_top_6')
// (3, 21, 'local_g3_6')
// (3, 21, 'lutff_4/in_1')
// (3, 21, 'lutff_6/out')
// (3, 21, 'lutff_7/in_0')
// (3, 22, 'neigh_op_bot_6')
// (4, 20, 'neigh_op_tnl_6')
// (4, 21, 'neigh_op_lft_6')
// (4, 22, 'neigh_op_bnl_6')

wire n487;
// (2, 20, 'neigh_op_tnr_7')
// (2, 21, 'neigh_op_rgt_7')
// (2, 22, 'neigh_op_bnr_7')
// (3, 20, 'neigh_op_top_7')
// (3, 21, 'local_g2_7')
// (3, 21, 'lutff_0/in_1')
// (3, 21, 'lutff_7/out')
// (3, 22, 'neigh_op_bot_7')
// (4, 20, 'neigh_op_tnl_7')
// (4, 21, 'neigh_op_lft_7')
// (4, 22, 'neigh_op_bnl_7')

reg n488 = 0;
// (2, 20, 'sp4_h_r_10')
// (3, 19, 'local_g2_1')
// (3, 19, 'lutff_4/in_1')
// (3, 19, 'neigh_op_tnr_1')
// (3, 20, 'neigh_op_rgt_1')
// (3, 20, 'sp4_h_r_23')
// (3, 20, 'sp4_h_r_7')
// (3, 21, 'neigh_op_bnr_1')
// (4, 17, 'sp4_r_v_b_38')
// (4, 18, 'sp4_r_v_b_27')
// (4, 19, 'local_g0_1')
// (4, 19, 'lutff_3/in_2')
// (4, 19, 'neigh_op_top_1')
// (4, 19, 'sp4_r_v_b_14')
// (4, 19, 'sp4_r_v_b_46')
// (4, 20, 'local_g2_1')
// (4, 20, 'lutff_1/out')
// (4, 20, 'lutff_2/in_1')
// (4, 20, 'sp4_h_r_18')
// (4, 20, 'sp4_h_r_34')
// (4, 20, 'sp4_r_v_b_3')
// (4, 20, 'sp4_r_v_b_35')
// (4, 21, 'neigh_op_bot_1')
// (4, 21, 'sp4_r_v_b_22')
// (4, 22, 'local_g2_3')
// (4, 22, 'lutff_0/in_1')
// (4, 22, 'sp4_r_v_b_11')
// (5, 16, 'sp4_h_r_3')
// (5, 16, 'sp4_v_t_38')
// (5, 17, 'sp4_v_b_38')
// (5, 18, 'sp4_v_b_27')
// (5, 18, 'sp4_v_t_46')
// (5, 19, 'neigh_op_tnl_1')
// (5, 19, 'sp4_v_b_14')
// (5, 19, 'sp4_v_b_46')
// (5, 20, 'neigh_op_lft_1')
// (5, 20, 'sp4_h_r_31')
// (5, 20, 'sp4_h_r_47')
// (5, 20, 'sp4_v_b_3')
// (5, 20, 'sp4_v_b_35')
// (5, 21, 'neigh_op_bnl_1')
// (5, 21, 'sp4_v_b_22')
// (5, 22, 'sp4_v_b_11')
// (6, 16, 'sp4_h_r_14')
// (6, 17, 'sp4_r_v_b_36')
// (6, 18, 'sp4_r_v_b_25')
// (6, 19, 'sp4_r_v_b_12')
// (6, 20, 'sp4_h_l_47')
// (6, 20, 'sp4_h_r_1')
// (6, 20, 'sp4_h_r_42')
// (6, 20, 'sp4_r_v_b_1')
// (7, 16, 'local_g3_3')
// (7, 16, 'lutff_7/in_3')
// (7, 16, 'sp4_h_r_27')
// (7, 16, 'sp4_v_t_36')
// (7, 17, 'sp4_v_b_36')
// (7, 18, 'sp4_v_b_25')
// (7, 19, 'local_g0_4')
// (7, 19, 'lutff_7/in_1')
// (7, 19, 'sp4_v_b_12')
// (7, 20, 'sp4_h_l_42')
// (7, 20, 'sp4_h_r_12')
// (7, 20, 'sp4_v_b_1')
// (8, 9, 'sp4_r_v_b_46')
// (8, 10, 'sp4_r_v_b_35')
// (8, 11, 'sp4_r_v_b_22')
// (8, 12, 'sp4_r_v_b_11')
// (8, 13, 'sp4_r_v_b_38')
// (8, 14, 'sp4_r_v_b_27')
// (8, 15, 'sp4_r_v_b_14')
// (8, 16, 'sp4_h_r_38')
// (8, 16, 'sp4_r_v_b_3')
// (8, 20, 'sp4_h_r_25')
// (9, 8, 'sp4_v_t_46')
// (9, 9, 'local_g3_6')
// (9, 9, 'lutff_7/in_2')
// (9, 9, 'sp4_v_b_46')
// (9, 10, 'sp4_v_b_35')
// (9, 11, 'sp4_v_b_22')
// (9, 12, 'sp4_v_b_11')
// (9, 12, 'sp4_v_t_38')
// (9, 13, 'sp4_v_b_38')
// (9, 14, 'sp4_v_b_27')
// (9, 15, 'local_g0_6')
// (9, 15, 'lutff_4/in_0')
// (9, 15, 'sp4_v_b_14')
// (9, 16, 'sp4_h_l_38')
// (9, 16, 'sp4_v_b_3')
// (9, 17, 'sp4_r_v_b_36')
// (9, 18, 'sp4_r_v_b_25')
// (9, 19, 'local_g2_4')
// (9, 19, 'lutff_6/in_2')
// (9, 19, 'sp4_r_v_b_12')
// (9, 20, 'sp4_h_r_36')
// (9, 20, 'sp4_r_v_b_1')
// (10, 16, 'sp4_v_t_36')
// (10, 17, 'sp4_v_b_36')
// (10, 18, 'sp4_v_b_25')
// (10, 19, 'sp4_v_b_12')
// (10, 20, 'sp4_h_l_36')
// (10, 20, 'sp4_v_b_1')

wire n489;
// (2, 20, 'sp4_h_r_4')
// (3, 19, 'neigh_op_tnr_6')
// (3, 20, 'local_g0_1')
// (3, 20, 'lutff_0/in_1')
// (3, 20, 'neigh_op_rgt_6')
// (3, 20, 'sp4_h_r_17')
// (3, 21, 'neigh_op_bnr_6')
// (4, 19, 'neigh_op_top_6')
// (4, 20, 'lutff_6/out')
// (4, 20, 'sp4_h_r_28')
// (4, 21, 'neigh_op_bot_6')
// (5, 19, 'neigh_op_tnl_6')
// (5, 20, 'neigh_op_lft_6')
// (5, 20, 'sp4_h_r_41')
// (5, 21, 'neigh_op_bnl_6')
// (6, 20, 'sp4_h_l_41')

reg n490 = 0;
// (2, 20, 'sp4_h_r_8')
// (3, 19, 'local_g3_0')
// (3, 19, 'lutff_5/in_2')
// (3, 19, 'neigh_op_tnr_0')
// (3, 20, 'neigh_op_rgt_0')
// (3, 20, 'sp4_h_r_21')
// (3, 21, 'neigh_op_bnr_0')
// (4, 18, 'sp4_r_v_b_41')
// (4, 19, 'local_g1_0')
// (4, 19, 'lutff_4/in_1')
// (4, 19, 'neigh_op_top_0')
// (4, 19, 'sp4_r_v_b_28')
// (4, 19, 'sp4_r_v_b_44')
// (4, 20, 'lutff_0/out')
// (4, 20, 'sp4_h_r_0')
// (4, 20, 'sp4_h_r_32')
// (4, 20, 'sp4_r_v_b_17')
// (4, 20, 'sp4_r_v_b_33')
// (4, 21, 'neigh_op_bot_0')
// (4, 21, 'sp4_r_v_b_20')
// (4, 21, 'sp4_r_v_b_4')
// (4, 22, 'local_g2_1')
// (4, 22, 'lutff_1/in_0')
// (4, 22, 'sp4_r_v_b_9')
// (5, 17, 'sp4_h_r_9')
// (5, 17, 'sp4_v_t_41')
// (5, 18, 'sp4_v_b_41')
// (5, 18, 'sp4_v_t_44')
// (5, 19, 'neigh_op_tnl_0')
// (5, 19, 'sp4_v_b_28')
// (5, 19, 'sp4_v_b_44')
// (5, 20, 'neigh_op_lft_0')
// (5, 20, 'sp4_h_r_13')
// (5, 20, 'sp4_h_r_45')
// (5, 20, 'sp4_v_b_17')
// (5, 20, 'sp4_v_b_33')
// (5, 21, 'neigh_op_bnl_0')
// (5, 21, 'sp4_v_b_20')
// (5, 21, 'sp4_v_b_4')
// (5, 22, 'sp4_v_b_9')
// (6, 17, 'sp4_h_r_20')
// (6, 20, 'sp4_h_l_45')
// (6, 20, 'sp4_h_r_24')
// (6, 20, 'sp4_h_r_4')
// (7, 17, 'sp4_h_r_33')
// (7, 17, 'sp4_r_v_b_37')
// (7, 18, 'sp4_r_v_b_24')
// (7, 19, 'local_g2_5')
// (7, 19, 'lutff_4/in_3')
// (7, 19, 'lutff_7/in_2')
// (7, 19, 'sp4_r_v_b_13')
// (7, 20, 'sp4_h_r_17')
// (7, 20, 'sp4_h_r_37')
// (7, 20, 'sp4_r_v_b_0')
// (8, 16, 'sp4_v_t_37')
// (8, 17, 'sp4_h_r_44')
// (8, 17, 'sp4_v_b_37')
// (8, 18, 'sp4_v_b_24')
// (8, 19, 'sp4_v_b_13')
// (8, 20, 'sp4_h_l_37')
// (8, 20, 'sp4_h_r_28')
// (8, 20, 'sp4_v_b_0')
// (9, 17, 'local_g1_1')
// (9, 17, 'lutff_3/in_3')
// (9, 17, 'sp4_h_l_44')
// (9, 17, 'sp4_h_r_9')
// (9, 17, 'sp4_r_v_b_47')
// (9, 18, 'sp4_r_v_b_34')
// (9, 19, 'local_g3_7')
// (9, 19, 'lutff_6/in_0')
// (9, 19, 'sp4_r_v_b_23')
// (9, 20, 'sp4_h_r_41')
// (9, 20, 'sp4_r_v_b_10')
// (10, 16, 'sp4_v_t_47')
// (10, 17, 'sp4_h_r_20')
// (10, 17, 'sp4_v_b_47')
// (10, 18, 'sp4_v_b_34')
// (10, 19, 'sp4_v_b_23')
// (10, 20, 'sp4_h_l_41')
// (10, 20, 'sp4_v_b_10')
// (11, 17, 'sp4_h_r_33')
// (12, 17, 'sp4_h_r_44')
// (13, 17, 'sp4_h_l_44')

wire n491;
// (2, 21, 'lutff_1/cout')
// (2, 21, 'lutff_2/in_3')

reg n492 = 0;
// (3, 0, 'logic_op_tnr_0')
// (3, 1, 'neigh_op_rgt_0')
// (3, 2, 'neigh_op_bnr_0')
// (4, 0, 'logic_op_top_0')
// (4, 1, 'lutff_0/out')
// (4, 2, 'neigh_op_bot_0')
// (5, 0, 'logic_op_tnl_0')
// (5, 1, 'local_g0_0')
// (5, 1, 'lutff_7/in_1')
// (5, 1, 'neigh_op_lft_0')
// (5, 2, 'neigh_op_bnl_0')

wire n493;
// (3, 0, 'logic_op_tnr_1')
// (3, 1, 'neigh_op_rgt_1')
// (3, 2, 'neigh_op_bnr_1')
// (4, 0, 'logic_op_top_1')
// (4, 1, 'lutff_1/out')
// (4, 2, 'neigh_op_bot_1')
// (5, 0, 'logic_op_tnl_1')
// (5, 1, 'neigh_op_lft_1')
// (5, 2, 'local_g3_1')
// (5, 2, 'lutff_5/in_3')
// (5, 2, 'neigh_op_bnl_1')

wire n494;
// (3, 0, 'logic_op_tnr_2')
// (3, 1, 'neigh_op_rgt_2')
// (3, 2, 'neigh_op_bnr_2')
// (4, 0, 'logic_op_top_2')
// (4, 1, 'lutff_2/out')
// (4, 2, 'neigh_op_bot_2')
// (5, 0, 'logic_op_tnl_2')
// (5, 1, 'local_g1_2')
// (5, 1, 'lutff_2/in_3')
// (5, 1, 'neigh_op_lft_2')
// (5, 2, 'neigh_op_bnl_2')

wire n495;
// (3, 0, 'logic_op_tnr_3')
// (3, 1, 'neigh_op_rgt_3')
// (3, 2, 'neigh_op_bnr_3')
// (4, 0, 'logic_op_top_3')
// (4, 1, 'lutff_3/out')
// (4, 2, 'local_g0_3')
// (4, 2, 'lutff_1/in_2')
// (4, 2, 'neigh_op_bot_3')
// (5, 0, 'logic_op_tnl_3')
// (5, 1, 'neigh_op_lft_3')
// (5, 2, 'neigh_op_bnl_3')

reg n496 = 0;
// (3, 0, 'logic_op_tnr_4')
// (3, 1, 'neigh_op_rgt_4')
// (3, 2, 'neigh_op_bnr_4')
// (4, 0, 'logic_op_top_4')
// (4, 1, 'lutff_4/out')
// (4, 2, 'neigh_op_bot_4')
// (5, 0, 'logic_op_tnl_4')
// (5, 1, 'local_g1_4')
// (5, 1, 'lutff_7/in_0')
// (5, 1, 'neigh_op_lft_4')
// (5, 2, 'neigh_op_bnl_4')

wire n497;
// (3, 0, 'logic_op_tnr_5')
// (3, 1, 'neigh_op_rgt_5')
// (3, 2, 'neigh_op_bnr_5')
// (4, 0, 'logic_op_top_5')
// (4, 1, 'lutff_5/out')
// (4, 2, 'neigh_op_bot_5')
// (5, 0, 'logic_op_tnl_5')
// (5, 1, 'neigh_op_lft_5')
// (5, 2, 'local_g2_5')
// (5, 2, 'lutff_7/in_0')
// (5, 2, 'neigh_op_bnl_5')

wire n498;
// (3, 0, 'logic_op_tnr_6')
// (3, 1, 'neigh_op_rgt_6')
// (3, 2, 'neigh_op_bnr_6')
// (4, 0, 'logic_op_top_6')
// (4, 1, 'lutff_6/out')
// (4, 2, 'neigh_op_bot_6')
// (5, 0, 'logic_op_tnl_6')
// (5, 1, 'local_g0_6')
// (5, 1, 'lutff_2/in_2')
// (5, 1, 'neigh_op_lft_6')
// (5, 2, 'neigh_op_bnl_6')

wire n499;
// (3, 0, 'logic_op_tnr_7')
// (3, 1, 'neigh_op_rgt_7')
// (3, 2, 'neigh_op_bnr_7')
// (4, 0, 'logic_op_top_7')
// (4, 1, 'lutff_7/out')
// (4, 1, 'sp4_r_v_b_15')
// (4, 2, 'neigh_op_bot_7')
// (4, 2, 'sp4_r_v_b_2')
// (5, 0, 'logic_op_tnl_7')
// (5, 0, 'span4_vert_15')
// (5, 1, 'neigh_op_lft_7')
// (5, 1, 'sp4_v_b_15')
// (5, 2, 'neigh_op_bnl_7')
// (5, 2, 'sp4_h_r_8')
// (5, 2, 'sp4_v_b_2')
// (6, 2, 'sp4_h_r_21')
// (7, 2, 'local_g2_0')
// (7, 2, 'lutff_0/in_0')
// (7, 2, 'sp4_h_r_32')
// (8, 2, 'sp4_h_r_45')
// (9, 2, 'sp4_h_l_45')

wire n500;
// (3, 1, 'local_g1_3')
// (3, 1, 'lutff_global/cen')
// (3, 1, 'sp4_h_r_11')
// (3, 2, 'local_g0_2')
// (3, 2, 'lutff_global/cen')
// (3, 2, 'sp4_h_r_2')
// (4, 1, 'sp4_h_r_22')
// (4, 2, 'sp4_h_r_15')
// (5, 1, 'sp4_h_r_35')
// (5, 2, 'sp4_h_r_26')
// (6, 1, 'sp4_h_r_46')
// (6, 2, 'sp4_h_r_39')
// (6, 2, 'sp4_r_v_b_40')
// (6, 3, 'neigh_op_tnr_0')
// (6, 3, 'sp4_r_v_b_29')
// (6, 3, 'sp4_r_v_b_45')
// (6, 4, 'neigh_op_rgt_0')
// (6, 4, 'sp4_r_v_b_16')
// (6, 4, 'sp4_r_v_b_32')
// (6, 5, 'neigh_op_bnr_0')
// (6, 5, 'sp4_r_v_b_21')
// (6, 5, 'sp4_r_v_b_5')
// (6, 6, 'sp4_r_v_b_8')
// (7, 1, 'sp4_h_l_46')
// (7, 1, 'sp4_v_t_40')
// (7, 2, 'sp4_h_l_39')
// (7, 2, 'sp4_v_b_40')
// (7, 2, 'sp4_v_t_45')
// (7, 3, 'neigh_op_top_0')
// (7, 3, 'sp4_v_b_29')
// (7, 3, 'sp4_v_b_45')
// (7, 4, 'lutff_0/out')
// (7, 4, 'sp4_v_b_16')
// (7, 4, 'sp4_v_b_32')
// (7, 5, 'neigh_op_bot_0')
// (7, 5, 'sp4_v_b_21')
// (7, 5, 'sp4_v_b_5')
// (7, 6, 'sp4_v_b_8')
// (8, 3, 'neigh_op_tnl_0')
// (8, 4, 'neigh_op_lft_0')
// (8, 5, 'neigh_op_bnl_0')

reg n501 = 0;
// (3, 1, 'neigh_op_tnr_0')
// (3, 2, 'neigh_op_rgt_0')
// (3, 3, 'neigh_op_bnr_0')
// (4, 1, 'local_g0_0')
// (4, 1, 'lutff_3/in_1')
// (4, 1, 'neigh_op_top_0')
// (4, 2, 'local_g3_0')
// (4, 2, 'lutff_0/out')
// (4, 2, 'lutff_3/in_2')
// (4, 3, 'neigh_op_bot_0')
// (5, 1, 'local_g2_0')
// (5, 1, 'lutff_3/in_3')
// (5, 1, 'neigh_op_tnl_0')
// (5, 2, 'neigh_op_lft_0')
// (5, 3, 'neigh_op_bnl_0')

wire n502;
// (3, 1, 'neigh_op_tnr_1')
// (3, 2, 'neigh_op_rgt_1')
// (3, 3, 'neigh_op_bnr_1')
// (4, 1, 'local_g0_1')
// (4, 1, 'lutff_1/in_0')
// (4, 1, 'neigh_op_top_1')
// (4, 2, 'lutff_1/out')
// (4, 3, 'neigh_op_bot_1')
// (5, 1, 'local_g3_1')
// (5, 1, 'lutff_5/in_3')
// (5, 1, 'neigh_op_tnl_1')
// (5, 2, 'neigh_op_lft_1')
// (5, 3, 'neigh_op_bnl_1')

wire n503;
// (3, 1, 'neigh_op_tnr_2')
// (3, 2, 'neigh_op_rgt_2')
// (3, 3, 'neigh_op_bnr_2')
// (4, 1, 'neigh_op_top_2')
// (4, 2, 'lutff_2/out')
// (4, 3, 'neigh_op_bot_2')
// (5, 1, 'local_g3_2')
// (5, 1, 'lutff_5/in_2')
// (5, 1, 'neigh_op_tnl_2')
// (5, 2, 'neigh_op_lft_2')
// (5, 3, 'neigh_op_bnl_2')

wire n504;
// (3, 1, 'neigh_op_tnr_3')
// (3, 2, 'neigh_op_rgt_3')
// (3, 3, 'neigh_op_bnr_3')
// (4, 1, 'neigh_op_top_3')
// (4, 2, 'lutff_3/out')
// (4, 3, 'local_g0_3')
// (4, 3, 'lutff_2/in_1')
// (4, 3, 'neigh_op_bot_3')
// (5, 1, 'neigh_op_tnl_3')
// (5, 2, 'neigh_op_lft_3')
// (5, 3, 'neigh_op_bnl_3')

wire n505;
// (3, 1, 'neigh_op_tnr_4')
// (3, 2, 'neigh_op_rgt_4')
// (3, 3, 'neigh_op_bnr_4')
// (4, 1, 'neigh_op_top_4')
// (4, 2, 'lutff_4/out')
// (4, 3, 'local_g1_4')
// (4, 3, 'lutff_3/in_0')
// (4, 3, 'neigh_op_bot_4')
// (5, 1, 'neigh_op_tnl_4')
// (5, 2, 'neigh_op_lft_4')
// (5, 3, 'neigh_op_bnl_4')

reg n506 = 0;
// (3, 1, 'neigh_op_tnr_5')
// (3, 2, 'neigh_op_rgt_5')
// (3, 2, 'sp4_r_v_b_42')
// (3, 3, 'neigh_op_bnr_5')
// (3, 3, 'sp4_r_v_b_31')
// (3, 4, 'sp4_r_v_b_18')
// (3, 5, 'sp4_r_v_b_7')
// (4, 1, 'neigh_op_top_5')
// (4, 1, 'sp4_v_t_42')
// (4, 2, 'lutff_5/out')
// (4, 2, 'sp4_r_v_b_43')
// (4, 2, 'sp4_v_b_42')
// (4, 3, 'local_g2_7')
// (4, 3, 'lutff_1/in_2')
// (4, 3, 'neigh_op_bot_5')
// (4, 3, 'sp4_r_v_b_30')
// (4, 3, 'sp4_v_b_31')
// (4, 4, 'sp4_r_v_b_19')
// (4, 4, 'sp4_v_b_18')
// (4, 5, 'sp4_r_v_b_6')
// (4, 5, 'sp4_v_b_7')
// (5, 1, 'neigh_op_tnl_5')
// (5, 1, 'sp4_v_t_43')
// (5, 2, 'neigh_op_lft_5')
// (5, 2, 'sp4_v_b_43')
// (5, 3, 'neigh_op_bnl_5')
// (5, 3, 'sp4_v_b_30')
// (5, 4, 'local_g0_3')
// (5, 4, 'lutff_2/in_3')
// (5, 4, 'lutff_4/in_1')
// (5, 4, 'sp4_v_b_19')
// (5, 5, 'sp4_v_b_6')

wire n507;
// (3, 1, 'neigh_op_tnr_6')
// (3, 2, 'neigh_op_rgt_6')
// (3, 3, 'neigh_op_bnr_6')
// (4, 1, 'neigh_op_top_6')
// (4, 2, 'lutff_6/out')
// (4, 3, 'local_g1_6')
// (4, 3, 'lutff_4/in_3')
// (4, 3, 'neigh_op_bot_6')
// (5, 1, 'neigh_op_tnl_6')
// (5, 2, 'neigh_op_lft_6')
// (5, 3, 'neigh_op_bnl_6')

wire n508;
// (3, 1, 'neigh_op_tnr_7')
// (3, 2, 'neigh_op_rgt_7')
// (3, 3, 'neigh_op_bnr_7')
// (4, 1, 'neigh_op_top_7')
// (4, 2, 'lutff_7/out')
// (4, 3, 'local_g1_7')
// (4, 3, 'lutff_4/in_2')
// (4, 3, 'neigh_op_bot_7')
// (5, 1, 'neigh_op_tnl_7')
// (5, 2, 'neigh_op_lft_7')
// (5, 3, 'neigh_op_bnl_7')

wire n509;
// (3, 1, 'sp4_r_v_b_42')
// (3, 2, 'sp4_r_v_b_31')
// (3, 3, 'sp4_r_v_b_18')
// (3, 4, 'sp4_r_v_b_7')
// (4, 0, 'span4_vert_42')
// (4, 1, 'sp4_r_v_b_23')
// (4, 1, 'sp4_v_b_42')
// (4, 2, 'local_g2_2')
// (4, 2, 'lutff_global/cen')
// (4, 2, 'sp4_r_v_b_10')
// (4, 2, 'sp4_v_b_31')
// (4, 3, 'local_g0_2')
// (4, 3, 'lutff_global/cen')
// (4, 3, 'sp4_v_b_18')
// (4, 4, 'sp4_h_r_2')
// (4, 4, 'sp4_v_b_7')
// (5, 0, 'span4_vert_23')
// (5, 1, 'sp4_v_b_23')
// (5, 2, 'local_g1_3')
// (5, 2, 'lutff_global/cen')
// (5, 2, 'sp4_h_r_11')
// (5, 2, 'sp4_h_r_5')
// (5, 2, 'sp4_v_b_10')
// (5, 4, 'sp4_h_r_15')
// (6, 2, 'sp4_h_r_16')
// (6, 2, 'sp4_h_r_22')
// (6, 4, 'sp4_h_r_26')
// (7, 2, 'local_g3_3')
// (7, 2, 'lutff_global/cen')
// (7, 2, 'sp4_h_r_29')
// (7, 2, 'sp4_h_r_35')
// (7, 4, 'sp4_h_r_39')
// (7, 5, 'neigh_op_tnr_5')
// (7, 5, 'sp4_r_v_b_39')
// (7, 6, 'neigh_op_rgt_5')
// (7, 6, 'sp4_r_v_b_26')
// (7, 7, 'neigh_op_bnr_5')
// (7, 7, 'sp4_r_v_b_15')
// (7, 8, 'sp4_r_v_b_2')
// (8, 2, 'sp4_h_r_40')
// (8, 2, 'sp4_h_r_46')
// (8, 3, 'sp4_r_v_b_46')
// (8, 4, 'sp4_h_l_39')
// (8, 4, 'sp4_r_v_b_35')
// (8, 4, 'sp4_v_t_39')
// (8, 5, 'neigh_op_top_5')
// (8, 5, 'sp4_r_v_b_22')
// (8, 5, 'sp4_v_b_39')
// (8, 6, 'lutff_5/out')
// (8, 6, 'sp4_r_v_b_11')
// (8, 6, 'sp4_v_b_26')
// (8, 7, 'neigh_op_bot_5')
// (8, 7, 'sp4_v_b_15')
// (8, 8, 'sp4_v_b_2')
// (9, 2, 'sp4_h_l_40')
// (9, 2, 'sp4_h_l_46')
// (9, 2, 'sp4_v_t_46')
// (9, 3, 'sp4_v_b_46')
// (9, 4, 'sp4_v_b_35')
// (9, 5, 'neigh_op_tnl_5')
// (9, 5, 'sp4_v_b_22')
// (9, 6, 'neigh_op_lft_5')
// (9, 6, 'sp4_v_b_11')
// (9, 7, 'neigh_op_bnl_5')

wire n510;
// (3, 2, 'neigh_op_tnr_0')
// (3, 3, 'neigh_op_rgt_0')
// (3, 3, 'sp4_h_r_5')
// (3, 4, 'neigh_op_bnr_0')
// (4, 2, 'local_g0_0')
// (4, 2, 'lutff_2/in_2')
// (4, 2, 'neigh_op_top_0')
// (4, 3, 'lutff_0/out')
// (4, 3, 'sp4_h_r_16')
// (4, 4, 'neigh_op_bot_0')
// (5, 2, 'neigh_op_tnl_0')
// (5, 3, 'local_g2_5')
// (5, 3, 'lutff_6/in_3')
// (5, 3, 'neigh_op_lft_0')
// (5, 3, 'sp4_h_r_29')
// (5, 4, 'neigh_op_bnl_0')
// (6, 3, 'sp4_h_r_40')
// (7, 3, 'sp4_h_l_40')

wire n511;
// (3, 2, 'neigh_op_tnr_1')
// (3, 3, 'neigh_op_rgt_1')
// (3, 4, 'neigh_op_bnr_1')
// (4, 2, 'local_g1_1')
// (4, 2, 'lutff_1/in_1')
// (4, 2, 'neigh_op_top_1')
// (4, 3, 'lutff_1/out')
// (4, 4, 'neigh_op_bot_1')
// (5, 2, 'neigh_op_tnl_1')
// (5, 3, 'neigh_op_lft_1')
// (5, 4, 'neigh_op_bnl_1')

wire n512;
// (3, 2, 'neigh_op_tnr_2')
// (3, 3, 'neigh_op_rgt_2')
// (3, 4, 'local_g0_2')
// (3, 4, 'lutff_6/in_2')
// (3, 4, 'neigh_op_bnr_2')
// (4, 2, 'neigh_op_top_2')
// (4, 3, 'lutff_2/out')
// (4, 4, 'neigh_op_bot_2')
// (5, 2, 'neigh_op_tnl_2')
// (5, 3, 'neigh_op_lft_2')
// (5, 4, 'neigh_op_bnl_2')

wire n513;
// (3, 2, 'neigh_op_tnr_3')
// (3, 3, 'neigh_op_rgt_3')
// (3, 4, 'neigh_op_bnr_3')
// (4, 2, 'local_g1_3')
// (4, 2, 'lutff_2/in_0')
// (4, 2, 'neigh_op_top_3')
// (4, 3, 'lutff_3/out')
// (4, 4, 'neigh_op_bot_3')
// (5, 2, 'neigh_op_tnl_3')
// (5, 3, 'local_g1_3')
// (5, 3, 'lutff_6/in_2')
// (5, 3, 'neigh_op_lft_3')
// (5, 4, 'neigh_op_bnl_3')

wire n514;
// (3, 2, 'neigh_op_tnr_4')
// (3, 3, 'local_g2_4')
// (3, 3, 'lutff_5/in_1')
// (3, 3, 'neigh_op_rgt_4')
// (3, 4, 'neigh_op_bnr_4')
// (4, 2, 'neigh_op_top_4')
// (4, 3, 'lutff_4/out')
// (4, 4, 'neigh_op_bot_4')
// (5, 2, 'neigh_op_tnl_4')
// (5, 3, 'neigh_op_lft_4')
// (5, 4, 'neigh_op_bnl_4')

reg n515 = 0;
// (3, 2, 'neigh_op_tnr_5')
// (3, 3, 'neigh_op_rgt_5')
// (3, 4, 'neigh_op_bnr_5')
// (4, 1, 'local_g2_3')
// (4, 1, 'lutff_2/in_3')
// (4, 1, 'sp4_r_v_b_35')
// (4, 2, 'neigh_op_top_5')
// (4, 2, 'sp4_r_v_b_22')
// (4, 2, 'sp4_r_v_b_38')
// (4, 3, 'lutff_5/out')
// (4, 3, 'sp4_r_v_b_11')
// (4, 3, 'sp4_r_v_b_27')
// (4, 4, 'neigh_op_bot_5')
// (4, 4, 'sp4_r_v_b_14')
// (4, 5, 'sp4_r_v_b_3')
// (5, 0, 'span4_vert_35')
// (5, 1, 'sp4_h_r_3')
// (5, 1, 'sp4_v_b_35')
// (5, 1, 'sp4_v_t_38')
// (5, 2, 'neigh_op_tnl_5')
// (5, 2, 'sp4_v_b_22')
// (5, 2, 'sp4_v_b_38')
// (5, 3, 'neigh_op_lft_5')
// (5, 3, 'sp4_v_b_11')
// (5, 3, 'sp4_v_b_27')
// (5, 4, 'neigh_op_bnl_5')
// (5, 4, 'sp4_v_b_14')
// (5, 5, 'sp4_v_b_3')
// (6, 1, 'sp4_h_r_14')
// (7, 1, 'local_g2_3')
// (7, 1, 'lutff_5/in_2')
// (7, 1, 'sp4_h_r_27')
// (8, 1, 'sp4_h_r_38')
// (9, 1, 'sp4_h_l_38')

reg n516 = 0;
// (3, 2, 'neigh_op_tnr_6')
// (3, 3, 'local_g3_6')
// (3, 3, 'lutff_3/in_2')
// (3, 3, 'neigh_op_rgt_6')
// (3, 4, 'neigh_op_bnr_6')
// (4, 2, 'local_g1_6')
// (4, 2, 'lutff_3/in_0')
// (4, 2, 'neigh_op_top_6')
// (4, 3, 'local_g2_6')
// (4, 3, 'lutff_1/in_3')
// (4, 3, 'lutff_6/out')
// (4, 4, 'neigh_op_bot_6')
// (5, 2, 'neigh_op_tnl_6')
// (5, 3, 'neigh_op_lft_6')
// (5, 4, 'neigh_op_bnl_6')

wire n517;
// (3, 2, 'neigh_op_tnr_7')
// (3, 3, 'neigh_op_rgt_7')
// (3, 4, 'neigh_op_bnr_7')
// (4, 2, 'neigh_op_top_7')
// (4, 3, 'local_g3_7')
// (4, 3, 'lutff_2/in_2')
// (4, 3, 'lutff_7/out')
// (4, 4, 'neigh_op_bot_7')
// (5, 2, 'neigh_op_tnl_7')
// (5, 3, 'neigh_op_lft_7')
// (5, 4, 'neigh_op_bnl_7')

wire n518;
// (3, 2, 'sp4_h_r_1')
// (4, 2, 'local_g1_4')
// (4, 2, 'lutff_7/in_2')
// (4, 2, 'sp4_h_r_12')
// (4, 2, 'sp4_h_r_3')
// (5, 2, 'local_g0_6')
// (5, 2, 'lutff_7/in_1')
// (5, 2, 'sp4_h_r_14')
// (5, 2, 'sp4_h_r_25')
// (6, 2, 'sp4_h_r_27')
// (6, 2, 'sp4_h_r_36')
// (7, 1, 'neigh_op_tnr_0')
// (7, 2, 'neigh_op_rgt_0')
// (7, 2, 'sp4_h_l_36')
// (7, 2, 'sp4_h_r_38')
// (7, 2, 'sp4_h_r_5')
// (7, 3, 'neigh_op_bnr_0')
// (8, 1, 'neigh_op_top_0')
// (8, 2, 'lutff_0/out')
// (8, 2, 'sp4_h_l_38')
// (8, 2, 'sp4_h_r_0')
// (8, 2, 'sp4_h_r_16')
// (8, 3, 'neigh_op_bot_0')
// (9, 1, 'neigh_op_tnl_0')
// (9, 2, 'neigh_op_lft_0')
// (9, 2, 'sp4_h_r_13')
// (9, 2, 'sp4_h_r_29')
// (9, 3, 'neigh_op_bnl_0')
// (10, 2, 'sp4_h_r_24')
// (10, 2, 'sp4_h_r_40')
// (11, 2, 'sp4_h_l_40')
// (11, 2, 'sp4_h_r_37')
// (12, 2, 'sp4_h_l_37')

wire n519;
// (3, 3, 'neigh_op_tnr_0')
// (3, 4, 'neigh_op_rgt_0')
// (3, 5, 'neigh_op_bnr_0')
// (4, 3, 'neigh_op_top_0')
// (4, 4, 'lutff_0/out')
// (4, 5, 'neigh_op_bot_0')
// (5, 3, 'local_g2_0')
// (5, 3, 'lutff_2/in_0')
// (5, 3, 'neigh_op_tnl_0')
// (5, 4, 'neigh_op_lft_0')
// (5, 5, 'neigh_op_bnl_0')

wire n520;
// (3, 3, 'neigh_op_tnr_1')
// (3, 4, 'neigh_op_rgt_1')
// (3, 5, 'neigh_op_bnr_1')
// (4, 3, 'neigh_op_top_1')
// (4, 4, 'local_g3_1')
// (4, 4, 'lutff_0/in_2')
// (4, 4, 'lutff_1/out')
// (4, 5, 'neigh_op_bot_1')
// (5, 3, 'neigh_op_tnl_1')
// (5, 4, 'neigh_op_lft_1')
// (5, 5, 'neigh_op_bnl_1')

wire n521;
// (3, 3, 'neigh_op_tnr_2')
// (3, 4, 'local_g3_2')
// (3, 4, 'lutff_6/in_1')
// (3, 4, 'neigh_op_rgt_2')
// (3, 5, 'neigh_op_bnr_2')
// (4, 3, 'neigh_op_top_2')
// (4, 4, 'lutff_2/out')
// (4, 5, 'neigh_op_bot_2')
// (5, 3, 'neigh_op_tnl_2')
// (5, 4, 'neigh_op_lft_2')
// (5, 5, 'neigh_op_bnl_2')

wire n522;
// (3, 3, 'neigh_op_tnr_3')
// (3, 4, 'neigh_op_rgt_3')
// (3, 5, 'neigh_op_bnr_3')
// (4, 3, 'neigh_op_top_3')
// (4, 4, 'lutff_3/out')
// (4, 4, 'sp4_r_v_b_39')
// (4, 5, 'local_g0_2')
// (4, 5, 'lutff_3/in_3')
// (4, 5, 'neigh_op_bot_3')
// (4, 5, 'sp4_r_v_b_26')
// (4, 6, 'sp4_r_v_b_15')
// (4, 7, 'sp4_r_v_b_2')
// (5, 3, 'neigh_op_tnl_3')
// (5, 3, 'sp4_v_t_39')
// (5, 4, 'neigh_op_lft_3')
// (5, 4, 'sp4_v_b_39')
// (5, 5, 'neigh_op_bnl_3')
// (5, 5, 'sp4_v_b_26')
// (5, 6, 'sp4_v_b_15')
// (5, 7, 'sp4_v_b_2')

wire n523;
// (3, 3, 'neigh_op_tnr_7')
// (3, 4, 'local_g2_7')
// (3, 4, 'lutff_6/in_3')
// (3, 4, 'neigh_op_rgt_7')
// (3, 5, 'neigh_op_bnr_7')
// (4, 3, 'neigh_op_top_7')
// (4, 4, 'lutff_7/out')
// (4, 5, 'neigh_op_bot_7')
// (5, 3, 'neigh_op_tnl_7')
// (5, 4, 'neigh_op_lft_7')
// (5, 5, 'neigh_op_bnl_7')

wire n524;
// (3, 4, 'local_g1_3')
// (3, 4, 'lutff_global/cen')
// (3, 4, 'sp4_h_r_11')
// (4, 4, 'sp4_h_r_22')
// (4, 5, 'local_g1_3')
// (4, 5, 'lutff_global/cen')
// (4, 5, 'sp12_h_r_1')
// (4, 5, 'sp4_h_r_11')
// (5, 4, 'sp4_h_r_35')
// (5, 5, 'local_g0_2')
// (5, 5, 'lutff_global/cen')
// (5, 5, 'sp12_h_r_2')
// (5, 5, 'sp4_h_r_22')
// (6, 4, 'neigh_op_tnr_7')
// (6, 4, 'sp4_h_r_46')
// (6, 5, 'neigh_op_rgt_7')
// (6, 5, 'sp12_h_r_5')
// (6, 5, 'sp4_h_r_35')
// (6, 5, 'sp4_r_v_b_46')
// (6, 6, 'neigh_op_bnr_7')
// (6, 6, 'sp4_r_v_b_35')
// (6, 7, 'sp4_r_v_b_22')
// (6, 8, 'sp4_r_v_b_11')
// (7, 4, 'neigh_op_top_7')
// (7, 4, 'sp4_h_l_46')
// (7, 4, 'sp4_v_t_46')
// (7, 5, 'lutff_7/out')
// (7, 5, 'sp12_h_r_6')
// (7, 5, 'sp4_h_r_46')
// (7, 5, 'sp4_v_b_46')
// (7, 6, 'neigh_op_bot_7')
// (7, 6, 'sp4_v_b_35')
// (7, 7, 'sp4_v_b_22')
// (7, 8, 'sp4_v_b_11')
// (8, 4, 'neigh_op_tnl_7')
// (8, 5, 'neigh_op_lft_7')
// (8, 5, 'sp12_h_r_9')
// (8, 5, 'sp4_h_l_46')
// (8, 6, 'neigh_op_bnl_7')
// (9, 5, 'sp12_h_r_10')
// (10, 5, 'sp12_h_r_13')
// (11, 5, 'sp12_h_r_14')
// (12, 5, 'sp12_h_r_17')
// (13, 5, 'sp12_h_r_18')
// (14, 5, 'sp12_h_r_21')
// (15, 5, 'sp12_h_r_22')
// (16, 5, 'sp12_h_l_22')

wire n525;
// (3, 4, 'local_g2_4')
// (3, 4, 'lutff_3/in_3')
// (3, 4, 'neigh_op_tnr_4')
// (3, 5, 'neigh_op_rgt_4')
// (3, 6, 'neigh_op_bnr_4')
// (4, 4, 'neigh_op_top_4')
// (4, 5, 'lutff_4/out')
// (4, 6, 'neigh_op_bot_4')
// (5, 4, 'neigh_op_tnl_4')
// (5, 5, 'neigh_op_lft_4')
// (5, 6, 'neigh_op_bnl_4')

wire n526;
// (3, 4, 'local_g3_0')
// (3, 4, 'lutff_1/in_2')
// (3, 4, 'neigh_op_tnr_0')
// (3, 5, 'neigh_op_rgt_0')
// (3, 6, 'neigh_op_bnr_0')
// (4, 4, 'neigh_op_top_0')
// (4, 5, 'lutff_0/out')
// (4, 6, 'neigh_op_bot_0')
// (5, 4, 'neigh_op_tnl_0')
// (5, 5, 'neigh_op_lft_0')
// (5, 6, 'neigh_op_bnl_0')

reg n527 = 0;
// (3, 4, 'neigh_op_tnr_1')
// (3, 5, 'neigh_op_rgt_1')
// (3, 6, 'neigh_op_bnr_1')
// (4, 3, 'sp4_r_v_b_43')
// (4, 4, 'neigh_op_top_1')
// (4, 4, 'sp4_r_v_b_30')
// (4, 5, 'lutff_1/out')
// (4, 5, 'sp4_r_v_b_19')
// (4, 6, 'neigh_op_bot_1')
// (4, 6, 'sp4_r_v_b_6')
// (5, 2, 'sp4_v_t_43')
// (5, 3, 'sp4_v_b_43')
// (5, 4, 'local_g2_1')
// (5, 4, 'lutff_7/in_0')
// (5, 4, 'neigh_op_tnl_1')
// (5, 4, 'sp4_v_b_30')
// (5, 5, 'local_g0_1')
// (5, 5, 'lutff_0/in_1')
// (5, 5, 'neigh_op_lft_1')
// (5, 5, 'sp4_v_b_19')
// (5, 6, 'neigh_op_bnl_1')
// (5, 6, 'sp4_h_r_6')
// (5, 6, 'sp4_v_b_6')
// (6, 6, 'sp4_h_r_19')
// (7, 6, 'local_g2_6')
// (7, 6, 'lutff_7/in_1')
// (7, 6, 'sp4_h_r_30')
// (8, 6, 'sp4_h_r_43')
// (9, 6, 'sp4_h_l_43')

wire n528;
// (3, 4, 'neigh_op_tnr_2')
// (3, 5, 'neigh_op_rgt_2')
// (3, 6, 'local_g0_2')
// (3, 6, 'lutff_5/in_3')
// (3, 6, 'neigh_op_bnr_2')
// (4, 4, 'neigh_op_top_2')
// (4, 5, 'lutff_2/out')
// (4, 6, 'neigh_op_bot_2')
// (5, 4, 'neigh_op_tnl_2')
// (5, 5, 'neigh_op_lft_2')
// (5, 6, 'neigh_op_bnl_2')

wire n529;
// (3, 4, 'neigh_op_tnr_3')
// (3, 5, 'neigh_op_rgt_3')
// (3, 5, 'sp4_h_r_11')
// (3, 6, 'neigh_op_bnr_3')
// (4, 4, 'neigh_op_top_3')
// (4, 5, 'local_g0_6')
// (4, 5, 'lutff_0/in_2')
// (4, 5, 'lutff_3/out')
// (4, 5, 'sp4_h_r_22')
// (4, 6, 'neigh_op_bot_3')
// (5, 4, 'neigh_op_tnl_3')
// (5, 5, 'neigh_op_lft_3')
// (5, 5, 'sp4_h_r_35')
// (5, 6, 'neigh_op_bnl_3')
// (6, 5, 'sp4_h_r_46')
// (7, 5, 'sp4_h_l_46')

wire n530;
// (3, 4, 'neigh_op_tnr_5')
// (3, 5, 'neigh_op_rgt_5')
// (3, 6, 'local_g0_5')
// (3, 6, 'lutff_2/in_3')
// (3, 6, 'lutff_7/in_2')
// (3, 6, 'neigh_op_bnr_5')
// (4, 4, 'neigh_op_top_5')
// (4, 5, 'lutff_5/out')
// (4, 6, 'neigh_op_bot_5')
// (5, 4, 'neigh_op_tnl_5')
// (5, 5, 'neigh_op_lft_5')
// (5, 6, 'neigh_op_bnl_5')

wire n531;
// (3, 4, 'neigh_op_tnr_6')
// (3, 5, 'neigh_op_rgt_6')
// (3, 6, 'neigh_op_bnr_6')
// (4, 4, 'neigh_op_top_6')
// (4, 5, 'lutff_6/out')
// (4, 6, 'neigh_op_bot_6')
// (5, 4, 'local_g3_6')
// (5, 4, 'lutff_0/in_3')
// (5, 4, 'neigh_op_tnl_6')
// (5, 5, 'neigh_op_lft_6')
// (5, 6, 'neigh_op_bnl_6')

wire n532;
// (3, 4, 'sp4_r_v_b_47')
// (3, 5, 'local_g2_2')
// (3, 5, 'lutff_global/cen')
// (3, 5, 'sp4_r_v_b_34')
// (3, 6, 'sp12_h_r_0')
// (3, 6, 'sp4_r_v_b_23')
// (3, 7, 'sp4_h_r_10')
// (3, 7, 'sp4_h_r_7')
// (3, 7, 'sp4_r_v_b_10')
// (4, 3, 'sp4_h_r_10')
// (4, 3, 'sp4_v_t_47')
// (4, 4, 'sp4_v_b_47')
// (4, 5, 'sp4_v_b_34')
// (4, 6, 'local_g1_3')
// (4, 6, 'lutff_global/cen')
// (4, 6, 'sp12_h_r_3')
// (4, 6, 'sp4_v_b_23')
// (4, 7, 'local_g0_2')
// (4, 7, 'lutff_global/cen')
// (4, 7, 'sp4_h_r_18')
// (4, 7, 'sp4_h_r_23')
// (4, 7, 'sp4_v_b_10')
// (5, 3, 'sp4_h_r_23')
// (5, 6, 'sp12_h_r_4')
// (5, 7, 'local_g2_2')
// (5, 7, 'lutff_global/cen')
// (5, 7, 'sp4_h_r_31')
// (5, 7, 'sp4_h_r_34')
// (6, 3, 'sp4_h_r_34')
// (6, 4, 'sp4_r_v_b_40')
// (6, 5, 'neigh_op_tnr_0')
// (6, 5, 'sp4_r_v_b_29')
// (6, 6, 'neigh_op_rgt_0')
// (6, 6, 'sp12_h_r_7')
// (6, 6, 'sp4_r_v_b_16')
// (6, 7, 'neigh_op_bnr_0')
// (6, 7, 'sp4_h_r_42')
// (6, 7, 'sp4_h_r_47')
// (6, 7, 'sp4_r_v_b_5')
// (7, 3, 'sp4_h_r_47')
// (7, 3, 'sp4_v_t_40')
// (7, 4, 'sp4_r_v_b_41')
// (7, 4, 'sp4_v_b_40')
// (7, 5, 'neigh_op_top_0')
// (7, 5, 'sp4_r_v_b_28')
// (7, 5, 'sp4_v_b_29')
// (7, 6, 'lutff_0/out')
// (7, 6, 'sp12_h_r_8')
// (7, 6, 'sp4_r_v_b_17')
// (7, 6, 'sp4_v_b_16')
// (7, 7, 'neigh_op_bot_0')
// (7, 7, 'sp4_h_l_42')
// (7, 7, 'sp4_h_l_47')
// (7, 7, 'sp4_h_r_11')
// (7, 7, 'sp4_r_v_b_4')
// (7, 7, 'sp4_v_b_5')
// (8, 3, 'sp4_h_l_47')
// (8, 3, 'sp4_v_t_41')
// (8, 4, 'sp4_v_b_41')
// (8, 5, 'neigh_op_tnl_0')
// (8, 5, 'sp4_v_b_28')
// (8, 6, 'neigh_op_lft_0')
// (8, 6, 'sp12_h_r_11')
// (8, 6, 'sp4_v_b_17')
// (8, 7, 'neigh_op_bnl_0')
// (8, 7, 'sp4_h_r_22')
// (8, 7, 'sp4_v_b_4')
// (9, 6, 'sp12_h_r_12')
// (9, 7, 'sp4_h_r_35')
// (10, 6, 'sp12_h_r_15')
// (10, 7, 'sp4_h_r_46')
// (11, 6, 'sp12_h_r_16')
// (11, 7, 'sp4_h_l_46')
// (12, 6, 'sp12_h_r_19')
// (13, 6, 'sp12_h_r_20')
// (14, 6, 'sp12_h_r_23')
// (15, 6, 'sp12_h_l_23')

wire n533;
// (3, 5, 'local_g2_0')
// (3, 5, 'lutff_4/in_2')
// (3, 5, 'neigh_op_tnr_0')
// (3, 6, 'neigh_op_rgt_0')
// (3, 7, 'neigh_op_bnr_0')
// (4, 5, 'neigh_op_top_0')
// (4, 6, 'lutff_0/out')
// (4, 7, 'neigh_op_bot_0')
// (5, 5, 'neigh_op_tnl_0')
// (5, 6, 'neigh_op_lft_0')
// (5, 7, 'neigh_op_bnl_0')

wire n534;
// (3, 5, 'local_g2_4')
// (3, 5, 'lutff_4/in_0')
// (3, 5, 'neigh_op_tnr_4')
// (3, 6, 'neigh_op_rgt_4')
// (3, 7, 'neigh_op_bnr_4')
// (4, 5, 'neigh_op_top_4')
// (4, 6, 'lutff_4/out')
// (4, 7, 'neigh_op_bot_4')
// (5, 5, 'neigh_op_tnl_4')
// (5, 6, 'neigh_op_lft_4')
// (5, 7, 'neigh_op_bnl_4')

wire n535;
// (3, 5, 'local_g2_7')
// (3, 5, 'lutff_5/in_2')
// (3, 5, 'neigh_op_tnr_7')
// (3, 6, 'neigh_op_rgt_7')
// (3, 7, 'neigh_op_bnr_7')
// (4, 5, 'neigh_op_top_7')
// (4, 6, 'lutff_7/out')
// (4, 7, 'neigh_op_bot_7')
// (5, 5, 'neigh_op_tnl_7')
// (5, 6, 'neigh_op_lft_7')
// (5, 7, 'neigh_op_bnl_7')

wire n536;
// (3, 5, 'local_g3_3')
// (3, 5, 'lutff_5/in_3')
// (3, 5, 'neigh_op_tnr_3')
// (3, 6, 'neigh_op_rgt_3')
// (3, 7, 'neigh_op_bnr_3')
// (4, 5, 'neigh_op_top_3')
// (4, 6, 'lutff_3/out')
// (4, 7, 'neigh_op_bot_3')
// (5, 5, 'neigh_op_tnl_3')
// (5, 6, 'neigh_op_lft_3')
// (5, 7, 'neigh_op_bnl_3')

reg n537 = 0;
// (3, 5, 'neigh_op_tnr_1')
// (3, 6, 'neigh_op_rgt_1')
// (3, 7, 'neigh_op_bnr_1')
// (4, 5, 'neigh_op_top_1')
// (4, 5, 'sp4_r_v_b_46')
// (4, 6, 'lutff_1/out')
// (4, 6, 'sp4_r_v_b_35')
// (4, 7, 'neigh_op_bot_1')
// (4, 7, 'sp4_r_v_b_22')
// (4, 8, 'sp4_r_v_b_11')
// (4, 9, 'sp4_r_v_b_46')
// (4, 10, 'sp4_r_v_b_35')
// (4, 11, 'sp4_r_v_b_22')
// (4, 12, 'sp4_r_v_b_11')
// (5, 4, 'sp4_v_t_46')
// (5, 5, 'neigh_op_tnl_1')
// (5, 5, 'sp4_v_b_46')
// (5, 6, 'neigh_op_lft_1')
// (5, 6, 'sp4_v_b_35')
// (5, 7, 'local_g3_1')
// (5, 7, 'lutff_5/in_3')
// (5, 7, 'neigh_op_bnl_1')
// (5, 7, 'sp4_v_b_22')
// (5, 8, 'sp4_v_b_11')
// (5, 8, 'sp4_v_t_46')
// (5, 9, 'local_g3_6')
// (5, 9, 'lutff_1/in_0')
// (5, 9, 'sp4_v_b_46')
// (5, 10, 'sp4_v_b_35')
// (5, 11, 'sp4_v_b_22')
// (5, 12, 'sp4_v_b_11')

wire n538;
// (3, 5, 'neigh_op_tnr_2')
// (3, 6, 'neigh_op_rgt_2')
// (3, 7, 'neigh_op_bnr_2')
// (4, 5, 'neigh_op_top_2')
// (4, 6, 'local_g3_2')
// (4, 6, 'lutff_2/out')
// (4, 6, 'lutff_7/in_0')
// (4, 7, 'neigh_op_bot_2')
// (5, 5, 'neigh_op_tnl_2')
// (5, 6, 'neigh_op_lft_2')
// (5, 7, 'neigh_op_bnl_2')

wire n539;
// (3, 5, 'neigh_op_tnr_5')
// (3, 6, 'local_g2_5')
// (3, 6, 'lutff_0/in_3')
// (3, 6, 'neigh_op_rgt_5')
// (3, 7, 'neigh_op_bnr_5')
// (4, 5, 'neigh_op_top_5')
// (4, 6, 'lutff_5/out')
// (4, 7, 'neigh_op_bot_5')
// (5, 5, 'neigh_op_tnl_5')
// (5, 6, 'neigh_op_lft_5')
// (5, 7, 'neigh_op_bnl_5')

wire n540;
// (3, 5, 'neigh_op_tnr_6')
// (3, 6, 'neigh_op_rgt_6')
// (3, 7, 'neigh_op_bnr_6')
// (4, 5, 'neigh_op_top_6')
// (4, 6, 'lutff_6/out')
// (4, 7, 'neigh_op_bot_6')
// (5, 5, 'neigh_op_tnl_6')
// (5, 6, 'neigh_op_lft_6')
// (5, 7, 'local_g2_6')
// (5, 7, 'lutff_6/in_0')
// (5, 7, 'neigh_op_bnl_6')

reg n541 = 0;
// (3, 5, 'sp4_h_r_0')
// (4, 4, 'neigh_op_tnr_4')
// (4, 5, 'neigh_op_rgt_4')
// (4, 5, 'sp4_h_r_13')
// (4, 6, 'neigh_op_bnr_4')
// (5, 4, 'local_g1_4')
// (5, 4, 'lutff_1/in_2')
// (5, 4, 'neigh_op_top_4')
// (5, 5, 'local_g2_4')
// (5, 5, 'lutff_0/in_0')
// (5, 5, 'lutff_4/out')
// (5, 5, 'sp4_h_r_24')
// (5, 6, 'neigh_op_bot_4')
// (6, 4, 'neigh_op_tnl_4')
// (6, 5, 'neigh_op_lft_4')
// (6, 5, 'sp4_h_r_37')
// (6, 6, 'neigh_op_bnl_4')
// (6, 6, 'sp4_r_v_b_37')
// (6, 7, 'sp4_r_v_b_24')
// (6, 8, 'sp4_r_v_b_13')
// (6, 9, 'sp4_r_v_b_0')
// (7, 5, 'sp4_h_l_37')
// (7, 5, 'sp4_v_t_37')
// (7, 6, 'local_g3_5')
// (7, 6, 'lutff_4/in_0')
// (7, 6, 'sp4_v_b_37')
// (7, 7, 'sp4_v_b_24')
// (7, 8, 'sp4_v_b_13')
// (7, 9, 'sp4_v_b_0')

reg n542 = 0;
// (3, 6, 'local_g3_0')
// (3, 6, 'lutff_1/in_0')
// (3, 6, 'neigh_op_tnr_0')
// (3, 7, 'local_g2_0')
// (3, 7, 'lutff_4/in_2')
// (3, 7, 'neigh_op_rgt_0')
// (3, 8, 'neigh_op_bnr_0')
// (4, 6, 'neigh_op_top_0')
// (4, 7, 'lutff_0/out')
// (4, 8, 'neigh_op_bot_0')
// (5, 6, 'local_g2_0')
// (5, 6, 'lutff_2/in_0')
// (5, 6, 'neigh_op_tnl_0')
// (5, 7, 'neigh_op_lft_0')
// (5, 8, 'local_g2_0')
// (5, 8, 'lutff_1/in_1')
// (5, 8, 'neigh_op_bnl_0')

wire n543;
// (3, 6, 'local_g3_3')
// (3, 6, 'lutff_2/in_0')
// (3, 6, 'neigh_op_tnr_3')
// (3, 7, 'neigh_op_rgt_3')
// (3, 8, 'neigh_op_bnr_3')
// (4, 6, 'neigh_op_top_3')
// (4, 7, 'lutff_3/out')
// (4, 8, 'neigh_op_bot_3')
// (5, 6, 'neigh_op_tnl_3')
// (5, 7, 'neigh_op_lft_3')
// (5, 8, 'neigh_op_bnl_3')

wire n544;
// (3, 6, 'local_g3_6')
// (3, 6, 'lutff_0/in_1')
// (3, 6, 'neigh_op_tnr_6')
// (3, 7, 'neigh_op_rgt_6')
// (3, 8, 'neigh_op_bnr_6')
// (4, 6, 'neigh_op_top_6')
// (4, 7, 'lutff_6/out')
// (4, 8, 'neigh_op_bot_6')
// (5, 6, 'neigh_op_tnl_6')
// (5, 7, 'neigh_op_lft_6')
// (5, 8, 'neigh_op_bnl_6')

reg n545 = 0;
// (3, 6, 'neigh_op_tnr_2')
// (3, 7, 'neigh_op_rgt_2')
// (3, 8, 'neigh_op_bnr_2')
// (4, 6, 'local_g0_2')
// (4, 6, 'lutff_4/in_2')
// (4, 6, 'neigh_op_top_2')
// (4, 7, 'local_g2_2')
// (4, 7, 'lutff_2/out')
// (4, 7, 'lutff_6/in_2')
// (4, 7, 'sp4_r_v_b_37')
// (4, 8, 'neigh_op_bot_2')
// (4, 8, 'sp4_r_v_b_24')
// (4, 9, 'sp4_r_v_b_13')
// (4, 10, 'sp4_r_v_b_0')
// (5, 6, 'neigh_op_tnl_2')
// (5, 6, 'sp4_v_t_37')
// (5, 7, 'neigh_op_lft_2')
// (5, 7, 'sp4_v_b_37')
// (5, 8, 'neigh_op_bnl_2')
// (5, 8, 'sp4_v_b_24')
// (5, 9, 'local_g0_5')
// (5, 9, 'lutff_0/in_3')
// (5, 9, 'sp4_v_b_13')
// (5, 10, 'sp4_v_b_0')

wire n546;
// (3, 6, 'neigh_op_tnr_5')
// (3, 7, 'neigh_op_rgt_5')
// (3, 8, 'neigh_op_bnr_5')
// (4, 6, 'local_g1_5')
// (4, 6, 'lutff_6/in_2')
// (4, 6, 'neigh_op_top_5')
// (4, 7, 'lutff_5/out')
// (4, 8, 'neigh_op_bot_5')
// (5, 6, 'neigh_op_tnl_5')
// (5, 7, 'neigh_op_lft_5')
// (5, 8, 'neigh_op_bnl_5')

wire n547;
// (3, 6, 'neigh_op_tnr_7')
// (3, 7, 'neigh_op_rgt_7')
// (3, 8, 'neigh_op_bnr_7')
// (4, 6, 'local_g1_7')
// (4, 6, 'lutff_5/in_3')
// (4, 6, 'neigh_op_top_7')
// (4, 7, 'lutff_7/out')
// (4, 8, 'neigh_op_bot_7')
// (5, 6, 'neigh_op_tnl_7')
// (5, 7, 'neigh_op_lft_7')
// (5, 8, 'neigh_op_bnl_7')

wire n548;
// (3, 7, 'neigh_op_tnr_1')
// (3, 8, 'neigh_op_rgt_1')
// (3, 9, 'neigh_op_bnr_1')
// (4, 7, 'neigh_op_top_1')
// (4, 8, 'local_g3_1')
// (4, 8, 'lutff_1/out')
// (4, 8, 'lutff_6/in_0')
// (4, 9, 'neigh_op_bot_1')
// (5, 7, 'neigh_op_tnl_1')
// (5, 8, 'neigh_op_lft_1')
// (5, 9, 'neigh_op_bnl_1')

wire n549;
// (3, 7, 'neigh_op_tnr_2')
// (3, 8, 'neigh_op_rgt_2')
// (3, 9, 'neigh_op_bnr_2')
// (4, 7, 'neigh_op_top_2')
// (4, 8, 'local_g0_2')
// (4, 8, 'lutff_2/out')
// (4, 8, 'lutff_7/in_3')
// (4, 9, 'neigh_op_bot_2')
// (5, 7, 'neigh_op_tnl_2')
// (5, 8, 'neigh_op_lft_2')
// (5, 9, 'neigh_op_bnl_2')

reg n550 = 0;
// (3, 7, 'neigh_op_tnr_3')
// (3, 8, 'neigh_op_rgt_3')
// (3, 9, 'neigh_op_bnr_3')
// (4, 7, 'neigh_op_top_3')
// (4, 8, 'lutff_3/out')
// (4, 8, 'sp4_h_r_6')
// (4, 9, 'neigh_op_bot_3')
// (5, 7, 'neigh_op_tnl_3')
// (5, 8, 'neigh_op_lft_3')
// (5, 8, 'sp4_h_r_19')
// (5, 9, 'neigh_op_bnl_3')
// (6, 8, 'sp4_h_r_30')
// (7, 5, 'sp4_r_v_b_43')
// (7, 6, 'sp4_r_v_b_30')
// (7, 7, 'local_g3_3')
// (7, 7, 'lutff_5/in_3')
// (7, 7, 'sp4_r_v_b_19')
// (7, 8, 'sp4_h_r_43')
// (7, 8, 'sp4_r_v_b_6')
// (8, 4, 'sp4_v_t_43')
// (8, 5, 'sp4_v_b_43')
// (8, 6, 'sp4_v_b_30')
// (8, 7, 'sp4_v_b_19')
// (8, 8, 'sp4_h_l_43')
// (8, 8, 'sp4_v_b_6')

reg n551 = 0;
// (3, 7, 'neigh_op_tnr_4')
// (3, 8, 'neigh_op_rgt_4')
// (3, 9, 'neigh_op_bnr_4')
// (4, 7, 'neigh_op_top_4')
// (4, 8, 'lutff_4/out')
// (4, 9, 'neigh_op_bot_4')
// (5, 7, 'neigh_op_tnl_4')
// (5, 8, 'local_g0_4')
// (5, 8, 'lutff_6/in_2')
// (5, 8, 'neigh_op_lft_4')
// (5, 9, 'neigh_op_bnl_4')

wire n552;
// (3, 7, 'neigh_op_tnr_5')
// (3, 8, 'neigh_op_rgt_5')
// (3, 9, 'neigh_op_bnr_5')
// (4, 7, 'neigh_op_top_5')
// (4, 8, 'lutff_5/out')
// (4, 9, 'neigh_op_bot_5')
// (5, 7, 'local_g2_5')
// (5, 7, 'lutff_6/in_3')
// (5, 7, 'neigh_op_tnl_5')
// (5, 8, 'neigh_op_lft_5')
// (5, 9, 'neigh_op_bnl_5')

wire n553;
// (3, 7, 'neigh_op_tnr_6')
// (3, 8, 'neigh_op_rgt_6')
// (3, 9, 'neigh_op_bnr_6')
// (4, 7, 'neigh_op_top_6')
// (4, 8, 'local_g1_6')
// (4, 8, 'lutff_6/out')
// (4, 8, 'lutff_7/in_2')
// (4, 9, 'neigh_op_bot_6')
// (5, 7, 'neigh_op_tnl_6')
// (5, 8, 'neigh_op_lft_6')
// (5, 9, 'neigh_op_bnl_6')

wire n554;
// (3, 7, 'neigh_op_tnr_7')
// (3, 8, 'neigh_op_rgt_7')
// (3, 9, 'neigh_op_bnr_7')
// (4, 7, 'neigh_op_top_7')
// (4, 8, 'local_g1_7')
// (4, 8, 'lutff_5/in_1')
// (4, 8, 'lutff_7/out')
// (4, 9, 'neigh_op_bot_7')
// (5, 7, 'neigh_op_tnl_7')
// (5, 8, 'neigh_op_lft_7')
// (5, 9, 'neigh_op_bnl_7')

wire n555;
// (3, 8, 'lutff_1/cout')
// (3, 8, 'lutff_2/in_3')

wire n556;
// (3, 8, 'lutff_2/cout')
// (3, 8, 'lutff_3/in_3')

reg n557 = 0;
// (3, 8, 'neigh_op_tnr_1')
// (3, 9, 'neigh_op_rgt_1')
// (3, 10, 'neigh_op_bnr_1')
// (4, 8, 'neigh_op_top_1')
// (4, 9, 'lutff_1/out')
// (4, 10, 'neigh_op_bot_1')
// (5, 8, 'local_g3_1')
// (5, 8, 'lutff_3/in_3')
// (5, 8, 'neigh_op_tnl_1')
// (5, 9, 'neigh_op_lft_1')
// (5, 10, 'neigh_op_bnl_1')

reg n558 = 0;
// (3, 8, 'neigh_op_tnr_2')
// (3, 9, 'neigh_op_rgt_2')
// (3, 10, 'neigh_op_bnr_2')
// (4, 8, 'neigh_op_top_2')
// (4, 9, 'lutff_2/out')
// (4, 10, 'neigh_op_bot_2')
// (5, 8, 'local_g3_2')
// (5, 8, 'lutff_5/in_2')
// (5, 8, 'neigh_op_tnl_2')
// (5, 9, 'neigh_op_lft_2')
// (5, 10, 'neigh_op_bnl_2')

wire n559;
// (3, 8, 'neigh_op_tnr_3')
// (3, 9, 'neigh_op_rgt_3')
// (3, 10, 'neigh_op_bnr_3')
// (4, 8, 'local_g0_3')
// (4, 8, 'lutff_3/in_2')
// (4, 8, 'lutff_4/in_3')
// (4, 8, 'neigh_op_top_3')
// (4, 9, 'local_g2_3')
// (4, 9, 'lutff_1/in_2')
// (4, 9, 'lutff_2/in_3')
// (4, 9, 'lutff_3/out')
// (4, 9, 'lutff_4/in_3')
// (4, 9, 'lutff_5/in_0')
// (4, 9, 'lutff_6/in_1')
// (4, 10, 'neigh_op_bot_3')
// (5, 8, 'local_g2_3')
// (5, 8, 'lutff_0/in_3')
// (5, 8, 'neigh_op_tnl_3')
// (5, 9, 'neigh_op_lft_3')
// (5, 10, 'neigh_op_bnl_3')

reg n560 = 0;
// (3, 8, 'neigh_op_tnr_4')
// (3, 9, 'neigh_op_rgt_4')
// (3, 10, 'neigh_op_bnr_4')
// (4, 8, 'neigh_op_top_4')
// (4, 9, 'lutff_4/out')
// (4, 10, 'neigh_op_bot_4')
// (5, 8, 'neigh_op_tnl_4')
// (5, 9, 'local_g1_4')
// (5, 9, 'lutff_4/in_1')
// (5, 9, 'neigh_op_lft_4')
// (5, 10, 'neigh_op_bnl_4')

reg n561 = 0;
// (3, 8, 'neigh_op_tnr_5')
// (3, 9, 'neigh_op_rgt_5')
// (3, 10, 'neigh_op_bnr_5')
// (4, 8, 'neigh_op_top_5')
// (4, 9, 'lutff_5/out')
// (4, 10, 'neigh_op_bot_5')
// (5, 8, 'neigh_op_tnl_5')
// (5, 9, 'local_g1_5')
// (5, 9, 'lutff_7/in_1')
// (5, 9, 'neigh_op_lft_5')
// (5, 10, 'neigh_op_bnl_5')

reg n562 = 0;
// (3, 8, 'neigh_op_tnr_6')
// (3, 9, 'neigh_op_rgt_6')
// (3, 10, 'neigh_op_bnr_6')
// (4, 8, 'neigh_op_top_6')
// (4, 9, 'lutff_6/out')
// (4, 10, 'neigh_op_bot_6')
// (5, 8, 'neigh_op_tnl_6')
// (5, 9, 'local_g1_6')
// (5, 9, 'lutff_6/in_3')
// (5, 9, 'neigh_op_lft_6')
// (5, 10, 'neigh_op_bnl_6')

wire n563;
// (3, 8, 'neigh_op_tnr_7')
// (3, 9, 'local_g3_7')
// (3, 9, 'lutff_5/in_1')
// (3, 9, 'neigh_op_rgt_7')
// (3, 10, 'neigh_op_bnr_7')
// (4, 8, 'neigh_op_top_7')
// (4, 9, 'lutff_7/out')
// (4, 10, 'neigh_op_bot_7')
// (5, 8, 'neigh_op_tnl_7')
// (5, 9, 'neigh_op_lft_7')
// (5, 10, 'neigh_op_bnl_7')

wire n564;
// (3, 8, 'sp4_h_r_7')
// (4, 8, 'sp4_h_r_18')
// (4, 9, 'sp4_h_r_6')
// (4, 12, 'sp4_h_r_6')
// (5, 6, 'local_g1_2')
// (5, 6, 'lutff_5/in_2')
// (5, 6, 'lutff_6/in_3')
// (5, 6, 'sp4_h_r_2')
// (5, 8, 'local_g3_7')
// (5, 8, 'lutff_1/in_3')
// (5, 8, 'lutff_4/in_0')
// (5, 8, 'lutff_7/in_1')
// (5, 8, 'sp4_h_r_31')
// (5, 9, 'local_g0_3')
// (5, 9, 'lutff_0/in_1')
// (5, 9, 'lutff_1/in_2')
// (5, 9, 'lutff_3/in_0')
// (5, 9, 'sp4_h_r_19')
// (5, 12, 'local_g0_3')
// (5, 12, 'lutff_0/in_1')
// (5, 12, 'sp4_h_r_19')
// (6, 5, 'neigh_op_tnr_5')
// (6, 5, 'sp4_r_v_b_39')
// (6, 6, 'neigh_op_rgt_5')
// (6, 6, 'sp4_h_r_15')
// (6, 6, 'sp4_r_v_b_26')
// (6, 6, 'sp4_r_v_b_42')
// (6, 7, 'neigh_op_bnr_5')
// (6, 7, 'sp4_r_v_b_15')
// (6, 7, 'sp4_r_v_b_31')
// (6, 7, 'sp4_r_v_b_41')
// (6, 8, 'sp4_h_r_42')
// (6, 8, 'sp4_r_v_b_18')
// (6, 8, 'sp4_r_v_b_2')
// (6, 8, 'sp4_r_v_b_28')
// (6, 9, 'sp4_h_r_30')
// (6, 9, 'sp4_r_v_b_17')
// (6, 9, 'sp4_r_v_b_7')
// (6, 10, 'sp4_r_v_b_4')
// (6, 10, 'sp4_r_v_b_47')
// (6, 11, 'sp4_r_v_b_34')
// (6, 11, 'sp4_r_v_b_41')
// (6, 12, 'sp4_h_r_30')
// (6, 12, 'sp4_r_v_b_23')
// (6, 12, 'sp4_r_v_b_28')
// (6, 13, 'sp4_r_v_b_10')
// (6, 13, 'sp4_r_v_b_17')
// (6, 14, 'sp4_r_v_b_4')
// (7, 0, 'span12_vert_21')
// (7, 1, 'sp12_v_b_21')
// (7, 2, 'sp12_v_b_18')
// (7, 3, 'sp12_v_b_17')
// (7, 3, 'sp4_r_v_b_46')
// (7, 4, 'sp12_v_b_14')
// (7, 4, 'sp4_r_v_b_35')
// (7, 4, 'sp4_v_t_39')
// (7, 5, 'neigh_op_top_5')
// (7, 5, 'sp12_v_b_13')
// (7, 5, 'sp4_r_v_b_22')
// (7, 5, 'sp4_r_v_b_38')
// (7, 5, 'sp4_v_b_39')
// (7, 5, 'sp4_v_t_42')
// (7, 6, 'lutff_5/out')
// (7, 6, 'sp12_v_b_10')
// (7, 6, 'sp4_h_r_10')
// (7, 6, 'sp4_h_r_26')
// (7, 6, 'sp4_r_v_b_11')
// (7, 6, 'sp4_r_v_b_27')
// (7, 6, 'sp4_r_v_b_43')
// (7, 6, 'sp4_v_b_26')
// (7, 6, 'sp4_v_b_42')
// (7, 6, 'sp4_v_t_41')
// (7, 7, 'local_g1_5')
// (7, 7, 'lutff_3/in_3')
// (7, 7, 'neigh_op_bot_5')
// (7, 7, 'sp12_v_b_9')
// (7, 7, 'sp4_r_v_b_14')
// (7, 7, 'sp4_r_v_b_30')
// (7, 7, 'sp4_r_v_b_46')
// (7, 7, 'sp4_v_b_15')
// (7, 7, 'sp4_v_b_31')
// (7, 7, 'sp4_v_b_41')
// (7, 8, 'sp12_v_b_6')
// (7, 8, 'sp4_h_l_42')
// (7, 8, 'sp4_r_v_b_19')
// (7, 8, 'sp4_r_v_b_3')
// (7, 8, 'sp4_r_v_b_35')
// (7, 8, 'sp4_v_b_18')
// (7, 8, 'sp4_v_b_2')
// (7, 8, 'sp4_v_b_28')
// (7, 9, 'sp12_v_b_5')
// (7, 9, 'sp4_h_r_43')
// (7, 9, 'sp4_r_v_b_22')
// (7, 9, 'sp4_r_v_b_43')
// (7, 9, 'sp4_r_v_b_6')
// (7, 9, 'sp4_v_b_17')
// (7, 9, 'sp4_v_b_7')
// (7, 9, 'sp4_v_t_47')
// (7, 10, 'sp12_v_b_2')
// (7, 10, 'sp4_r_v_b_11')
// (7, 10, 'sp4_r_v_b_30')
// (7, 10, 'sp4_v_b_4')
// (7, 10, 'sp4_v_b_47')
// (7, 10, 'sp4_v_t_41')
// (7, 11, 'local_g3_1')
// (7, 11, 'lutff_1/in_1')
// (7, 11, 'lutff_5/in_1')
// (7, 11, 'sp12_v_b_1')
// (7, 11, 'sp4_r_v_b_19')
// (7, 11, 'sp4_v_b_34')
// (7, 11, 'sp4_v_b_41')
// (7, 12, 'sp4_h_r_43')
// (7, 12, 'sp4_r_v_b_6')
// (7, 12, 'sp4_v_b_23')
// (7, 12, 'sp4_v_b_28')
// (7, 13, 'local_g0_2')
// (7, 13, 'lutff_2/in_2')
// (7, 13, 'lutff_3/in_1')
// (7, 13, 'lutff_5/in_1')
// (7, 13, 'lutff_6/in_0')
// (7, 13, 'sp4_v_b_10')
// (7, 13, 'sp4_v_b_17')
// (7, 14, 'local_g1_4')
// (7, 14, 'lutff_1/in_2')
// (7, 14, 'sp4_v_b_4')
// (8, 2, 'sp4_v_t_46')
// (8, 3, 'sp4_v_b_46')
// (8, 4, 'sp4_v_b_35')
// (8, 4, 'sp4_v_t_38')
// (8, 5, 'neigh_op_tnl_5')
// (8, 5, 'sp4_v_b_22')
// (8, 5, 'sp4_v_b_38')
// (8, 5, 'sp4_v_t_43')
// (8, 6, 'neigh_op_lft_5')
// (8, 6, 'sp4_h_r_23')
// (8, 6, 'sp4_h_r_39')
// (8, 6, 'sp4_v_b_11')
// (8, 6, 'sp4_v_b_27')
// (8, 6, 'sp4_v_b_43')
// (8, 6, 'sp4_v_t_46')
// (8, 7, 'neigh_op_bnl_5')
// (8, 7, 'sp4_r_v_b_42')
// (8, 7, 'sp4_v_b_14')
// (8, 7, 'sp4_v_b_30')
// (8, 7, 'sp4_v_b_46')
// (8, 8, 'sp4_r_v_b_31')
// (8, 8, 'sp4_v_b_19')
// (8, 8, 'sp4_v_b_3')
// (8, 8, 'sp4_v_b_35')
// (8, 8, 'sp4_v_t_43')
// (8, 9, 'sp4_h_l_43')
// (8, 9, 'sp4_r_v_b_18')
// (8, 9, 'sp4_v_b_22')
// (8, 9, 'sp4_v_b_43')
// (8, 9, 'sp4_v_b_6')
// (8, 10, 'local_g0_3')
// (8, 10, 'lutff_0/in_3')
// (8, 10, 'lutff_1/in_2')
// (8, 10, 'lutff_3/in_0')
// (8, 10, 'sp4_r_v_b_7')
// (8, 10, 'sp4_v_b_11')
// (8, 10, 'sp4_v_b_30')
// (8, 11, 'local_g1_3')
// (8, 11, 'lutff_0/in_0')
// (8, 11, 'sp4_r_v_b_38')
// (8, 11, 'sp4_v_b_19')
// (8, 12, 'sp4_h_l_43')
// (8, 12, 'sp4_r_v_b_27')
// (8, 12, 'sp4_v_b_6')
// (8, 13, 'sp4_r_v_b_14')
// (8, 14, 'sp4_r_v_b_3')
// (9, 6, 'sp4_h_l_39')
// (9, 6, 'sp4_h_r_34')
// (9, 6, 'sp4_v_t_42')
// (9, 7, 'sp4_v_b_42')
// (9, 8, 'sp4_v_b_31')
// (9, 9, 'sp4_v_b_18')
// (9, 10, 'sp4_v_b_7')
// (9, 10, 'sp4_v_t_38')
// (9, 11, 'local_g2_6')
// (9, 11, 'lutff_2/in_2')
// (9, 11, 'lutff_4/in_2')
// (9, 11, 'sp4_v_b_38')
// (9, 12, 'sp4_v_b_27')
// (9, 13, 'sp4_v_b_14')
// (9, 14, 'sp4_v_b_3')
// (10, 6, 'sp4_h_r_47')
// (11, 6, 'sp4_h_l_47')

reg n565 = 0;
// (3, 9, 'local_g2_0')
// (3, 9, 'lutff_0/in_2')
// (3, 9, 'neigh_op_tnr_0')
// (3, 10, 'neigh_op_rgt_0')
// (3, 11, 'neigh_op_bnr_0')
// (4, 9, 'local_g1_0')
// (4, 9, 'lutff_7/in_2')
// (4, 9, 'neigh_op_top_0')
// (4, 10, 'lutff_0/out')
// (4, 10, 'sp4_h_r_0')
// (4, 11, 'neigh_op_bot_0')
// (5, 9, 'local_g3_0')
// (5, 9, 'lutff_2/in_1')
// (5, 9, 'neigh_op_tnl_0')
// (5, 10, 'neigh_op_lft_0')
// (5, 10, 'sp4_h_r_13')
// (5, 11, 'neigh_op_bnl_0')
// (6, 10, 'sp4_h_r_24')
// (7, 10, 'sp4_h_r_37')
// (8, 10, 'sp4_h_l_37')
// (8, 10, 'sp4_h_r_8')
// (9, 10, 'local_g1_5')
// (9, 10, 'lutff_0/in_2')
// (9, 10, 'sp4_h_r_21')
// (10, 10, 'sp4_h_r_32')
// (11, 10, 'sp4_h_r_45')
// (12, 10, 'sp4_h_l_45')

reg n566 = 0;
// (3, 9, 'local_g2_3')
// (3, 9, 'lutff_1/in_2')
// (3, 9, 'neigh_op_tnr_3')
// (3, 10, 'neigh_op_rgt_3')
// (3, 11, 'neigh_op_bnr_3')
// (4, 8, 'sp4_r_v_b_47')
// (4, 9, 'neigh_op_top_3')
// (4, 9, 'sp4_r_v_b_34')
// (4, 10, 'lutff_3/out')
// (4, 10, 'sp4_r_v_b_23')
// (4, 11, 'neigh_op_bot_3')
// (4, 11, 'sp4_r_v_b_10')
// (5, 7, 'sp4_v_t_47')
// (5, 8, 'sp4_v_b_47')
// (5, 9, 'neigh_op_tnl_3')
// (5, 9, 'sp4_v_b_34')
// (5, 10, 'local_g0_3')
// (5, 10, 'lutff_2/in_1')
// (5, 10, 'neigh_op_lft_3')
// (5, 10, 'sp4_v_b_23')
// (5, 11, 'neigh_op_bnl_3')
// (5, 11, 'sp4_h_r_10')
// (5, 11, 'sp4_v_b_10')
// (6, 11, 'sp4_h_r_23')
// (7, 11, 'sp4_h_r_34')
// (8, 11, 'local_g3_7')
// (8, 11, 'lutff_1/in_3')
// (8, 11, 'sp4_h_r_47')
// (9, 11, 'sp4_h_l_47')

reg n567 = 0;
// (3, 9, 'local_g2_7')
// (3, 9, 'lutff_3/in_2')
// (3, 9, 'neigh_op_tnr_7')
// (3, 10, 'neigh_op_rgt_7')
// (3, 10, 'sp4_h_r_3')
// (3, 11, 'neigh_op_bnr_7')
// (4, 8, 'sp4_r_v_b_39')
// (4, 9, 'neigh_op_top_7')
// (4, 9, 'sp4_r_v_b_26')
// (4, 10, 'lutff_7/out')
// (4, 10, 'sp4_h_r_14')
// (4, 10, 'sp4_r_v_b_15')
// (4, 11, 'neigh_op_bot_7')
// (4, 11, 'sp4_r_v_b_2')
// (5, 7, 'sp4_v_t_39')
// (5, 8, 'sp4_v_b_39')
// (5, 9, 'neigh_op_tnl_7')
// (5, 9, 'sp4_v_b_26')
// (5, 10, 'neigh_op_lft_7')
// (5, 10, 'sp4_h_r_27')
// (5, 10, 'sp4_v_b_15')
// (5, 11, 'neigh_op_bnl_7')
// (5, 11, 'sp4_h_r_2')
// (5, 11, 'sp4_v_b_2')
// (6, 10, 'sp4_h_r_38')
// (6, 11, 'sp4_h_r_15')
// (7, 10, 'local_g0_3')
// (7, 10, 'lutff_1/in_0')
// (7, 10, 'sp4_h_l_38')
// (7, 10, 'sp4_h_r_11')
// (7, 11, 'local_g3_2')
// (7, 11, 'lutff_2/in_3')
// (7, 11, 'sp4_h_r_26')
// (8, 10, 'sp4_h_r_22')
// (8, 11, 'sp4_h_r_39')
// (9, 10, 'sp4_h_r_35')
// (9, 11, 'sp4_h_l_39')
// (10, 10, 'sp4_h_r_46')
// (11, 10, 'sp4_h_l_46')

reg n568 = 0;
// (3, 9, 'local_g3_2')
// (3, 9, 'lutff_2/in_1')
// (3, 9, 'neigh_op_tnr_2')
// (3, 10, 'neigh_op_rgt_2')
// (3, 11, 'neigh_op_bnr_2')
// (4, 9, 'neigh_op_top_2')
// (4, 10, 'lutff_2/out')
// (4, 10, 'sp4_h_r_4')
// (4, 11, 'neigh_op_bot_2')
// (5, 9, 'local_g3_2')
// (5, 9, 'lutff_5/in_2')
// (5, 9, 'neigh_op_tnl_2')
// (5, 10, 'neigh_op_lft_2')
// (5, 10, 'sp4_h_r_17')
// (5, 11, 'neigh_op_bnl_2')
// (6, 10, 'sp4_h_r_28')
// (7, 10, 'sp4_h_r_41')
// (8, 10, 'local_g1_0')
// (8, 10, 'lutff_7/in_2')
// (8, 10, 'sp4_h_l_41')
// (8, 10, 'sp4_h_r_0')
// (9, 10, 'sp4_h_r_13')
// (10, 10, 'sp4_h_r_24')
// (11, 10, 'sp4_h_r_37')
// (12, 10, 'sp4_h_l_37')

wire n569;
// (3, 9, 'lutff_0/cout')
// (3, 9, 'lutff_1/in_3')

wire n570;
// (3, 9, 'lutff_1/cout')
// (3, 9, 'lutff_2/in_3')

wire n571;
// (3, 9, 'lutff_2/cout')
// (3, 9, 'lutff_3/in_3')

wire n572;
// (3, 9, 'lutff_3/cout')
// (3, 9, 'lutff_4/in_3')

reg n573 = 0;
// (3, 9, 'neigh_op_tnr_1')
// (3, 9, 'sp4_r_v_b_47')
// (3, 10, 'neigh_op_rgt_1')
// (3, 10, 'sp4_r_v_b_34')
// (3, 11, 'neigh_op_bnr_1')
// (3, 11, 'sp4_r_v_b_23')
// (3, 12, 'local_g2_2')
// (3, 12, 'lutff_3/in_3')
// (3, 12, 'sp4_r_v_b_10')
// (4, 7, 'sp4_r_v_b_38')
// (4, 8, 'sp4_h_r_10')
// (4, 8, 'sp4_r_v_b_27')
// (4, 8, 'sp4_v_t_47')
// (4, 9, 'neigh_op_top_1')
// (4, 9, 'sp4_r_v_b_14')
// (4, 9, 'sp4_v_b_47')
// (4, 10, 'lutff_1/out')
// (4, 10, 'sp4_r_v_b_3')
// (4, 10, 'sp4_v_b_34')
// (4, 11, 'neigh_op_bot_1')
// (4, 11, 'sp4_v_b_23')
// (4, 12, 'sp4_v_b_10')
// (5, 6, 'sp4_h_r_8')
// (5, 6, 'sp4_v_t_38')
// (5, 7, 'sp4_v_b_38')
// (5, 8, 'sp4_h_r_23')
// (5, 8, 'sp4_v_b_27')
// (5, 9, 'neigh_op_tnl_1')
// (5, 9, 'sp4_v_b_14')
// (5, 10, 'neigh_op_lft_1')
// (5, 10, 'sp4_v_b_3')
// (5, 11, 'neigh_op_bnl_1')
// (6, 6, 'sp4_h_r_21')
// (6, 8, 'sp4_h_r_34')
// (7, 6, 'sp4_h_r_32')
// (7, 8, 'sp4_h_r_47')
// (8, 6, 'sp4_h_r_45')
// (8, 7, 'sp4_r_v_b_45')
// (8, 8, 'sp4_h_l_47')
// (8, 8, 'sp4_h_r_6')
// (8, 8, 'sp4_r_v_b_32')
// (8, 9, 'sp4_r_v_b_21')
// (8, 10, 'sp4_r_v_b_8')
// (9, 6, 'sp4_h_l_45')
// (9, 6, 'sp4_v_t_45')
// (9, 7, 'sp4_v_b_45')
// (9, 8, 'local_g1_3')
// (9, 8, 'lutff_1/in_3')
// (9, 8, 'sp4_h_r_19')
// (9, 8, 'sp4_v_b_32')
// (9, 9, 'local_g0_5')
// (9, 9, 'lutff_4/in_3')
// (9, 9, 'sp4_v_b_21')
// (9, 10, 'sp4_v_b_8')
// (10, 8, 'sp4_h_r_30')
// (11, 8, 'sp4_h_r_43')
// (12, 8, 'sp4_h_l_43')

reg n574 = 0;
// (3, 9, 'sp4_h_r_5')
// (4, 9, 'sp4_h_r_16')
// (5, 9, 'local_g2_5')
// (5, 9, 'lutff_7/in_2')
// (5, 9, 'sp4_h_r_29')
// (6, 5, 'neigh_op_tnr_4')
// (6, 6, 'neigh_op_rgt_4')
// (6, 6, 'sp4_r_v_b_40')
// (6, 7, 'neigh_op_bnr_4')
// (6, 7, 'sp4_r_v_b_29')
// (6, 8, 'sp4_r_v_b_16')
// (6, 9, 'sp4_h_r_40')
// (6, 9, 'sp4_r_v_b_5')
// (7, 5, 'neigh_op_top_4')
// (7, 5, 'sp4_v_t_40')
// (7, 6, 'lutff_4/out')
// (7, 6, 'sp4_v_b_40')
// (7, 7, 'neigh_op_bot_4')
// (7, 7, 'sp4_v_b_29')
// (7, 8, 'sp4_v_b_16')
// (7, 9, 'sp4_h_l_40')
// (7, 9, 'sp4_v_b_5')
// (8, 5, 'neigh_op_tnl_4')
// (8, 6, 'neigh_op_lft_4')
// (8, 7, 'neigh_op_bnl_4')

wire n575;
// (3, 9, 'sp4_r_v_b_38')
// (3, 10, 'sp4_r_v_b_27')
// (3, 11, 'local_g2_6')
// (3, 11, 'lutff_6/in_2')
// (3, 11, 'sp4_r_v_b_14')
// (3, 12, 'sp4_r_v_b_3')
// (4, 8, 'sp4_v_t_38')
// (4, 9, 'sp4_v_b_38')
// (4, 10, 'sp4_v_b_27')
// (4, 11, 'neigh_op_tnr_7')
// (4, 11, 'sp4_v_b_14')
// (4, 12, 'neigh_op_rgt_7')
// (4, 12, 'sp4_h_r_3')
// (4, 12, 'sp4_v_b_3')
// (4, 13, 'local_g0_7')
// (4, 13, 'lutff_5/in_2')
// (4, 13, 'neigh_op_bnr_7')
// (5, 11, 'neigh_op_top_7')
// (5, 12, 'lutff_7/out')
// (5, 12, 'sp4_h_r_14')
// (5, 13, 'neigh_op_bot_7')
// (6, 11, 'neigh_op_tnl_7')
// (6, 12, 'neigh_op_lft_7')
// (6, 12, 'sp4_h_r_27')
// (6, 13, 'neigh_op_bnl_7')
// (7, 12, 'sp4_h_r_38')
// (8, 12, 'sp4_h_l_38')

wire n576;
// (3, 10, 'local_g0_2')
// (3, 10, 'lutff_global/cen')
// (3, 10, 'sp4_h_r_10')
// (3, 10, 'sp4_h_r_6')
// (4, 10, 'local_g1_3')
// (4, 10, 'lutff_global/cen')
// (4, 10, 'sp4_h_r_19')
// (4, 10, 'sp4_h_r_23')
// (5, 10, 'sp4_h_r_30')
// (5, 10, 'sp4_h_r_34')
// (6, 9, 'neigh_op_tnr_5')
// (6, 10, 'neigh_op_rgt_5')
// (6, 10, 'sp4_h_r_43')
// (6, 10, 'sp4_h_r_47')
// (6, 11, 'neigh_op_bnr_5')
// (7, 9, 'neigh_op_top_5')
// (7, 10, 'lutff_5/out')
// (7, 10, 'sp4_h_l_43')
// (7, 10, 'sp4_h_l_47')
// (7, 10, 'sp4_h_r_10')
// (7, 11, 'neigh_op_bot_5')
// (8, 9, 'neigh_op_tnl_5')
// (8, 10, 'neigh_op_lft_5')
// (8, 10, 'sp4_h_r_23')
// (8, 11, 'neigh_op_bnl_5')
// (9, 10, 'sp4_h_r_34')
// (10, 10, 'sp4_h_r_47')
// (11, 10, 'sp4_h_l_47')

reg n577 = 0;
// (3, 10, 'neigh_op_tnr_0')
// (3, 11, 'neigh_op_rgt_0')
// (3, 12, 'neigh_op_bnr_0')
// (4, 9, 'sp4_r_v_b_41')
// (4, 10, 'neigh_op_top_0')
// (4, 10, 'sp4_r_v_b_28')
// (4, 11, 'lutff_0/out')
// (4, 11, 'sp4_h_r_0')
// (4, 11, 'sp4_r_v_b_17')
// (4, 12, 'neigh_op_bot_0')
// (4, 12, 'sp4_r_v_b_4')
// (5, 8, 'sp4_h_r_9')
// (5, 8, 'sp4_v_t_41')
// (5, 9, 'sp4_v_b_41')
// (5, 10, 'neigh_op_tnl_0')
// (5, 10, 'sp4_v_b_28')
// (5, 11, 'neigh_op_lft_0')
// (5, 11, 'sp4_h_r_13')
// (5, 11, 'sp4_v_b_17')
// (5, 12, 'neigh_op_bnl_0')
// (5, 12, 'sp4_v_b_4')
// (6, 8, 'sp4_h_r_20')
// (6, 11, 'sp4_h_r_24')
// (7, 8, 'sp4_h_r_33')
// (7, 11, 'sp4_h_r_37')
// (8, 8, 'sp4_h_r_44')
// (8, 11, 'sp4_h_l_37')
// (8, 11, 'sp4_h_r_0')
// (9, 8, 'sp4_h_l_44')
// (9, 8, 'sp4_h_r_5')
// (9, 11, 'sp4_h_r_13')
// (10, 8, 'sp4_h_r_16')
// (10, 11, 'sp4_h_r_24')
// (11, 8, 'sp4_h_r_29')
// (11, 11, 'sp4_h_r_37')
// (12, 8, 'sp4_h_r_40')
// (12, 11, 'sp4_h_l_37')
// (12, 11, 'sp4_h_r_0')
// (13, 8, 'sp4_h_l_40')
// (13, 8, 'sp4_h_r_5')
// (13, 11, 'sp4_h_r_13')
// (14, 8, 'sp4_h_r_16')
// (14, 11, 'local_g3_0')
// (14, 11, 'lutff_6/in_1')
// (14, 11, 'sp4_h_r_24')
// (15, 8, 'sp4_h_r_29')
// (15, 11, 'sp4_h_r_37')
// (16, 8, 'sp4_h_r_40')
// (16, 11, 'sp4_h_l_37')
// (16, 11, 'sp4_h_r_3')
// (16, 11, 'sp4_h_r_8')
// (17, 8, 'sp4_h_l_40')
// (17, 8, 'sp4_h_r_5')
// (17, 11, 'local_g0_5')
// (17, 11, 'lutff_1/in_0')
// (17, 11, 'lutff_2/in_1')
// (17, 11, 'sp4_h_r_14')
// (17, 11, 'sp4_h_r_21')
// (18, 8, 'local_g1_0')
// (18, 8, 'lutff_2/in_1')
// (18, 8, 'lutff_4/in_1')
// (18, 8, 'sp4_h_r_16')
// (18, 11, 'sp4_h_r_27')
// (18, 11, 'sp4_h_r_32')
// (19, 8, 'sp4_h_r_29')
// (19, 8, 'sp4_r_v_b_44')
// (19, 9, 'sp4_r_v_b_33')
// (19, 10, 'sp4_r_v_b_20')
// (19, 11, 'sp4_h_r_38')
// (19, 11, 'sp4_h_r_45')
// (19, 11, 'sp4_r_v_b_9')
// (20, 7, 'sp4_v_t_44')
// (20, 8, 'sp4_h_r_40')
// (20, 8, 'sp4_v_b_44')
// (20, 9, 'local_g2_1')
// (20, 9, 'local_g3_1')
// (20, 9, 'lutff_0/in_2')
// (20, 9, 'lutff_5/in_0')
// (20, 9, 'sp4_v_b_33')
// (20, 10, 'local_g0_4')
// (20, 10, 'lutff_0/in_2')
// (20, 10, 'sp4_v_b_20')
// (20, 11, 'sp4_h_l_38')
// (20, 11, 'sp4_h_l_45')
// (20, 11, 'sp4_v_b_9')
// (21, 8, 'sp4_h_l_40')

wire n578;
// (3, 10, 'sp4_r_v_b_44')
// (3, 11, 'sp4_r_v_b_33')
// (3, 12, 'local_g3_4')
// (3, 12, 'lutff_1/in_0')
// (3, 12, 'sp4_r_v_b_20')
// (3, 13, 'sp4_r_v_b_9')
// (4, 9, 'sp4_v_t_44')
// (4, 10, 'sp4_v_b_44')
// (4, 11, 'sp4_v_b_33')
// (4, 12, 'neigh_op_tnr_2')
// (4, 12, 'sp4_v_b_20')
// (4, 13, 'neigh_op_rgt_2')
// (4, 13, 'sp4_h_r_9')
// (4, 13, 'sp4_v_b_9')
// (4, 14, 'neigh_op_bnr_2')
// (5, 12, 'neigh_op_top_2')
// (5, 13, 'lutff_2/out')
// (5, 13, 'sp4_h_r_20')
// (5, 14, 'local_g0_2')
// (5, 14, 'lutff_0/in_0')
// (5, 14, 'lutff_2/in_0')
// (5, 14, 'neigh_op_bot_2')
// (6, 12, 'neigh_op_tnl_2')
// (6, 13, 'neigh_op_lft_2')
// (6, 13, 'sp4_h_r_33')
// (6, 14, 'neigh_op_bnl_2')
// (7, 13, 'sp4_h_r_44')
// (8, 13, 'sp4_h_l_44')

reg n579 = 0;
// (3, 11, 'local_g2_2')
// (3, 11, 'lutff_1/in_3')
// (3, 11, 'neigh_op_tnr_2')
// (3, 12, 'neigh_op_rgt_2')
// (3, 13, 'neigh_op_bnr_2')
// (4, 11, 'neigh_op_top_2')
// (4, 12, 'local_g2_2')
// (4, 12, 'lutff_2/in_2')
// (4, 12, 'lutff_2/out')
// (4, 13, 'neigh_op_bot_2')
// (5, 11, 'neigh_op_tnl_2')
// (5, 12, 'local_g1_2')
// (5, 12, 'lutff_5/in_0')
// (5, 12, 'lutff_7/in_2')
// (5, 12, 'neigh_op_lft_2')
// (5, 13, 'local_g3_2')
// (5, 13, 'lutff_4/in_3')
// (5, 13, 'lutff_6/in_1')
// (5, 13, 'neigh_op_bnl_2')

reg n580 = 0;
// (3, 11, 'neigh_op_tnr_3')
// (3, 12, 'neigh_op_rgt_3')
// (3, 13, 'local_g1_3')
// (3, 13, 'lutff_7/in_3')
// (3, 13, 'neigh_op_bnr_3')
// (4, 11, 'neigh_op_top_3')
// (4, 12, 'local_g0_3')
// (4, 12, 'lutff_3/in_2')
// (4, 12, 'lutff_3/out')
// (4, 13, 'neigh_op_bot_3')
// (5, 11, 'neigh_op_tnl_3')
// (5, 12, 'local_g1_3')
// (5, 12, 'lutff_3/in_1')
// (5, 12, 'lutff_7/in_3')
// (5, 12, 'neigh_op_lft_3')
// (5, 13, 'local_g3_3')
// (5, 13, 'lutff_4/in_2')
// (5, 13, 'lutff_6/in_2')
// (5, 13, 'neigh_op_bnl_3')

reg n581 = 0;
// (3, 11, 'neigh_op_tnr_4')
// (3, 12, 'neigh_op_rgt_4')
// (3, 13, 'neigh_op_bnr_4')
// (4, 11, 'neigh_op_top_4')
// (4, 12, 'local_g0_4')
// (4, 12, 'lutff_4/in_2')
// (4, 12, 'lutff_4/out')
// (4, 12, 'sp4_h_r_8')
// (4, 13, 'neigh_op_bot_4')
// (5, 11, 'neigh_op_tnl_4')
// (5, 12, 'neigh_op_lft_4')
// (5, 12, 'sp4_h_r_21')
// (5, 13, 'local_g2_4')
// (5, 13, 'lutff_1/in_3')
// (5, 13, 'lutff_3/in_1')
// (5, 13, 'lutff_6/in_0')
// (5, 13, 'neigh_op_bnl_4')
// (6, 12, 'sp4_h_r_32')
// (7, 12, 'local_g3_5')
// (7, 12, 'lutff_6/in_0')
// (7, 12, 'sp4_h_r_45')
// (8, 12, 'sp4_h_l_45')

reg n582 = 0;
// (3, 11, 'neigh_op_tnr_5')
// (3, 12, 'neigh_op_rgt_5')
// (3, 13, 'neigh_op_bnr_5')
// (4, 11, 'neigh_op_top_5')
// (4, 12, 'local_g3_5')
// (4, 12, 'lutff_5/in_1')
// (4, 12, 'lutff_5/out')
// (4, 12, 'sp4_h_r_10')
// (4, 12, 'sp4_r_v_b_43')
// (4, 13, 'neigh_op_bot_5')
// (4, 13, 'sp4_r_v_b_30')
// (4, 14, 'local_g3_3')
// (4, 14, 'lutff_4/in_2')
// (4, 14, 'sp4_r_v_b_19')
// (4, 15, 'sp4_r_v_b_6')
// (5, 11, 'neigh_op_tnl_5')
// (5, 11, 'sp4_v_t_43')
// (5, 12, 'neigh_op_lft_5')
// (5, 12, 'sp4_h_r_23')
// (5, 12, 'sp4_v_b_43')
// (5, 13, 'local_g2_5')
// (5, 13, 'lutff_3/in_2')
// (5, 13, 'neigh_op_bnl_5')
// (5, 13, 'sp4_v_b_30')
// (5, 14, 'sp4_v_b_19')
// (5, 15, 'sp4_v_b_6')
// (6, 12, 'sp4_h_r_34')
// (7, 12, 'local_g2_7')
// (7, 12, 'lutff_6/in_3')
// (7, 12, 'sp4_h_r_47')
// (8, 12, 'sp4_h_l_47')

reg n583 = 0;
// (3, 11, 'sp4_h_r_0')
// (4, 10, 'neigh_op_tnr_4')
// (4, 11, 'neigh_op_rgt_4')
// (4, 11, 'sp4_h_r_13')
// (4, 12, 'neigh_op_bnr_4')
// (5, 10, 'neigh_op_top_4')
// (5, 11, 'local_g2_4')
// (5, 11, 'lutff_4/in_2')
// (5, 11, 'lutff_4/out')
// (5, 11, 'sp4_h_r_24')
// (5, 12, 'neigh_op_bot_4')
// (6, 10, 'neigh_op_tnl_4')
// (6, 11, 'neigh_op_lft_4')
// (6, 11, 'sp4_h_r_37')
// (6, 12, 'neigh_op_bnl_4')
// (6, 12, 'sp4_r_v_b_40')
// (6, 13, 'sp4_r_v_b_29')
// (6, 14, 'sp4_r_v_b_16')
// (6, 15, 'sp4_r_v_b_5')
// (7, 11, 'sp4_h_l_37')
// (7, 11, 'sp4_v_t_40')
// (7, 12, 'local_g2_0')
// (7, 12, 'lutff_4/in_0')
// (7, 12, 'sp4_v_b_40')
// (7, 13, 'sp4_v_b_29')
// (7, 14, 'sp4_v_b_16')
// (7, 15, 'sp4_v_b_5')

wire n584;
// (3, 11, 'sp4_r_v_b_36')
// (3, 12, 'local_g2_6')
// (3, 12, 'lutff_4/in_2')
// (3, 12, 'lutff_5/in_3')
// (3, 12, 'neigh_op_tnr_6')
// (3, 12, 'sp4_r_v_b_25')
// (3, 13, 'neigh_op_rgt_6')
// (3, 13, 'sp4_r_v_b_12')
// (3, 14, 'neigh_op_bnr_6')
// (3, 14, 'sp4_r_v_b_1')
// (3, 15, 'sp4_r_v_b_41')
// (3, 16, 'sp4_r_v_b_28')
// (3, 17, 'local_g3_1')
// (3, 17, 'lutff_7/in_1')
// (3, 17, 'sp4_r_v_b_17')
// (3, 18, 'sp4_r_v_b_4')
// (4, 10, 'sp4_v_t_36')
// (4, 11, 'sp4_v_b_36')
// (4, 12, 'neigh_op_top_6')
// (4, 12, 'sp4_v_b_25')
// (4, 13, 'lutff_6/out')
// (4, 13, 'sp4_v_b_12')
// (4, 14, 'neigh_op_bot_6')
// (4, 14, 'sp4_v_b_1')
// (4, 14, 'sp4_v_t_41')
// (4, 15, 'sp4_v_b_41')
// (4, 16, 'sp4_v_b_28')
// (4, 17, 'sp4_v_b_17')
// (4, 18, 'sp4_v_b_4')
// (5, 12, 'neigh_op_tnl_6')
// (5, 13, 'neigh_op_lft_6')
// (5, 14, 'neigh_op_bnl_6')

wire n585;
// (3, 12, 'neigh_op_tnr_5')
// (3, 13, 'neigh_op_rgt_5')
// (3, 13, 'sp4_r_v_b_42')
// (3, 14, 'neigh_op_bnr_5')
// (3, 14, 'sp4_r_v_b_31')
// (3, 15, 'sp4_r_v_b_18')
// (3, 16, 'sp4_r_v_b_7')
// (4, 12, 'neigh_op_top_5')
// (4, 12, 'sp4_v_t_42')
// (4, 13, 'lutff_5/out')
// (4, 13, 'sp4_v_b_42')
// (4, 14, 'neigh_op_bot_5')
// (4, 14, 'sp4_v_b_31')
// (4, 15, 'local_g1_2')
// (4, 15, 'lutff_5/in_0')
// (4, 15, 'sp4_v_b_18')
// (4, 16, 'sp4_v_b_7')
// (5, 12, 'neigh_op_tnl_5')
// (5, 13, 'neigh_op_lft_5')
// (5, 14, 'neigh_op_bnl_5')

reg n586 = 0;
// (3, 12, 'sp4_r_v_b_45')
// (3, 13, 'sp4_r_v_b_32')
// (3, 14, 'neigh_op_tnr_4')
// (3, 14, 'sp4_r_v_b_21')
// (3, 15, 'neigh_op_rgt_4')
// (3, 15, 'sp4_r_v_b_8')
// (3, 16, 'neigh_op_bnr_4')
// (4, 11, 'sp4_h_r_8')
// (4, 11, 'sp4_v_t_45')
// (4, 12, 'sp4_v_b_45')
// (4, 13, 'sp4_v_b_32')
// (4, 14, 'neigh_op_top_4')
// (4, 14, 'sp4_v_b_21')
// (4, 15, 'lutff_4/out')
// (4, 15, 'sp4_v_b_8')
// (4, 16, 'neigh_op_bot_4')
// (5, 11, 'sp4_h_r_21')
// (5, 14, 'neigh_op_tnl_4')
// (5, 15, 'neigh_op_lft_4')
// (5, 16, 'neigh_op_bnl_4')
// (6, 11, 'sp4_h_r_32')
// (7, 11, 'sp4_h_r_45')
// (8, 11, 'local_g1_0')
// (8, 11, 'lutff_0/in_1')
// (8, 11, 'sp4_h_l_45')
// (8, 11, 'sp4_h_r_8')
// (9, 11, 'sp4_h_r_21')
// (10, 11, 'sp4_h_r_32')
// (11, 11, 'sp4_h_r_45')
// (12, 11, 'sp4_h_l_45')

reg n587 = 0;
// (3, 12, 'sp4_r_v_b_47')
// (3, 13, 'sp4_r_v_b_34')
// (3, 14, 'neigh_op_tnr_5')
// (3, 14, 'sp4_r_v_b_23')
// (3, 15, 'neigh_op_rgt_5')
// (3, 15, 'sp4_r_v_b_10')
// (3, 16, 'neigh_op_bnr_5')
// (4, 11, 'sp4_h_r_3')
// (4, 11, 'sp4_v_t_47')
// (4, 12, 'sp4_v_b_47')
// (4, 13, 'sp4_v_b_34')
// (4, 14, 'neigh_op_top_5')
// (4, 14, 'sp4_v_b_23')
// (4, 15, 'lutff_5/out')
// (4, 15, 'sp4_v_b_10')
// (4, 16, 'neigh_op_bot_5')
// (5, 11, 'sp4_h_r_14')
// (5, 14, 'neigh_op_tnl_5')
// (5, 15, 'neigh_op_lft_5')
// (5, 16, 'neigh_op_bnl_5')
// (6, 11, 'sp4_h_r_27')
// (7, 11, 'sp4_h_r_38')
// (8, 11, 'sp4_h_l_38')
// (8, 11, 'sp4_h_r_3')
// (9, 11, 'local_g1_6')
// (9, 11, 'lutff_2/in_3')
// (9, 11, 'sp4_h_r_14')
// (10, 11, 'sp4_h_r_27')
// (11, 11, 'sp4_h_r_38')
// (12, 11, 'sp4_h_l_38')

wire n588;
// (3, 13, 'local_g2_4')
// (3, 13, 'lutff_5/in_1')
// (3, 13, 'neigh_op_tnr_4')
// (3, 14, 'local_g2_4')
// (3, 14, 'lutff_2/in_2')
// (3, 14, 'neigh_op_rgt_4')
// (3, 15, 'neigh_op_bnr_4')
// (4, 13, 'local_g0_4')
// (4, 13, 'lutff_4/in_2')
// (4, 13, 'neigh_op_top_4')
// (4, 14, 'lutff_4/out')
// (4, 15, 'neigh_op_bot_4')
// (5, 13, 'neigh_op_tnl_4')
// (5, 14, 'neigh_op_lft_4')
// (5, 15, 'neigh_op_bnl_4')

wire n589;
// (3, 13, 'local_g2_6')
// (3, 13, 'lutff_0/in_2')
// (3, 13, 'sp4_r_v_b_38')
// (3, 14, 'neigh_op_tnr_7')
// (3, 14, 'sp4_r_v_b_27')
// (3, 15, 'neigh_op_rgt_7')
// (3, 15, 'sp4_r_v_b_14')
// (3, 16, 'neigh_op_bnr_7')
// (3, 16, 'sp4_r_v_b_3')
// (4, 12, 'sp4_v_t_38')
// (4, 13, 'sp4_v_b_38')
// (4, 14, 'neigh_op_top_7')
// (4, 14, 'sp4_v_b_27')
// (4, 15, 'lutff_7/out')
// (4, 15, 'sp4_v_b_14')
// (4, 16, 'neigh_op_bot_7')
// (4, 16, 'sp4_v_b_3')
// (5, 14, 'neigh_op_tnl_7')
// (5, 15, 'neigh_op_lft_7')
// (5, 16, 'neigh_op_bnl_7')

wire n590;
// (3, 13, 'lutff_5/cout')
// (3, 13, 'lutff_6/in_3')

wire n591;
// (3, 13, 'neigh_op_tnr_1')
// (3, 14, 'neigh_op_rgt_1')
// (3, 15, 'neigh_op_bnr_1')
// (4, 13, 'neigh_op_top_1')
// (4, 14, 'lutff_1/out')
// (4, 15, 'local_g1_1')
// (4, 15, 'lutff_5/in_3')
// (4, 15, 'neigh_op_bot_1')
// (5, 13, 'neigh_op_tnl_1')
// (5, 14, 'neigh_op_lft_1')
// (5, 15, 'neigh_op_bnl_1')

wire n592;
// (3, 13, 'neigh_op_tnr_2')
// (3, 14, 'neigh_op_rgt_2')
// (3, 14, 'sp4_r_v_b_36')
// (3, 15, 'neigh_op_bnr_2')
// (3, 15, 'sp4_r_v_b_25')
// (3, 16, 'local_g2_4')
// (3, 16, 'lutff_1/in_1')
// (3, 16, 'sp4_r_v_b_12')
// (3, 17, 'sp4_r_v_b_1')
// (4, 13, 'local_g0_2')
// (4, 13, 'local_g1_2')
// (4, 13, 'lutff_6/in_3')
// (4, 13, 'lutff_7/in_1')
// (4, 13, 'neigh_op_top_2')
// (4, 13, 'sp4_v_t_36')
// (4, 14, 'lutff_2/out')
// (4, 14, 'sp4_v_b_36')
// (4, 15, 'neigh_op_bot_2')
// (4, 15, 'sp4_v_b_25')
// (4, 16, 'local_g0_4')
// (4, 16, 'lutff_5/in_3')
// (4, 16, 'sp4_v_b_12')
// (4, 17, 'sp4_v_b_1')
// (5, 13, 'neigh_op_tnl_2')
// (5, 14, 'neigh_op_lft_2')
// (5, 15, 'neigh_op_bnl_2')

wire n593;
// (3, 13, 'neigh_op_tnr_3')
// (3, 14, 'neigh_op_rgt_3')
// (3, 15, 'neigh_op_bnr_3')
// (4, 13, 'neigh_op_top_3')
// (4, 14, 'lutff_3/out')
// (4, 15, 'local_g0_3')
// (4, 15, 'lutff_4/in_3')
// (4, 15, 'neigh_op_bot_3')
// (5, 13, 'neigh_op_tnl_3')
// (5, 14, 'neigh_op_lft_3')
// (5, 15, 'neigh_op_bnl_3')

reg n594 = 0;
// (3, 13, 'neigh_op_tnr_5')
// (3, 14, 'neigh_op_rgt_5')
// (3, 15, 'neigh_op_bnr_5')
// (4, 13, 'neigh_op_top_5')
// (4, 14, 'local_g0_5')
// (4, 14, 'local_g3_5')
// (4, 14, 'lutff_1/in_0')
// (4, 14, 'lutff_3/in_0')
// (4, 14, 'lutff_5/in_1')
// (4, 14, 'lutff_5/out')
// (4, 14, 'lutff_6/in_2')
// (4, 15, 'local_g0_5')
// (4, 15, 'lutff_6/in_1')
// (4, 15, 'neigh_op_bot_5')
// (5, 13, 'neigh_op_tnl_5')
// (5, 14, 'neigh_op_lft_5')
// (5, 15, 'neigh_op_bnl_5')

wire n595;
// (3, 13, 'neigh_op_tnr_6')
// (3, 14, 'neigh_op_rgt_6')
// (3, 15, 'local_g1_6')
// (3, 15, 'lutff_1/in_0')
// (3, 15, 'neigh_op_bnr_6')
// (4, 13, 'neigh_op_top_6')
// (4, 14, 'local_g2_6')
// (4, 14, 'lutff_0/in_2')
// (4, 14, 'lutff_6/out')
// (4, 15, 'neigh_op_bot_6')
// (5, 13, 'neigh_op_tnl_6')
// (5, 14, 'neigh_op_lft_6')
// (5, 15, 'neigh_op_bnl_6')

wire n596;
// (3, 13, 'neigh_op_tnr_7')
// (3, 14, 'neigh_op_rgt_7')
// (3, 15, 'neigh_op_bnr_7')
// (4, 13, 'neigh_op_top_7')
// (4, 14, 'local_g1_7')
// (4, 14, 'lutff_1/in_3')
// (4, 14, 'lutff_7/out')
// (4, 15, 'neigh_op_bot_7')
// (5, 13, 'neigh_op_tnl_7')
// (5, 14, 'neigh_op_lft_7')
// (5, 15, 'neigh_op_bnl_7')

wire n597;
// (3, 13, 'sp4_r_v_b_43')
// (3, 14, 'sp4_r_v_b_30')
// (3, 15, 'local_g3_3')
// (3, 15, 'lutff_0/in_0')
// (3, 15, 'sp4_r_v_b_19')
// (3, 16, 'neigh_op_tnr_3')
// (3, 16, 'sp4_r_v_b_6')
// (3, 17, 'neigh_op_rgt_3')
// (3, 17, 'sp4_r_v_b_38')
// (3, 18, 'neigh_op_bnr_3')
// (3, 18, 'sp4_r_v_b_27')
// (3, 19, 'sp4_r_v_b_14')
// (3, 20, 'sp4_r_v_b_3')
// (4, 12, 'sp4_v_t_43')
// (4, 13, 'sp4_v_b_43')
// (4, 14, 'local_g3_2')
// (4, 14, 'lutff_2/in_3')
// (4, 14, 'sp4_r_v_b_42')
// (4, 14, 'sp4_v_b_30')
// (4, 15, 'sp4_r_v_b_31')
// (4, 15, 'sp4_v_b_19')
// (4, 16, 'neigh_op_top_3')
// (4, 16, 'sp4_r_v_b_18')
// (4, 16, 'sp4_v_b_6')
// (4, 16, 'sp4_v_t_38')
// (4, 17, 'lutff_3/out')
// (4, 17, 'sp4_r_v_b_7')
// (4, 17, 'sp4_v_b_38')
// (4, 18, 'neigh_op_bot_3')
// (4, 18, 'sp4_v_b_27')
// (4, 19, 'sp4_v_b_14')
// (4, 20, 'sp4_v_b_3')
// (5, 13, 'sp4_v_t_42')
// (5, 14, 'sp4_v_b_42')
// (5, 15, 'local_g3_7')
// (5, 15, 'lutff_5/in_3')
// (5, 15, 'lutff_7/in_1')
// (5, 15, 'sp4_v_b_31')
// (5, 16, 'neigh_op_tnl_3')
// (5, 16, 'sp4_v_b_18')
// (5, 17, 'neigh_op_lft_3')
// (5, 17, 'sp4_v_b_7')
// (5, 18, 'neigh_op_bnl_3')

wire n598;
// (3, 13, 'sp4_r_v_b_47')
// (3, 14, 'sp4_r_v_b_34')
// (3, 15, 'local_g3_7')
// (3, 15, 'lutff_5/in_1')
// (3, 15, 'sp4_r_v_b_23')
// (3, 16, 'sp4_r_v_b_10')
// (4, 12, 'sp4_v_t_47')
// (4, 13, 'sp4_r_v_b_37')
// (4, 13, 'sp4_v_b_47')
// (4, 14, 'local_g0_0')
// (4, 14, 'lutff_2/in_2')
// (4, 14, 'sp4_r_v_b_24')
// (4, 14, 'sp4_v_b_34')
// (4, 15, 'neigh_op_tnr_0')
// (4, 15, 'sp4_r_v_b_13')
// (4, 15, 'sp4_v_b_23')
// (4, 16, 'neigh_op_rgt_0')
// (4, 16, 'sp4_h_r_5')
// (4, 16, 'sp4_r_v_b_0')
// (4, 16, 'sp4_v_b_10')
// (4, 17, 'neigh_op_bnr_0')
// (5, 12, 'sp4_v_t_37')
// (5, 13, 'sp4_v_b_37')
// (5, 14, 'sp4_v_b_24')
// (5, 15, 'neigh_op_top_0')
// (5, 15, 'sp4_v_b_13')
// (5, 16, 'local_g3_0')
// (5, 16, 'lutff_0/out')
// (5, 16, 'lutff_7/in_0')
// (5, 16, 'sp4_h_r_16')
// (5, 16, 'sp4_v_b_0')
// (5, 17, 'neigh_op_bot_0')
// (6, 15, 'neigh_op_tnl_0')
// (6, 16, 'neigh_op_lft_0')
// (6, 16, 'sp4_h_r_29')
// (6, 17, 'neigh_op_bnl_0')
// (7, 16, 'sp4_h_r_40')
// (8, 16, 'sp4_h_l_40')

wire n599;
// (3, 14, 'lutff_2/cout')
// (3, 14, 'lutff_3/in_3')

wire n600;
// (3, 14, 'neigh_op_tnr_0')
// (3, 15, 'neigh_op_rgt_0')
// (3, 16, 'neigh_op_bnr_0')
// (4, 14, 'neigh_op_top_0')
// (4, 15, 'local_g1_0')
// (4, 15, 'lutff_0/out')
// (4, 15, 'lutff_5/in_2')
// (4, 16, 'neigh_op_bot_0')
// (5, 14, 'neigh_op_tnl_0')
// (5, 15, 'neigh_op_lft_0')
// (5, 16, 'neigh_op_bnl_0')

wire n601;
// (3, 14, 'neigh_op_tnr_1')
// (3, 15, 'neigh_op_rgt_1')
// (3, 16, 'neigh_op_bnr_1')
// (4, 14, 'neigh_op_top_1')
// (4, 15, 'lutff_1/out')
// (4, 16, 'neigh_op_bot_1')
// (5, 14, 'neigh_op_tnl_1')
// (5, 15, 'local_g1_1')
// (5, 15, 'lutff_2/in_2')
// (5, 15, 'neigh_op_lft_1')
// (5, 16, 'neigh_op_bnl_1')

wire n602;
// (3, 14, 'neigh_op_tnr_2')
// (3, 15, 'local_g2_2')
// (3, 15, 'lutff_7/in_1')
// (3, 15, 'neigh_op_rgt_2')
// (3, 16, 'neigh_op_bnr_2')
// (4, 14, 'neigh_op_top_2')
// (4, 15, 'lutff_2/out')
// (4, 16, 'neigh_op_bot_2')
// (5, 14, 'neigh_op_tnl_2')
// (5, 15, 'neigh_op_lft_2')
// (5, 16, 'neigh_op_bnl_2')

wire n603;
// (3, 14, 'neigh_op_tnr_3')
// (3, 15, 'neigh_op_rgt_3')
// (3, 16, 'neigh_op_bnr_3')
// (4, 14, 'neigh_op_top_3')
// (4, 15, 'lutff_3/out')
// (4, 16, 'neigh_op_bot_3')
// (5, 14, 'neigh_op_tnl_3')
// (5, 15, 'local_g0_3')
// (5, 15, 'lutff_5/in_2')
// (5, 15, 'lutff_7/in_0')
// (5, 15, 'neigh_op_lft_3')
// (5, 16, 'neigh_op_bnl_3')

wire n604;
// (3, 14, 'sp4_h_r_4')
// (4, 13, 'neigh_op_tnr_6')
// (4, 14, 'neigh_op_rgt_6')
// (4, 14, 'sp4_h_r_17')
// (4, 15, 'neigh_op_bnr_6')
// (5, 13, 'neigh_op_top_6')
// (5, 14, 'local_g3_6')
// (5, 14, 'lutff_0/in_1')
// (5, 14, 'lutff_6/out')
// (5, 14, 'sp4_h_r_28')
// (5, 15, 'neigh_op_bot_6')
// (6, 13, 'neigh_op_tnl_6')
// (6, 14, 'neigh_op_lft_6')
// (6, 14, 'sp4_h_r_41')
// (6, 15, 'neigh_op_bnl_6')
// (7, 14, 'sp4_h_l_41')
// (7, 14, 'sp4_h_r_7')
// (8, 14, 'sp4_h_r_18')
// (9, 14, 'sp4_h_r_31')
// (10, 14, 'sp4_h_r_42')
// (11, 14, 'sp4_h_l_42')
// (11, 14, 'sp4_h_r_10')
// (12, 14, 'sp4_h_r_23')
// (13, 14, 'local_g2_2')
// (13, 14, 'lutff_global/cen')
// (13, 14, 'sp4_h_r_34')
// (14, 14, 'sp4_h_r_47')
// (15, 14, 'sp4_h_l_47')

reg n605 = 0;
// (3, 14, 'sp4_r_v_b_38')
// (3, 15, 'neigh_op_tnr_7')
// (3, 15, 'sp4_r_v_b_27')
// (3, 16, 'local_g3_7')
// (3, 16, 'lutff_7/in_1')
// (3, 16, 'neigh_op_rgt_7')
// (3, 16, 'sp4_r_v_b_14')
// (3, 17, 'neigh_op_bnr_7')
// (3, 17, 'sp4_r_v_b_3')
// (4, 13, 'sp4_v_t_38')
// (4, 14, 'sp4_v_b_38')
// (4, 15, 'neigh_op_top_7')
// (4, 15, 'sp4_v_b_27')
// (4, 16, 'local_g3_7')
// (4, 16, 'lutff_7/in_3')
// (4, 16, 'lutff_7/out')
// (4, 16, 'sp4_v_b_14')
// (4, 17, 'local_g1_7')
// (4, 17, 'lutff_6/in_2')
// (4, 17, 'neigh_op_bot_7')
// (4, 17, 'sp4_h_r_3')
// (4, 17, 'sp4_v_b_3')
// (5, 15, 'neigh_op_tnl_7')
// (5, 16, 'neigh_op_lft_7')
// (5, 17, 'neigh_op_bnl_7')
// (5, 17, 'sp4_h_r_14')
// (6, 17, 'sp4_h_r_27')
// (7, 17, 'local_g2_6')
// (7, 17, 'lutff_5/in_1')
// (7, 17, 'sp4_h_r_38')
// (8, 17, 'sp4_h_l_38')

wire n606;
// (3, 14, 'sp4_r_v_b_40')
// (3, 15, 'sp4_r_v_b_29')
// (3, 16, 'sp4_r_v_b_16')
// (3, 17, 'sp4_r_v_b_5')
// (4, 12, 'neigh_op_tnr_0')
// (4, 13, 'neigh_op_rgt_0')
// (4, 13, 'sp4_h_r_5')
// (4, 13, 'sp4_v_t_40')
// (4, 14, 'neigh_op_bnr_0')
// (4, 14, 'sp4_v_b_40')
// (4, 15, 'sp4_v_b_29')
// (4, 16, 'local_g0_0')
// (4, 16, 'lutff_0/in_2')
// (4, 16, 'lutff_3/in_1')
// (4, 16, 'sp4_v_b_16')
// (4, 17, 'sp4_v_b_5')
// (5, 12, 'neigh_op_top_0')
// (5, 13, 'lutff_0/out')
// (5, 13, 'sp4_h_r_16')
// (5, 14, 'neigh_op_bot_0')
// (6, 12, 'neigh_op_tnl_0')
// (6, 13, 'neigh_op_lft_0')
// (6, 13, 'sp4_h_r_29')
// (6, 14, 'neigh_op_bnl_0')
// (7, 13, 'sp4_h_r_40')
// (8, 13, 'sp4_h_l_40')

wire n607;
// (3, 15, 'neigh_op_tnr_2')
// (3, 16, 'local_g2_2')
// (3, 16, 'lutff_5/in_3')
// (3, 16, 'neigh_op_rgt_2')
// (3, 17, 'neigh_op_bnr_2')
// (4, 15, 'neigh_op_top_2')
// (4, 16, 'lutff_2/out')
// (4, 17, 'local_g1_2')
// (4, 17, 'lutff_3/in_2')
// (4, 17, 'neigh_op_bot_2')
// (5, 15, 'neigh_op_tnl_2')
// (5, 16, 'neigh_op_lft_2')
// (5, 17, 'neigh_op_bnl_2')

reg n608 = 0;
// (3, 15, 'neigh_op_tnr_3')
// (3, 16, 'neigh_op_rgt_3')
// (3, 17, 'neigh_op_bnr_3')
// (4, 13, 'sp4_r_v_b_42')
// (4, 14, 'sp4_r_v_b_31')
// (4, 15, 'neigh_op_top_3')
// (4, 15, 'sp4_r_v_b_18')
// (4, 16, 'local_g2_3')
// (4, 16, 'lutff_3/in_0')
// (4, 16, 'lutff_3/out')
// (4, 16, 'sp4_r_v_b_7')
// (4, 17, 'neigh_op_bot_3')
// (5, 12, 'sp4_v_t_42')
// (5, 13, 'sp4_v_b_42')
// (5, 14, 'local_g3_7')
// (5, 14, 'lutff_6/in_0')
// (5, 14, 'sp4_v_b_31')
// (5, 15, 'local_g3_3')
// (5, 15, 'lutff_1/in_3')
// (5, 15, 'neigh_op_tnl_3')
// (5, 15, 'sp4_v_b_18')
// (5, 16, 'neigh_op_lft_3')
// (5, 16, 'sp4_v_b_7')
// (5, 17, 'neigh_op_bnl_3')

wire n609;
// (3, 15, 'neigh_op_tnr_4')
// (3, 16, 'local_g3_4')
// (3, 16, 'lutff_2/in_3')
// (3, 16, 'neigh_op_rgt_4')
// (3, 17, 'neigh_op_bnr_4')
// (4, 15, 'neigh_op_top_4')
// (4, 16, 'lutff_4/out')
// (4, 17, 'neigh_op_bot_4')
// (5, 15, 'neigh_op_tnl_4')
// (5, 16, 'neigh_op_lft_4')
// (5, 17, 'neigh_op_bnl_4')

reg n610 = 0;
// (3, 15, 'sp4_h_r_0')
// (4, 14, 'neigh_op_tnr_4')
// (4, 15, 'neigh_op_rgt_4')
// (4, 15, 'sp4_h_r_13')
// (4, 16, 'neigh_op_bnr_4')
// (5, 14, 'neigh_op_top_4')
// (5, 15, 'lutff_4/out')
// (5, 15, 'sp4_h_r_24')
// (5, 16, 'neigh_op_bot_4')
// (6, 12, 'sp4_r_v_b_43')
// (6, 13, 'sp4_r_v_b_30')
// (6, 14, 'neigh_op_tnl_4')
// (6, 14, 'sp4_r_v_b_19')
// (6, 15, 'neigh_op_lft_4')
// (6, 15, 'sp4_h_r_37')
// (6, 15, 'sp4_r_v_b_6')
// (6, 16, 'neigh_op_bnl_4')
// (7, 11, 'sp4_v_t_43')
// (7, 12, 'sp4_v_b_43')
// (7, 13, 'local_g3_6')
// (7, 13, 'lutff_6/in_1')
// (7, 13, 'sp4_v_b_30')
// (7, 14, 'sp4_v_b_19')
// (7, 15, 'sp4_h_l_37')
// (7, 15, 'sp4_v_b_6')

wire n611;
// (3, 16, 'local_g0_4')
// (3, 16, 'lutff_6/in_0')
// (3, 16, 'sp4_h_r_4')
// (4, 15, 'neigh_op_tnr_6')
// (4, 16, 'neigh_op_rgt_6')
// (4, 16, 'sp4_h_r_17')
// (4, 17, 'neigh_op_bnr_6')
// (5, 15, 'neigh_op_top_6')
// (5, 16, 'local_g3_6')
// (5, 16, 'lutff_2/in_3')
// (5, 16, 'lutff_6/out')
// (5, 16, 'sp4_h_r_28')
// (5, 17, 'neigh_op_bot_6')
// (6, 15, 'neigh_op_tnl_6')
// (6, 16, 'neigh_op_lft_6')
// (6, 16, 'sp4_h_r_41')
// (6, 17, 'neigh_op_bnl_6')
// (7, 16, 'sp4_h_l_41')

wire n612;
// (3, 16, 'local_g2_1')
// (3, 16, 'lutff_3/in_2')
// (3, 16, 'lutff_7/in_2')
// (3, 16, 'neigh_op_tnr_1')
// (3, 17, 'neigh_op_rgt_1')
// (3, 18, 'neigh_op_bnr_1')
// (4, 16, 'local_g0_1')
// (4, 16, 'lutff_2/in_1')
// (4, 16, 'neigh_op_top_1')
// (4, 17, 'local_g0_1')
// (4, 17, 'lutff_0/in_1')
// (4, 17, 'lutff_1/out')
// (4, 17, 'lutff_5/in_2')
// (4, 17, 'lutff_7/in_2')
// (4, 18, 'neigh_op_bot_1')
// (5, 16, 'neigh_op_tnl_1')
// (5, 17, 'neigh_op_lft_1')
// (5, 18, 'neigh_op_bnl_1')

wire n613;
// (3, 16, 'neigh_op_tnr_2')
// (3, 17, 'neigh_op_rgt_2')
// (3, 18, 'neigh_op_bnr_2')
// (4, 16, 'neigh_op_top_2')
// (4, 17, 'lutff_2/out')
// (4, 18, 'neigh_op_bot_2')
// (5, 16, 'neigh_op_tnl_2')
// (5, 17, 'local_g1_2')
// (5, 17, 'lutff_4/in_1')
// (5, 17, 'neigh_op_lft_2')
// (5, 18, 'neigh_op_bnl_2')

reg n614 = 0;
// (3, 17, 'local_g0_1')
// (3, 17, 'lutff_1/in_2')
// (3, 17, 'lutff_4/in_1')
// (3, 17, 'sp4_h_r_9')
// (4, 17, 'sp4_h_r_20')
// (5, 17, 'sp4_h_r_33')
// (6, 14, 'sp4_r_v_b_41')
// (6, 15, 'sp4_r_v_b_28')
// (6, 16, 'neigh_op_tnr_2')
// (6, 16, 'sp4_r_v_b_17')
// (6, 17, 'neigh_op_rgt_2')
// (6, 17, 'sp4_h_r_44')
// (6, 17, 'sp4_r_v_b_4')
// (6, 18, 'neigh_op_bnr_2')
// (7, 13, 'sp4_v_t_41')
// (7, 14, 'sp4_v_b_41')
// (7, 15, 'sp4_v_b_28')
// (7, 16, 'neigh_op_top_2')
// (7, 16, 'sp4_v_b_17')
// (7, 17, 'lutff_2/out')
// (7, 17, 'sp4_h_l_44')
// (7, 17, 'sp4_v_b_4')
// (7, 18, 'neigh_op_bot_2')
// (8, 16, 'neigh_op_tnl_2')
// (8, 17, 'neigh_op_lft_2')
// (8, 18, 'neigh_op_bnl_2')

reg n615 = 0;
// (3, 17, 'local_g1_0')
// (3, 17, 'lutff_2/in_1')
// (3, 17, 'lutff_4/in_3')
// (3, 17, 'sp4_h_r_8')
// (4, 17, 'sp4_h_r_21')
// (5, 17, 'sp4_h_r_32')
// (6, 16, 'neigh_op_tnr_4')
// (6, 17, 'neigh_op_rgt_4')
// (6, 17, 'sp4_h_r_45')
// (6, 18, 'neigh_op_bnr_4')
// (7, 16, 'neigh_op_top_4')
// (7, 17, 'lutff_4/out')
// (7, 17, 'sp4_h_l_45')
// (7, 17, 'sp4_h_r_8')
// (7, 18, 'neigh_op_bot_4')
// (8, 16, 'neigh_op_tnl_4')
// (8, 17, 'neigh_op_lft_4')
// (8, 17, 'sp4_h_r_21')
// (8, 18, 'neigh_op_bnl_4')
// (9, 17, 'sp4_h_r_32')
// (10, 17, 'sp4_h_r_45')
// (11, 17, 'sp4_h_l_45')

wire n616;
// (3, 17, 'lutff_1/cout')
// (3, 17, 'lutff_2/in_3')

wire n617;
// (3, 17, 'neigh_op_tnr_2')
// (3, 18, 'neigh_op_rgt_2')
// (3, 19, 'neigh_op_bnr_2')
// (4, 17, 'neigh_op_top_2')
// (4, 18, 'lutff_2/out')
// (4, 19, 'neigh_op_bot_2')
// (5, 17, 'neigh_op_tnl_2')
// (5, 18, 'local_g1_2')
// (5, 18, 'lutff_4/in_3')
// (5, 18, 'neigh_op_lft_2')
// (5, 19, 'neigh_op_bnl_2')

wire n618;
// (3, 17, 'neigh_op_tnr_4')
// (3, 18, 'neigh_op_rgt_4')
// (3, 19, 'neigh_op_bnr_4')
// (4, 17, 'neigh_op_top_4')
// (4, 17, 'sp4_r_v_b_36')
// (4, 18, 'lutff_4/out')
// (4, 18, 'sp4_r_v_b_25')
// (4, 19, 'neigh_op_bot_4')
// (4, 19, 'sp4_r_v_b_12')
// (4, 20, 'sp4_r_v_b_1')
// (5, 16, 'sp4_v_t_36')
// (5, 17, 'neigh_op_tnl_4')
// (5, 17, 'sp4_v_b_36')
// (5, 18, 'neigh_op_lft_4')
// (5, 18, 'sp4_v_b_25')
// (5, 19, 'neigh_op_bnl_4')
// (5, 19, 'sp4_v_b_12')
// (5, 20, 'local_g0_1')
// (5, 20, 'lutff_1/in_2')
// (5, 20, 'sp4_v_b_1')

wire n619;
// (3, 17, 'neigh_op_tnr_6')
// (3, 18, 'neigh_op_rgt_6')
// (3, 19, 'neigh_op_bnr_6')
// (4, 17, 'neigh_op_top_6')
// (4, 17, 'sp4_r_v_b_40')
// (4, 18, 'lutff_6/out')
// (4, 18, 'sp4_r_v_b_29')
// (4, 19, 'neigh_op_bot_6')
// (4, 19, 'sp4_r_v_b_16')
// (4, 20, 'sp4_r_v_b_5')
// (5, 16, 'sp4_v_t_40')
// (5, 17, 'neigh_op_tnl_6')
// (5, 17, 'sp4_v_b_40')
// (5, 18, 'neigh_op_lft_6')
// (5, 18, 'sp4_v_b_29')
// (5, 19, 'neigh_op_bnl_6')
// (5, 19, 'sp4_v_b_16')
// (5, 20, 'local_g0_5')
// (5, 20, 'lutff_2/in_1')
// (5, 20, 'sp4_v_b_5')

reg n620 = 0;
// (3, 17, 'sp4_r_v_b_36')
// (3, 18, 'sp4_r_v_b_25')
// (3, 19, 'local_g2_4')
// (3, 19, 'lutff_1/in_1')
// (3, 19, 'sp4_r_v_b_12')
// (3, 20, 'sp4_r_v_b_1')
// (4, 16, 'sp4_v_t_36')
// (4, 17, 'sp4_v_b_36')
// (4, 18, 'local_g2_4')
// (4, 18, 'lutff_7/in_1')
// (4, 18, 'sp4_r_v_b_36')
// (4, 18, 'sp4_v_b_25')
// (4, 19, 'neigh_op_tnr_6')
// (4, 19, 'sp4_r_v_b_25')
// (4, 19, 'sp4_v_b_12')
// (4, 20, 'neigh_op_rgt_6')
// (4, 20, 'sp4_h_r_1')
// (4, 20, 'sp4_r_v_b_12')
// (4, 20, 'sp4_v_b_1')
// (4, 21, 'local_g0_6')
// (4, 21, 'lutff_5/in_1')
// (4, 21, 'neigh_op_bnr_6')
// (4, 21, 'sp4_r_v_b_1')
// (5, 14, 'sp4_r_v_b_38')
// (5, 15, 'sp4_r_v_b_27')
// (5, 16, 'sp4_r_v_b_14')
// (5, 17, 'sp4_r_v_b_3')
// (5, 17, 'sp4_v_t_36')
// (5, 18, 'sp4_r_v_b_37')
// (5, 18, 'sp4_v_b_36')
// (5, 19, 'neigh_op_top_6')
// (5, 19, 'sp4_r_v_b_24')
// (5, 19, 'sp4_v_b_25')
// (5, 20, 'local_g0_6')
// (5, 20, 'lutff_2/in_0')
// (5, 20, 'lutff_6/out')
// (5, 20, 'sp4_h_r_12')
// (5, 20, 'sp4_r_v_b_13')
// (5, 20, 'sp4_v_b_12')
// (5, 21, 'neigh_op_bot_6')
// (5, 21, 'sp4_r_v_b_0')
// (5, 21, 'sp4_v_b_1')
// (6, 13, 'sp4_h_r_8')
// (6, 13, 'sp4_v_t_38')
// (6, 14, 'sp4_v_b_38')
// (6, 15, 'sp4_v_b_27')
// (6, 16, 'sp4_v_b_14')
// (6, 17, 'sp4_h_r_5')
// (6, 17, 'sp4_v_b_3')
// (6, 17, 'sp4_v_t_37')
// (6, 18, 'sp4_v_b_37')
// (6, 19, 'neigh_op_tnl_6')
// (6, 19, 'sp4_v_b_24')
// (6, 20, 'neigh_op_lft_6')
// (6, 20, 'sp4_h_r_25')
// (6, 20, 'sp4_v_b_13')
// (6, 21, 'neigh_op_bnl_6')
// (6, 21, 'sp4_v_b_0')
// (7, 13, 'sp4_h_r_21')
// (7, 13, 'sp4_r_v_b_47')
// (7, 14, 'sp4_r_v_b_34')
// (7, 15, 'sp4_r_v_b_23')
// (7, 16, 'sp4_r_v_b_10')
// (7, 17, 'local_g1_0')
// (7, 17, 'lutff_3/in_2')
// (7, 17, 'sp4_h_r_16')
// (7, 17, 'sp4_r_v_b_42')
// (7, 18, 'sp4_r_v_b_31')
// (7, 19, 'sp4_r_v_b_18')
// (7, 20, 'sp4_h_r_36')
// (7, 20, 'sp4_r_v_b_7')
// (8, 12, 'sp4_v_t_47')
// (8, 13, 'sp4_h_r_32')
// (8, 13, 'sp4_v_b_47')
// (8, 14, 'local_g2_2')
// (8, 14, 'lutff_1/in_3')
// (8, 14, 'sp4_v_b_34')
// (8, 15, 'sp4_v_b_23')
// (8, 16, 'sp4_v_b_10')
// (8, 16, 'sp4_v_t_42')
// (8, 17, 'sp4_h_r_29')
// (8, 17, 'sp4_v_b_42')
// (8, 18, 'local_g3_7')
// (8, 18, 'lutff_3/in_1')
// (8, 18, 'lutff_4/in_0')
// (8, 18, 'sp4_v_b_31')
// (8, 19, 'sp4_v_b_18')
// (8, 20, 'sp4_h_l_36')
// (8, 20, 'sp4_v_b_7')
// (9, 13, 'local_g2_5')
// (9, 13, 'lutff_5/in_2')
// (9, 13, 'sp4_h_r_45')
// (9, 17, 'sp4_h_r_40')
// (10, 13, 'sp4_h_l_45')
// (10, 17, 'sp4_h_l_40')

reg n621 = 0;
// (3, 17, 'sp4_r_v_b_47')
// (3, 18, 'sp4_r_v_b_34')
// (3, 19, 'local_g3_7')
// (3, 19, 'lutff_0/in_2')
// (3, 19, 'lutff_1/in_3')
// (3, 19, 'sp4_r_v_b_23')
// (3, 20, 'sp4_r_v_b_10')
// (4, 16, 'sp4_v_t_47')
// (4, 17, 'sp4_r_v_b_37')
// (4, 17, 'sp4_v_b_47')
// (4, 18, 'local_g0_0')
// (4, 18, 'lutff_5/in_1')
// (4, 18, 'sp4_r_v_b_24')
// (4, 18, 'sp4_v_b_34')
// (4, 19, 'neigh_op_tnr_0')
// (4, 19, 'sp4_r_v_b_13')
// (4, 19, 'sp4_v_b_23')
// (4, 20, 'neigh_op_rgt_0')
// (4, 20, 'sp4_h_r_5')
// (4, 20, 'sp4_r_v_b_0')
// (4, 20, 'sp4_v_b_10')
// (4, 21, 'local_g1_0')
// (4, 21, 'lutff_4/in_1')
// (4, 21, 'neigh_op_bnr_0')
// (5, 14, 'sp4_r_v_b_42')
// (5, 15, 'sp4_r_v_b_31')
// (5, 15, 'sp4_r_v_b_40')
// (5, 16, 'sp4_r_v_b_18')
// (5, 16, 'sp4_r_v_b_29')
// (5, 16, 'sp4_v_t_37')
// (5, 17, 'sp4_r_v_b_16')
// (5, 17, 'sp4_r_v_b_7')
// (5, 17, 'sp4_v_b_37')
// (5, 18, 'sp4_r_v_b_41')
// (5, 18, 'sp4_r_v_b_5')
// (5, 18, 'sp4_v_b_24')
// (5, 19, 'neigh_op_top_0')
// (5, 19, 'sp4_r_v_b_28')
// (5, 19, 'sp4_r_v_b_44')
// (5, 19, 'sp4_v_b_13')
// (5, 20, 'local_g0_0')
// (5, 20, 'local_g3_0')
// (5, 20, 'lutff_0/out')
// (5, 20, 'lutff_1/in_1')
// (5, 20, 'lutff_7/in_2')
// (5, 20, 'sp4_h_r_16')
// (5, 20, 'sp4_r_v_b_17')
// (5, 20, 'sp4_r_v_b_33')
// (5, 20, 'sp4_v_b_0')
// (5, 21, 'neigh_op_bot_0')
// (5, 21, 'sp4_r_v_b_20')
// (5, 21, 'sp4_r_v_b_4')
// (5, 22, 'sp4_r_v_b_9')
// (6, 13, 'sp4_h_r_0')
// (6, 13, 'sp4_v_t_42')
// (6, 14, 'sp4_h_r_5')
// (6, 14, 'sp4_v_b_42')
// (6, 14, 'sp4_v_t_40')
// (6, 15, 'sp4_v_b_31')
// (6, 15, 'sp4_v_b_40')
// (6, 16, 'sp4_v_b_18')
// (6, 16, 'sp4_v_b_29')
// (6, 17, 'sp4_h_r_9')
// (6, 17, 'sp4_v_b_16')
// (6, 17, 'sp4_v_b_7')
// (6, 17, 'sp4_v_t_41')
// (6, 18, 'sp4_h_r_2')
// (6, 18, 'sp4_v_b_41')
// (6, 18, 'sp4_v_b_5')
// (6, 18, 'sp4_v_t_44')
// (6, 19, 'neigh_op_tnl_0')
// (6, 19, 'sp4_v_b_28')
// (6, 19, 'sp4_v_b_44')
// (6, 20, 'neigh_op_lft_0')
// (6, 20, 'sp4_h_r_29')
// (6, 20, 'sp4_v_b_17')
// (6, 20, 'sp4_v_b_33')
// (6, 21, 'neigh_op_bnl_0')
// (6, 21, 'sp4_v_b_20')
// (6, 21, 'sp4_v_b_4')
// (6, 22, 'sp4_v_b_9')
// (7, 13, 'local_g1_5')
// (7, 13, 'lutff_7/in_1')
// (7, 13, 'sp4_h_r_13')
// (7, 14, 'sp4_h_r_16')
// (7, 17, 'local_g0_4')
// (7, 17, 'lutff_7/in_1')
// (7, 17, 'sp4_h_r_20')
// (7, 18, 'sp4_h_r_15')
// (7, 20, 'sp4_h_r_40')
// (8, 13, 'sp4_h_r_24')
// (8, 14, 'local_g3_5')
// (8, 14, 'lutff_3/in_1')
// (8, 14, 'sp4_h_r_29')
// (8, 17, 'sp4_h_r_33')
// (8, 18, 'local_g3_2')
// (8, 18, 'lutff_7/in_0')
// (8, 18, 'sp4_h_r_26')
// (8, 20, 'sp4_h_l_40')
// (9, 13, 'sp4_h_r_37')
// (9, 14, 'sp4_h_r_40')
// (9, 17, 'sp4_h_r_44')
// (9, 18, 'sp4_h_r_39')
// (10, 13, 'sp4_h_l_37')
// (10, 14, 'sp4_h_l_40')
// (10, 17, 'sp4_h_l_44')
// (10, 18, 'sp4_h_l_39')

wire n622;
// (3, 18, 'lutff_1/cout')
// (3, 18, 'lutff_2/in_3')

wire n623;
// (3, 18, 'neigh_op_tnr_0')
// (3, 19, 'neigh_op_rgt_0')
// (3, 20, 'neigh_op_bnr_0')
// (4, 18, 'neigh_op_top_0')
// (4, 19, 'lutff_0/out')
// (4, 20, 'local_g0_0')
// (4, 20, 'lutff_6/in_2')
// (4, 20, 'neigh_op_bot_0')
// (5, 18, 'neigh_op_tnl_0')
// (5, 19, 'neigh_op_lft_0')
// (5, 20, 'neigh_op_bnl_0')

wire n624;
// (3, 18, 'neigh_op_tnr_1')
// (3, 19, 'neigh_op_rgt_1')
// (3, 20, 'neigh_op_bnr_1')
// (4, 18, 'neigh_op_top_1')
// (4, 19, 'lutff_1/out')
// (4, 20, 'local_g0_1')
// (4, 20, 'lutff_3/in_2')
// (4, 20, 'neigh_op_bot_1')
// (5, 18, 'neigh_op_tnl_1')
// (5, 19, 'neigh_op_lft_1')
// (5, 20, 'neigh_op_bnl_1')

wire n625;
// (3, 18, 'neigh_op_tnr_2')
// (3, 19, 'neigh_op_rgt_2')
// (3, 20, 'neigh_op_bnr_2')
// (4, 18, 'neigh_op_top_2')
// (4, 19, 'lutff_2/out')
// (4, 20, 'local_g0_2')
// (4, 20, 'lutff_2/in_2')
// (4, 20, 'neigh_op_bot_2')
// (5, 18, 'neigh_op_tnl_2')
// (5, 19, 'neigh_op_lft_2')
// (5, 20, 'neigh_op_bnl_2')

wire n626;
// (3, 18, 'neigh_op_tnr_4')
// (3, 19, 'neigh_op_rgt_4')
// (3, 20, 'neigh_op_bnr_4')
// (4, 18, 'neigh_op_top_4')
// (4, 19, 'lutff_4/out')
// (4, 20, 'local_g0_4')
// (4, 20, 'lutff_0/in_2')
// (4, 20, 'neigh_op_bot_4')
// (5, 18, 'neigh_op_tnl_4')
// (5, 19, 'neigh_op_lft_4')
// (5, 20, 'neigh_op_bnl_4')

wire n627;
// (3, 18, 'neigh_op_tnr_5')
// (3, 19, 'neigh_op_rgt_5')
// (3, 20, 'local_g1_5')
// (3, 20, 'lutff_2/in_0')
// (3, 20, 'lutff_3/in_1')
// (3, 20, 'lutff_6/in_2')
// (3, 20, 'neigh_op_bnr_5')
// (4, 18, 'neigh_op_top_5')
// (4, 19, 'local_g1_5')
// (4, 19, 'lutff_4/in_2')
// (4, 19, 'lutff_5/out')
// (4, 20, 'local_g1_5')
// (4, 20, 'lutff_2/in_0')
// (4, 20, 'lutff_3/in_3')
// (4, 20, 'lutff_4/in_0')
// (4, 20, 'lutff_6/in_0')
// (4, 20, 'lutff_7/in_1')
// (4, 20, 'neigh_op_bot_5')
// (5, 18, 'local_g2_5')
// (5, 18, 'lutff_1/in_2')
// (5, 18, 'lutff_3/in_2')
// (5, 18, 'lutff_4/in_1')
// (5, 18, 'neigh_op_tnl_5')
// (5, 19, 'local_g1_5')
// (5, 19, 'lutff_3/in_3')
// (5, 19, 'lutff_6/in_2')
// (5, 19, 'lutff_7/in_1')
// (5, 19, 'neigh_op_lft_5')
// (5, 20, 'local_g2_5')
// (5, 20, 'local_g3_5')
// (5, 20, 'lutff_1/in_3')
// (5, 20, 'lutff_2/in_2')
// (5, 20, 'lutff_3/in_2')
// (5, 20, 'lutff_7/in_3')
// (5, 20, 'neigh_op_bnl_5')

wire n628;
// (3, 18, 'neigh_op_tnr_6')
// (3, 19, 'neigh_op_rgt_6')
// (3, 20, 'local_g1_6')
// (3, 20, 'lutff_2/in_3')
// (3, 20, 'lutff_3/in_2')
// (3, 20, 'lutff_6/in_3')
// (3, 20, 'neigh_op_bnr_6')
// (4, 18, 'neigh_op_top_6')
// (4, 19, 'lutff_6/out')
// (4, 20, 'local_g1_6')
// (4, 20, 'lutff_4/in_3')
// (4, 20, 'lutff_7/in_2')
// (4, 20, 'neigh_op_bot_6')
// (5, 18, 'neigh_op_tnl_6')
// (5, 19, 'local_g1_6')
// (5, 19, 'lutff_6/in_3')
// (5, 19, 'lutff_7/in_2')
// (5, 19, 'neigh_op_lft_6')
// (5, 20, 'local_g2_6')
// (5, 20, 'lutff_3/in_1')
// (5, 20, 'lutff_7/in_1')
// (5, 20, 'neigh_op_bnl_6')

wire n629;
// (3, 18, 'neigh_op_tnr_7')
// (3, 18, 'sp4_r_v_b_43')
// (3, 19, 'neigh_op_rgt_7')
// (3, 19, 'sp4_r_v_b_30')
// (3, 20, 'local_g3_3')
// (3, 20, 'lutff_global/cen')
// (3, 20, 'neigh_op_bnr_7')
// (3, 20, 'sp4_r_v_b_19')
// (3, 21, 'sp4_r_v_b_6')
// (4, 17, 'sp4_r_v_b_39')
// (4, 17, 'sp4_v_t_43')
// (4, 18, 'neigh_op_top_7')
// (4, 18, 'sp4_r_v_b_26')
// (4, 18, 'sp4_v_b_43')
// (4, 19, 'lutff_7/out')
// (4, 19, 'sp4_r_v_b_15')
// (4, 19, 'sp4_v_b_30')
// (4, 20, 'local_g1_3')
// (4, 20, 'lutff_global/cen')
// (4, 20, 'neigh_op_bot_7')
// (4, 20, 'sp4_r_v_b_2')
// (4, 20, 'sp4_v_b_19')
// (4, 21, 'sp4_v_b_6')
// (5, 16, 'sp4_v_t_39')
// (5, 17, 'sp4_v_b_39')
// (5, 18, 'neigh_op_tnl_7')
// (5, 18, 'sp4_v_b_26')
// (5, 19, 'neigh_op_lft_7')
// (5, 19, 'sp4_v_b_15')
// (5, 20, 'local_g0_2')
// (5, 20, 'lutff_global/cen')
// (5, 20, 'neigh_op_bnl_7')
// (5, 20, 'sp4_v_b_2')

reg n630 = 0;
// (3, 18, 'sp4_h_r_4')
// (4, 13, 'sp4_r_v_b_41')
// (4, 14, 'sp4_r_v_b_28')
// (4, 15, 'sp4_r_v_b_17')
// (4, 16, 'sp4_r_v_b_4')
// (4, 17, 'neigh_op_tnr_6')
// (4, 17, 'sp4_r_v_b_41')
// (4, 18, 'local_g3_6')
// (4, 18, 'lutff_1/in_2')
// (4, 18, 'neigh_op_rgt_6')
// (4, 18, 'sp4_h_r_17')
// (4, 18, 'sp4_r_v_b_28')
// (4, 18, 'sp4_r_v_b_44')
// (4, 19, 'neigh_op_bnr_6')
// (4, 19, 'sp4_r_v_b_17')
// (4, 19, 'sp4_r_v_b_33')
// (4, 20, 'sp4_r_v_b_20')
// (4, 20, 'sp4_r_v_b_4')
// (4, 21, 'local_g2_1')
// (4, 21, 'lutff_1/in_2')
// (4, 21, 'sp4_r_v_b_9')
// (5, 12, 'sp4_v_t_41')
// (5, 13, 'local_g2_1')
// (5, 13, 'lutff_5/in_2')
// (5, 13, 'sp4_v_b_41')
// (5, 14, 'sp4_v_b_28')
// (5, 15, 'sp4_v_b_17')
// (5, 16, 'sp4_v_b_4')
// (5, 16, 'sp4_v_t_41')
// (5, 17, 'neigh_op_top_6')
// (5, 17, 'sp4_v_b_41')
// (5, 17, 'sp4_v_t_44')
// (5, 18, 'local_g2_6')
// (5, 18, 'lutff_3/in_3')
// (5, 18, 'lutff_6/out')
// (5, 18, 'sp4_h_r_28')
// (5, 18, 'sp4_v_b_28')
// (5, 18, 'sp4_v_b_44')
// (5, 19, 'local_g0_6')
// (5, 19, 'lutff_0/in_2')
// (5, 19, 'neigh_op_bot_6')
// (5, 19, 'sp4_v_b_17')
// (5, 19, 'sp4_v_b_33')
// (5, 20, 'sp4_v_b_20')
// (5, 20, 'sp4_v_b_4')
// (5, 21, 'sp4_v_b_9')
// (6, 15, 'sp4_r_v_b_41')
// (6, 16, 'sp4_r_v_b_28')
// (6, 17, 'neigh_op_tnl_6')
// (6, 17, 'sp4_r_v_b_17')
// (6, 18, 'neigh_op_lft_6')
// (6, 18, 'sp4_h_r_41')
// (6, 18, 'sp4_r_v_b_4')
// (6, 19, 'neigh_op_bnl_6')
// (7, 14, 'sp4_h_r_9')
// (7, 14, 'sp4_v_t_41')
// (7, 15, 'sp4_v_b_41')
// (7, 16, 'sp4_v_b_28')
// (7, 17, 'sp4_v_b_17')
// (7, 18, 'sp4_h_l_41')
// (7, 18, 'sp4_h_r_0')
// (7, 18, 'sp4_h_r_7')
// (7, 18, 'sp4_v_b_4')
// (8, 14, 'local_g1_4')
// (8, 14, 'lutff_1/in_0')
// (8, 14, 'sp4_h_r_20')
// (8, 18, 'local_g0_2')
// (8, 18, 'local_g0_5')
// (8, 18, 'lutff_2/in_3')
// (8, 18, 'lutff_7/in_1')
// (8, 18, 'sp4_h_r_13')
// (8, 18, 'sp4_h_r_18')
// (9, 14, 'sp4_h_r_33')
// (9, 18, 'sp4_h_r_24')
// (9, 18, 'sp4_h_r_31')
// (10, 14, 'sp4_h_r_44')
// (10, 18, 'sp4_h_r_37')
// (10, 18, 'sp4_h_r_42')
// (11, 14, 'sp4_h_l_44')
// (11, 18, 'sp4_h_l_37')
// (11, 18, 'sp4_h_l_42')

wire n631;
// (3, 18, 'sp4_r_v_b_36')
// (3, 18, 'sp4_r_v_b_42')
// (3, 19, 'sp4_r_v_b_25')
// (3, 19, 'sp4_r_v_b_31')
// (3, 20, 'local_g2_4')
// (3, 20, 'local_g3_2')
// (3, 20, 'lutff_0/in_3')
// (3, 20, 'lutff_5/in_3')
// (3, 20, 'sp4_r_v_b_12')
// (3, 20, 'sp4_r_v_b_18')
// (3, 21, 'sp4_r_v_b_1')
// (3, 21, 'sp4_r_v_b_7')
// (4, 12, 'sp4_r_v_b_41')
// (4, 13, 'sp4_r_v_b_28')
// (4, 14, 'sp4_r_v_b_17')
// (4, 15, 'sp4_r_v_b_4')
// (4, 16, 'sp4_r_v_b_37')
// (4, 16, 'sp4_r_v_b_42')
// (4, 17, 'sp4_h_r_1')
// (4, 17, 'sp4_r_v_b_24')
// (4, 17, 'sp4_r_v_b_31')
// (4, 17, 'sp4_v_t_36')
// (4, 17, 'sp4_v_t_42')
// (4, 18, 'sp4_r_v_b_13')
// (4, 18, 'sp4_r_v_b_18')
// (4, 18, 'sp4_v_b_36')
// (4, 18, 'sp4_v_b_42')
// (4, 19, 'sp4_r_v_b_0')
// (4, 19, 'sp4_r_v_b_7')
// (4, 19, 'sp4_v_b_25')
// (4, 19, 'sp4_v_b_31')
// (4, 20, 'local_g1_2')
// (4, 20, 'lutff_5/in_0')
// (4, 20, 'sp4_v_b_12')
// (4, 20, 'sp4_v_b_18')
// (4, 21, 'sp4_v_b_1')
// (4, 21, 'sp4_v_b_7')
// (5, 11, 'sp12_h_r_0')
// (5, 11, 'sp12_v_t_23')
// (5, 11, 'sp4_h_r_4')
// (5, 11, 'sp4_v_t_41')
// (5, 12, 'sp12_v_b_23')
// (5, 12, 'sp4_v_b_41')
// (5, 13, 'sp12_v_b_20')
// (5, 13, 'sp4_v_b_28')
// (5, 14, 'sp12_v_b_19')
// (5, 14, 'sp4_v_b_17')
// (5, 15, 'sp12_v_b_16')
// (5, 15, 'sp4_v_b_4')
// (5, 15, 'sp4_v_t_37')
// (5, 15, 'sp4_v_t_42')
// (5, 16, 'sp12_v_b_15')
// (5, 16, 'sp4_v_b_37')
// (5, 16, 'sp4_v_b_42')
// (5, 17, 'sp12_v_b_12')
// (5, 17, 'sp4_h_r_12')
// (5, 17, 'sp4_v_b_24')
// (5, 17, 'sp4_v_b_31')
// (5, 18, 'local_g0_5')
// (5, 18, 'lutff_0/in_1')
// (5, 18, 'lutff_6/in_1')
// (5, 18, 'sp12_v_b_11')
// (5, 18, 'sp4_v_b_13')
// (5, 18, 'sp4_v_b_18')
// (5, 19, 'local_g0_7')
// (5, 19, 'lutff_2/in_3')
// (5, 19, 'lutff_4/in_1')
// (5, 19, 'sp12_v_b_8')
// (5, 19, 'sp4_v_b_0')
// (5, 19, 'sp4_v_b_7')
// (5, 20, 'local_g2_7')
// (5, 20, 'lutff_4/in_3')
// (5, 20, 'lutff_5/in_0')
// (5, 20, 'sp12_v_b_7')
// (5, 21, 'sp12_v_b_4')
// (5, 22, 'sp12_v_b_3')
// (5, 23, 'sp12_v_b_0')
// (6, 10, 'neigh_op_tnr_6')
// (6, 11, 'neigh_op_rgt_6')
// (6, 11, 'sp12_h_r_3')
// (6, 11, 'sp4_h_r_17')
// (6, 12, 'neigh_op_bnr_6')
// (6, 17, 'sp4_h_r_25')
// (7, 10, 'neigh_op_top_6')
// (7, 10, 'sp4_r_v_b_40')
// (7, 11, 'lutff_6/out')
// (7, 11, 'sp12_h_r_4')
// (7, 11, 'sp4_h_r_28')
// (7, 11, 'sp4_r_v_b_29')
// (7, 12, 'neigh_op_bot_6')
// (7, 12, 'sp4_r_v_b_16')
// (7, 13, 'sp4_r_v_b_5')
// (7, 14, 'sp4_r_v_b_45')
// (7, 15, 'sp4_r_v_b_32')
// (7, 16, 'sp4_r_v_b_21')
// (7, 17, 'sp4_h_r_36')
// (7, 17, 'sp4_r_v_b_8')
// (8, 9, 'sp4_v_t_40')
// (8, 10, 'neigh_op_tnl_6')
// (8, 10, 'sp4_v_b_40')
// (8, 11, 'neigh_op_lft_6')
// (8, 11, 'sp12_h_r_7')
// (8, 11, 'sp4_h_r_41')
// (8, 11, 'sp4_v_b_29')
// (8, 12, 'neigh_op_bnl_6')
// (8, 12, 'sp4_v_b_16')
// (8, 13, 'sp4_v_b_5')
// (8, 13, 'sp4_v_t_45')
// (8, 14, 'sp4_v_b_45')
// (8, 15, 'sp4_v_b_32')
// (8, 16, 'sp4_v_b_21')
// (8, 17, 'sp4_h_l_36')
// (8, 17, 'sp4_v_b_8')
// (9, 11, 'sp12_h_r_8')
// (9, 11, 'sp4_h_l_41')
// (10, 11, 'sp12_h_r_11')
// (11, 11, 'sp12_h_r_12')
// (12, 11, 'sp12_h_r_15')
// (13, 11, 'sp12_h_r_16')
// (14, 11, 'sp12_h_r_19')
// (15, 11, 'sp12_h_r_20')
// (16, 11, 'sp12_h_r_23')
// (17, 11, 'sp12_h_l_23')

wire n632;
// (3, 19, 'lutff_1/cout')
// (3, 19, 'lutff_2/in_3')

wire n633;
// (3, 19, 'lutff_2/cout')
// (3, 19, 'lutff_3/in_3')

wire n634;
// (3, 19, 'lutff_3/cout')
// (3, 19, 'lutff_4/in_3')

wire n635;
// (3, 19, 'lutff_4/cout')
// (3, 19, 'lutff_5/in_3')

wire n636;
// (3, 19, 'neigh_op_tnr_2')
// (3, 20, 'neigh_op_rgt_2')
// (3, 21, 'neigh_op_bnr_2')
// (4, 19, 'neigh_op_top_2')
// (4, 20, 'local_g2_2')
// (4, 20, 'lutff_1/in_1')
// (4, 20, 'lutff_2/out')
// (4, 21, 'neigh_op_bot_2')
// (5, 19, 'neigh_op_tnl_2')
// (5, 20, 'neigh_op_lft_2')
// (5, 21, 'neigh_op_bnl_2')

wire n637;
// (3, 19, 'neigh_op_tnr_3')
// (3, 20, 'local_g2_3')
// (3, 20, 'lutff_5/in_0')
// (3, 20, 'neigh_op_rgt_3')
// (3, 21, 'neigh_op_bnr_3')
// (4, 19, 'neigh_op_top_3')
// (4, 20, 'lutff_3/out')
// (4, 21, 'neigh_op_bot_3')
// (5, 19, 'neigh_op_tnl_3')
// (5, 20, 'neigh_op_lft_3')
// (5, 21, 'neigh_op_bnl_3')

wire n638;
// (3, 19, 'neigh_op_tnr_4')
// (3, 20, 'neigh_op_rgt_4')
// (3, 21, 'neigh_op_bnr_4')
// (4, 19, 'neigh_op_top_4')
// (4, 20, 'local_g3_4')
// (4, 20, 'lutff_1/in_2')
// (4, 20, 'lutff_4/out')
// (4, 21, 'neigh_op_bot_4')
// (5, 19, 'neigh_op_tnl_4')
// (5, 20, 'neigh_op_lft_4')
// (5, 21, 'neigh_op_bnl_4')

wire n639;
// (3, 19, 'neigh_op_tnr_5')
// (3, 20, 'neigh_op_rgt_5')
// (3, 21, 'neigh_op_bnr_5')
// (4, 19, 'neigh_op_top_5')
// (4, 20, 'local_g3_5')
// (4, 20, 'lutff_1/in_3')
// (4, 20, 'lutff_5/out')
// (4, 21, 'neigh_op_bot_5')
// (5, 19, 'neigh_op_tnl_5')
// (5, 20, 'neigh_op_lft_5')
// (5, 21, 'neigh_op_bnl_5')

wire n640;
// (3, 19, 'neigh_op_tnr_7')
// (3, 20, 'neigh_op_rgt_7')
// (3, 21, 'neigh_op_bnr_7')
// (4, 19, 'neigh_op_top_7')
// (4, 20, 'lutff_7/out')
// (4, 21, 'neigh_op_bot_7')
// (5, 19, 'neigh_op_tnl_7')
// (5, 20, 'local_g1_7')
// (5, 20, 'lutff_6/in_2')
// (5, 20, 'neigh_op_lft_7')
// (5, 21, 'neigh_op_bnl_7')

wire n641;
// (3, 19, 'sp4_r_v_b_37')
// (3, 20, 'sp4_r_v_b_24')
// (3, 21, 'neigh_op_tnr_0')
// (3, 21, 'sp4_r_v_b_13')
// (3, 22, 'neigh_op_rgt_0')
// (3, 22, 'sp4_r_v_b_0')
// (3, 23, 'neigh_op_bnr_0')
// (4, 18, 'sp4_v_t_37')
// (4, 19, 'sp4_v_b_37')
// (4, 20, 'local_g3_0')
// (4, 20, 'lutff_4/in_1')
// (4, 20, 'sp4_v_b_24')
// (4, 21, 'neigh_op_top_0')
// (4, 21, 'sp4_v_b_13')
// (4, 22, 'lutff_0/out')
// (4, 22, 'sp4_v_b_0')
// (4, 23, 'neigh_op_bot_0')
// (5, 21, 'neigh_op_tnl_0')
// (5, 22, 'neigh_op_lft_0')
// (5, 23, 'neigh_op_bnl_0')

reg n642 = 0;
// (3, 19, 'sp4_r_v_b_46')
// (3, 20, 'sp4_r_v_b_35')
// (3, 21, 'sp4_r_v_b_22')
// (3, 22, 'sp4_r_v_b_11')
// (4, 17, 'neigh_op_tnr_0')
// (4, 18, 'local_g2_0')
// (4, 18, 'lutff_0/in_2')
// (4, 18, 'neigh_op_rgt_0')
// (4, 18, 'sp4_h_r_5')
// (4, 18, 'sp4_v_t_46')
// (4, 19, 'neigh_op_bnr_0')
// (4, 19, 'sp4_v_b_46')
// (4, 20, 'sp4_v_b_35')
// (4, 21, 'local_g1_6')
// (4, 21, 'lutff_0/in_1')
// (4, 21, 'sp4_v_b_22')
// (4, 22, 'sp4_v_b_11')
// (5, 15, 'sp4_r_v_b_36')
// (5, 16, 'sp4_r_v_b_25')
// (5, 17, 'neigh_op_top_0')
// (5, 17, 'sp4_r_v_b_12')
// (5, 18, 'local_g1_0')
// (5, 18, 'lutff_0/out')
// (5, 18, 'lutff_1/in_0')
// (5, 18, 'lutff_3/in_0')
// (5, 18, 'sp4_h_r_0')
// (5, 18, 'sp4_h_r_16')
// (5, 18, 'sp4_r_v_b_1')
// (5, 19, 'local_g0_0')
// (5, 19, 'lutff_0/in_0')
// (5, 19, 'neigh_op_bot_0')
// (6, 14, 'sp4_h_r_1')
// (6, 14, 'sp4_v_t_36')
// (6, 15, 'sp4_v_b_36')
// (6, 16, 'sp4_v_b_25')
// (6, 17, 'neigh_op_tnl_0')
// (6, 17, 'sp4_v_b_12')
// (6, 18, 'neigh_op_lft_0')
// (6, 18, 'sp4_h_r_13')
// (6, 18, 'sp4_h_r_29')
// (6, 18, 'sp4_v_b_1')
// (6, 19, 'neigh_op_bnl_0')
// (7, 14, 'sp4_h_r_12')
// (7, 18, 'sp4_h_r_24')
// (7, 18, 'sp4_h_r_40')
// (8, 14, 'sp4_h_r_25')
// (8, 15, 'sp4_r_v_b_37')
// (8, 16, 'sp4_r_v_b_24')
// (8, 17, 'sp4_r_v_b_13')
// (8, 18, 'local_g2_5')
// (8, 18, 'lutff_6/in_1')
// (8, 18, 'lutff_7/in_2')
// (8, 18, 'sp4_h_l_40')
// (8, 18, 'sp4_h_r_37')
// (8, 18, 'sp4_r_v_b_0')
// (9, 11, 'sp4_r_v_b_42')
// (9, 12, 'sp4_r_v_b_31')
// (9, 13, 'local_g3_2')
// (9, 13, 'lutff_6/in_3')
// (9, 13, 'sp4_r_v_b_18')
// (9, 14, 'sp4_h_r_36')
// (9, 14, 'sp4_r_v_b_7')
// (9, 14, 'sp4_v_t_37')
// (9, 15, 'local_g3_5')
// (9, 15, 'lutff_7/in_3')
// (9, 15, 'sp4_v_b_37')
// (9, 16, 'sp4_v_b_24')
// (9, 17, 'sp4_v_b_13')
// (9, 18, 'sp4_h_l_37')
// (9, 18, 'sp4_v_b_0')
// (10, 10, 'sp4_v_t_42')
// (10, 11, 'sp4_v_b_42')
// (10, 12, 'sp4_v_b_31')
// (10, 13, 'sp4_v_b_18')
// (10, 14, 'sp4_h_l_36')
// (10, 14, 'sp4_v_b_7')

wire n643;
// (3, 20, 'local_g3_6')
// (3, 20, 'lutff_2/in_1')
// (3, 20, 'neigh_op_tnr_6')
// (3, 21, 'neigh_op_rgt_6')
// (3, 22, 'neigh_op_bnr_6')
// (4, 20, 'neigh_op_top_6')
// (4, 21, 'lutff_6/out')
// (4, 22, 'neigh_op_bot_6')
// (5, 20, 'neigh_op_tnl_6')
// (5, 21, 'neigh_op_lft_6')
// (5, 22, 'neigh_op_bnl_6')

wire n644;
// (3, 20, 'local_g3_7')
// (3, 20, 'lutff_3/in_3')
// (3, 20, 'neigh_op_tnr_7')
// (3, 21, 'neigh_op_rgt_7')
// (3, 22, 'neigh_op_bnr_7')
// (4, 20, 'neigh_op_top_7')
// (4, 21, 'lutff_7/out')
// (4, 22, 'neigh_op_bot_7')
// (5, 20, 'neigh_op_tnl_7')
// (5, 21, 'neigh_op_lft_7')
// (5, 22, 'neigh_op_bnl_7')

wire n645;
// (3, 20, 'neigh_op_tnr_2')
// (3, 21, 'neigh_op_rgt_2')
// (3, 22, 'neigh_op_bnr_2')
// (4, 20, 'neigh_op_top_2')
// (4, 21, 'lutff_2/out')
// (4, 22, 'neigh_op_bot_2')
// (5, 20, 'local_g2_2')
// (5, 20, 'lutff_3/in_3')
// (5, 20, 'neigh_op_tnl_2')
// (5, 21, 'neigh_op_lft_2')
// (5, 22, 'neigh_op_bnl_2')

wire n646;
// (3, 20, 'neigh_op_tnr_3')
// (3, 21, 'neigh_op_rgt_3')
// (3, 22, 'neigh_op_bnr_3')
// (4, 20, 'neigh_op_top_3')
// (4, 21, 'lutff_3/out')
// (4, 22, 'neigh_op_bot_3')
// (5, 20, 'local_g2_3')
// (5, 20, 'lutff_7/in_0')
// (5, 20, 'neigh_op_tnl_3')
// (5, 21, 'neigh_op_lft_3')
// (5, 22, 'neigh_op_bnl_3')

wire n647;
// (3, 20, 'neigh_op_tnr_5')
// (3, 21, 'neigh_op_rgt_5')
// (3, 22, 'neigh_op_bnr_5')
// (4, 20, 'local_g0_5')
// (4, 20, 'lutff_7/in_0')
// (4, 20, 'neigh_op_top_5')
// (4, 21, 'lutff_5/out')
// (4, 22, 'neigh_op_bot_5')
// (5, 20, 'neigh_op_tnl_5')
// (5, 21, 'neigh_op_lft_5')
// (5, 22, 'neigh_op_bnl_5')

wire n648;
// (3, 20, 'sp4_r_v_b_40')
// (3, 21, 'sp4_r_v_b_29')
// (3, 22, 'sp4_r_v_b_16')
// (3, 23, 'sp4_r_v_b_5')
// (4, 16, 'sp4_r_v_b_46')
// (4, 17, 'sp4_r_v_b_35')
// (4, 18, 'sp4_r_v_b_22')
// (4, 19, 'local_g1_3')
// (4, 19, 'lutff_4/in_0')
// (4, 19, 'sp4_h_r_11')
// (4, 19, 'sp4_r_v_b_11')
// (4, 19, 'sp4_v_t_40')
// (4, 20, 'local_g0_7')
// (4, 20, 'local_g2_0')
// (4, 20, 'lutff_2/in_3')
// (4, 20, 'lutff_3/in_1')
// (4, 20, 'lutff_6/in_1')
// (4, 20, 'sp4_h_r_7')
// (4, 20, 'sp4_v_b_40')
// (4, 21, 'sp4_v_b_29')
// (4, 22, 'sp4_v_b_16')
// (4, 23, 'sp4_v_b_5')
// (5, 15, 'sp4_v_t_46')
// (5, 16, 'sp4_v_b_46')
// (5, 17, 'sp4_v_b_35')
// (5, 18, 'local_g0_6')
// (5, 18, 'lutff_1/in_3')
// (5, 18, 'lutff_3/in_1')
// (5, 18, 'lutff_4/in_2')
// (5, 18, 'sp4_v_b_22')
// (5, 19, 'sp4_h_r_22')
// (5, 19, 'sp4_h_r_6')
// (5, 19, 'sp4_v_b_11')
// (5, 20, 'local_g1_2')
// (5, 20, 'lutff_1/in_0')
// (5, 20, 'lutff_2/in_3')
// (5, 20, 'sp4_h_r_18')
// (6, 18, 'neigh_op_tnr_7')
// (6, 19, 'neigh_op_rgt_7')
// (6, 19, 'sp4_h_r_19')
// (6, 19, 'sp4_h_r_3')
// (6, 19, 'sp4_h_r_35')
// (6, 20, 'neigh_op_bnr_7')
// (6, 20, 'sp4_h_r_31')
// (7, 17, 'sp4_r_v_b_39')
// (7, 18, 'neigh_op_top_7')
// (7, 18, 'sp4_r_v_b_26')
// (7, 19, 'lutff_7/out')
// (7, 19, 'sp4_h_r_14')
// (7, 19, 'sp4_h_r_30')
// (7, 19, 'sp4_h_r_46')
// (7, 19, 'sp4_r_v_b_15')
// (7, 20, 'neigh_op_bot_7')
// (7, 20, 'sp4_h_r_42')
// (7, 20, 'sp4_r_v_b_2')
// (8, 16, 'sp4_v_t_39')
// (8, 17, 'sp4_v_b_39')
// (8, 18, 'local_g2_7')
// (8, 18, 'lutff_4/in_1')
// (8, 18, 'neigh_op_tnl_7')
// (8, 18, 'sp4_v_b_26')
// (8, 19, 'neigh_op_lft_7')
// (8, 19, 'sp4_h_l_46')
// (8, 19, 'sp4_h_r_27')
// (8, 19, 'sp4_h_r_43')
// (8, 19, 'sp4_v_b_15')
// (8, 20, 'neigh_op_bnl_7')
// (8, 20, 'sp4_h_l_42')
// (8, 20, 'sp4_v_b_2')
// (9, 19, 'sp4_h_l_43')
// (9, 19, 'sp4_h_r_38')
// (10, 19, 'local_g1_6')
// (10, 19, 'lutff_7/in_2')
// (10, 19, 'sp4_h_l_38')
// (10, 19, 'sp4_h_r_6')
// (11, 19, 'sp4_h_r_19')
// (12, 19, 'sp4_h_r_30')
// (13, 19, 'sp4_h_r_43')
// (14, 19, 'sp4_h_l_43')

wire n649;
// (4, 0, 'logic_op_tnr_0')
// (4, 1, 'local_g2_0')
// (4, 1, 'lutff_7/in_1')
// (4, 1, 'neigh_op_rgt_0')
// (4, 2, 'neigh_op_bnr_0')
// (5, 0, 'logic_op_top_0')
// (5, 1, 'lutff_0/out')
// (5, 2, 'neigh_op_bot_0')
// (6, 0, 'logic_op_tnl_0')
// (6, 1, 'neigh_op_lft_0')
// (6, 2, 'neigh_op_bnl_0')

reg n650 = 0;
// (4, 0, 'logic_op_tnr_1')
// (4, 1, 'neigh_op_rgt_1')
// (4, 2, 'neigh_op_bnr_1')
// (5, 0, 'logic_op_top_1')
// (5, 1, 'local_g0_1')
// (5, 1, 'lutff_0/in_1')
// (5, 1, 'lutff_1/out')
// (5, 2, 'neigh_op_bot_1')
// (6, 0, 'logic_op_tnl_1')
// (6, 1, 'neigh_op_lft_1')
// (6, 2, 'neigh_op_bnl_1')

wire n651;
// (4, 0, 'logic_op_tnr_2')
// (4, 1, 'local_g3_2')
// (4, 1, 'lutff_1/in_2')
// (4, 1, 'neigh_op_rgt_2')
// (4, 2, 'neigh_op_bnr_2')
// (5, 0, 'logic_op_top_2')
// (5, 1, 'local_g2_2')
// (5, 1, 'lutff_2/out')
// (5, 1, 'lutff_5/in_1')
// (5, 2, 'neigh_op_bot_2')
// (6, 0, 'logic_op_tnl_2')
// (6, 1, 'neigh_op_lft_2')
// (6, 2, 'neigh_op_bnl_2')

wire n652;
// (4, 0, 'logic_op_tnr_3')
// (4, 1, 'neigh_op_rgt_3')
// (4, 1, 'sp4_r_v_b_38')
// (4, 2, 'neigh_op_bnr_3')
// (4, 2, 'sp4_r_v_b_27')
// (4, 3, 'sp4_r_v_b_14')
// (4, 4, 'sp4_r_v_b_3')
// (5, 0, 'logic_op_top_3')
// (5, 0, 'span4_vert_38')
// (5, 1, 'lutff_3/out')
// (5, 1, 'sp4_v_b_38')
// (5, 2, 'neigh_op_bot_3')
// (5, 2, 'sp4_v_b_27')
// (5, 3, 'sp4_v_b_14')
// (5, 4, 'sp4_h_r_3')
// (5, 4, 'sp4_v_b_3')
// (6, 0, 'logic_op_tnl_3')
// (6, 1, 'neigh_op_lft_3')
// (6, 2, 'neigh_op_bnl_3')
// (6, 4, 'sp4_h_r_14')
// (7, 4, 'local_g2_3')
// (7, 4, 'lutff_3/in_2')
// (7, 4, 'sp4_h_r_27')
// (8, 4, 'sp4_h_r_38')
// (9, 4, 'sp4_h_l_38')

reg n653 = 0;
// (4, 0, 'logic_op_tnr_4')
// (4, 1, 'neigh_op_rgt_4')
// (4, 2, 'neigh_op_bnr_4')
// (5, 0, 'logic_op_top_4')
// (5, 1, 'local_g2_4')
// (5, 1, 'lutff_0/in_0')
// (5, 1, 'lutff_4/out')
// (5, 2, 'neigh_op_bot_4')
// (6, 0, 'logic_op_tnl_4')
// (6, 1, 'neigh_op_lft_4')
// (6, 2, 'neigh_op_bnl_4')

wire n654;
// (4, 0, 'logic_op_tnr_5')
// (4, 1, 'neigh_op_rgt_5')
// (4, 2, 'neigh_op_bnr_5')
// (5, 0, 'logic_op_top_5')
// (5, 1, 'lutff_5/out')
// (5, 2, 'local_g1_5')
// (5, 2, 'lutff_7/in_3')
// (5, 2, 'neigh_op_bot_5')
// (6, 0, 'logic_op_tnl_5')
// (6, 1, 'neigh_op_lft_5')
// (6, 2, 'neigh_op_bnl_5')

wire n655;
// (4, 0, 'logic_op_tnr_7')
// (4, 1, 'local_g2_7')
// (4, 1, 'lutff_7/in_0')
// (4, 1, 'neigh_op_rgt_7')
// (4, 2, 'neigh_op_bnr_7')
// (5, 0, 'logic_op_top_7')
// (5, 1, 'lutff_7/out')
// (5, 2, 'neigh_op_bot_7')
// (6, 0, 'logic_op_tnl_7')
// (6, 1, 'neigh_op_lft_7')
// (6, 2, 'neigh_op_bnl_7')

wire n656;
// (4, 1, 'local_g1_3')
// (4, 1, 'lutff_global/cen')
// (4, 1, 'sp4_h_r_11')
// (5, 1, 'local_g0_2')
// (5, 1, 'lutff_global/cen')
// (5, 1, 'sp4_h_r_10')
// (5, 1, 'sp4_h_r_22')
// (6, 1, 'sp4_h_r_23')
// (6, 1, 'sp4_h_r_35')
// (7, 1, 'sp4_h_r_34')
// (7, 1, 'sp4_h_r_46')
// (7, 2, 'sp4_r_v_b_46')
// (7, 3, 'neigh_op_tnr_3')
// (7, 3, 'sp4_r_v_b_35')
// (7, 4, 'neigh_op_rgt_3')
// (7, 4, 'sp4_r_v_b_22')
// (7, 5, 'neigh_op_bnr_3')
// (7, 5, 'sp4_r_v_b_11')
// (8, 1, 'local_g1_3')
// (8, 1, 'lutff_global/cen')
// (8, 1, 'sp4_h_l_46')
// (8, 1, 'sp4_h_r_11')
// (8, 1, 'sp4_h_r_47')
// (8, 1, 'sp4_v_t_46')
// (8, 2, 'sp4_r_v_b_47')
// (8, 2, 'sp4_v_b_46')
// (8, 3, 'neigh_op_top_3')
// (8, 3, 'sp4_r_v_b_34')
// (8, 3, 'sp4_v_b_35')
// (8, 4, 'lutff_3/out')
// (8, 4, 'sp4_r_v_b_23')
// (8, 4, 'sp4_v_b_22')
// (8, 5, 'neigh_op_bot_3')
// (8, 5, 'sp4_r_v_b_10')
// (8, 5, 'sp4_v_b_11')
// (9, 1, 'sp4_h_l_47')
// (9, 1, 'sp4_h_r_22')
// (9, 1, 'sp4_v_t_47')
// (9, 2, 'sp4_v_b_47')
// (9, 3, 'neigh_op_tnl_3')
// (9, 3, 'sp4_v_b_34')
// (9, 4, 'neigh_op_lft_3')
// (9, 4, 'sp4_v_b_23')
// (9, 5, 'neigh_op_bnl_3')
// (9, 5, 'sp4_v_b_10')
// (10, 1, 'sp4_h_r_35')
// (11, 1, 'sp4_h_r_46')
// (12, 1, 'sp4_h_l_46')

reg n657 = 0;
// (4, 1, 'local_g2_2')
// (4, 1, 'lutff_6/in_2')
// (4, 1, 'neigh_op_tnr_2')
// (4, 1, 'sp4_r_v_b_33')
// (4, 2, 'neigh_op_rgt_2')
// (4, 2, 'sp4_r_v_b_20')
// (4, 3, 'neigh_op_bnr_2')
// (4, 3, 'sp4_r_v_b_9')
// (5, 0, 'span4_vert_33')
// (5, 1, 'neigh_op_top_2')
// (5, 1, 'sp4_v_b_33')
// (5, 2, 'lutff_2/out')
// (5, 2, 'sp4_v_b_20')
// (5, 3, 'neigh_op_bot_2')
// (5, 3, 'sp4_h_r_9')
// (5, 3, 'sp4_v_b_9')
// (6, 1, 'neigh_op_tnl_2')
// (6, 2, 'neigh_op_lft_2')
// (6, 3, 'neigh_op_bnl_2')
// (6, 3, 'sp4_h_r_20')
// (7, 3, 'local_g3_1')
// (7, 3, 'lutff_7/in_3')
// (7, 3, 'sp4_h_r_33')
// (8, 3, 'sp4_h_r_44')
// (9, 3, 'sp4_h_l_44')

reg n658 = 0;
// (4, 1, 'local_g2_6')
// (4, 1, 'lutff_2/in_0')
// (4, 1, 'neigh_op_tnr_6')
// (4, 2, 'neigh_op_rgt_6')
// (4, 2, 'sp4_r_v_b_44')
// (4, 3, 'local_g0_6')
// (4, 3, 'lutff_7/in_1')
// (4, 3, 'neigh_op_bnr_6')
// (4, 3, 'sp4_r_v_b_33')
// (4, 4, 'sp4_r_v_b_20')
// (4, 5, 'sp4_r_v_b_9')
// (5, 1, 'neigh_op_top_6')
// (5, 1, 'sp4_h_r_9')
// (5, 1, 'sp4_v_t_44')
// (5, 2, 'lutff_6/out')
// (5, 2, 'sp4_v_b_44')
// (5, 3, 'neigh_op_bot_6')
// (5, 3, 'sp4_v_b_33')
// (5, 4, 'sp4_v_b_20')
// (5, 5, 'sp4_v_b_9')
// (6, 1, 'neigh_op_tnl_6')
// (6, 1, 'sp4_h_r_20')
// (6, 2, 'neigh_op_lft_6')
// (6, 3, 'neigh_op_bnl_6')
// (7, 1, 'local_g3_1')
// (7, 1, 'lutff_6/in_2')
// (7, 1, 'sp4_h_r_33')
// (8, 1, 'sp4_h_r_44')
// (9, 1, 'sp4_h_l_44')

reg n659 = 0;
// (4, 1, 'local_g3_6')
// (4, 1, 'lutff_6/in_1')
// (4, 1, 'sp4_r_v_b_22')
// (4, 2, 'sp4_r_v_b_11')
// (5, 0, 'span4_vert_22')
// (5, 1, 'sp4_v_b_22')
// (5, 2, 'sp4_h_r_6')
// (5, 2, 'sp4_v_b_11')
// (6, 1, 'neigh_op_tnr_7')
// (6, 2, 'neigh_op_rgt_7')
// (6, 2, 'sp4_h_r_19')
// (6, 3, 'neigh_op_bnr_7')
// (7, 1, 'neigh_op_top_7')
// (7, 2, 'lutff_7/out')
// (7, 2, 'sp4_h_r_30')
// (7, 3, 'neigh_op_bot_7')
// (8, 1, 'neigh_op_tnl_7')
// (8, 2, 'neigh_op_lft_7')
// (8, 2, 'sp4_h_r_43')
// (8, 3, 'local_g3_7')
// (8, 3, 'lutff_2/in_0')
// (8, 3, 'neigh_op_bnl_7')
// (9, 2, 'sp4_h_l_43')

wire n660;
// (4, 1, 'neigh_op_tnr_0')
// (4, 2, 'neigh_op_rgt_0')
// (4, 3, 'local_g0_0')
// (4, 3, 'lutff_0/in_0')
// (4, 3, 'neigh_op_bnr_0')
// (5, 1, 'neigh_op_top_0')
// (5, 2, 'lutff_0/out')
// (5, 3, 'neigh_op_bot_0')
// (6, 1, 'neigh_op_tnl_0')
// (6, 2, 'neigh_op_lft_0')
// (6, 3, 'neigh_op_bnl_0')

wire n661;
// (4, 1, 'neigh_op_tnr_5')
// (4, 2, 'local_g2_5')
// (4, 2, 'lutff_6/in_1')
// (4, 2, 'neigh_op_rgt_5')
// (4, 3, 'neigh_op_bnr_5')
// (5, 1, 'neigh_op_top_5')
// (5, 2, 'lutff_5/out')
// (5, 3, 'neigh_op_bot_5')
// (6, 1, 'neigh_op_tnl_5')
// (6, 2, 'neigh_op_lft_5')
// (6, 3, 'neigh_op_bnl_5')

wire n662;
// (4, 1, 'neigh_op_tnr_7')
// (4, 2, 'neigh_op_rgt_7')
// (4, 3, 'local_g0_7')
// (4, 3, 'lutff_4/in_1')
// (4, 3, 'neigh_op_bnr_7')
// (5, 1, 'neigh_op_top_7')
// (5, 2, 'lutff_7/out')
// (5, 3, 'neigh_op_bot_7')
// (6, 1, 'neigh_op_tnl_7')
// (6, 2, 'neigh_op_lft_7')
// (6, 3, 'neigh_op_bnl_7')

wire n663;
// (4, 1, 'sp4_h_r_6')
// (5, 1, 'sp4_h_r_19')
// (6, 1, 'sp4_h_r_30')
// (6, 2, 'sp4_r_v_b_46')
// (6, 3, 'sp4_r_v_b_35')
// (6, 4, 'sp4_r_v_b_22')
// (6, 5, 'sp4_r_v_b_11')
// (7, 1, 'local_g3_3')
// (7, 1, 'lutff_global/cen')
// (7, 1, 'sp4_h_r_43')
// (7, 1, 'sp4_v_t_46')
// (7, 2, 'sp4_r_v_b_43')
// (7, 2, 'sp4_v_b_46')
// (7, 3, 'local_g3_3')
// (7, 3, 'lutff_global/cen')
// (7, 3, 'sp4_r_v_b_30')
// (7, 3, 'sp4_v_b_35')
// (7, 4, 'neigh_op_tnr_3')
// (7, 4, 'sp4_r_v_b_19')
// (7, 4, 'sp4_v_b_22')
// (7, 5, 'neigh_op_rgt_3')
// (7, 5, 'sp4_h_r_11')
// (7, 5, 'sp4_r_v_b_6')
// (7, 5, 'sp4_v_b_11')
// (7, 6, 'neigh_op_bnr_3')
// (8, 1, 'sp4_h_l_43')
// (8, 1, 'sp4_v_t_43')
// (8, 2, 'sp4_v_b_43')
// (8, 3, 'sp4_v_b_30')
// (8, 4, 'local_g1_3')
// (8, 4, 'lutff_global/cen')
// (8, 4, 'neigh_op_top_3')
// (8, 4, 'sp4_v_b_19')
// (8, 5, 'local_g3_3')
// (8, 5, 'lutff_3/out')
// (8, 5, 'lutff_global/cen')
// (8, 5, 'sp4_h_r_22')
// (8, 5, 'sp4_v_b_6')
// (8, 6, 'neigh_op_bot_3')
// (9, 4, 'neigh_op_tnl_3')
// (9, 5, 'neigh_op_lft_3')
// (9, 5, 'sp4_h_r_35')
// (9, 6, 'neigh_op_bnl_3')
// (10, 5, 'sp4_h_r_46')
// (11, 5, 'sp4_h_l_46')

wire n664;
// (4, 2, 'local_g3_2')
// (4, 2, 'lutff_6/in_3')
// (4, 2, 'neigh_op_tnr_2')
// (4, 3, 'neigh_op_rgt_2')
// (4, 4, 'neigh_op_bnr_2')
// (5, 2, 'neigh_op_top_2')
// (5, 3, 'lutff_2/out')
// (5, 4, 'neigh_op_bot_2')
// (6, 2, 'neigh_op_tnl_2')
// (6, 3, 'neigh_op_lft_2')
// (6, 4, 'neigh_op_bnl_2')

reg n665 = 0;
// (4, 2, 'neigh_op_tnr_0')
// (4, 3, 'neigh_op_rgt_0')
// (4, 4, 'neigh_op_bnr_0')
// (5, 2, 'neigh_op_top_0')
// (5, 2, 'sp4_r_v_b_44')
// (5, 3, 'local_g1_0')
// (5, 3, 'lutff_0/out')
// (5, 3, 'lutff_5/in_2')
// (5, 3, 'sp4_r_v_b_33')
// (5, 4, 'local_g1_0')
// (5, 4, 'lutff_6/in_3')
// (5, 4, 'neigh_op_bot_0')
// (5, 4, 'sp4_r_v_b_20')
// (5, 5, 'sp4_r_v_b_9')
// (6, 1, 'sp4_v_t_44')
// (6, 2, 'neigh_op_tnl_0')
// (6, 2, 'sp4_v_b_44')
// (6, 3, 'neigh_op_lft_0')
// (6, 3, 'sp4_v_b_33')
// (6, 4, 'neigh_op_bnl_0')
// (6, 4, 'sp4_v_b_20')
// (6, 5, 'sp4_h_r_3')
// (6, 5, 'sp4_v_b_9')
// (7, 5, 'local_g1_6')
// (7, 5, 'lutff_0/in_1')
// (7, 5, 'sp4_h_r_14')
// (8, 5, 'sp4_h_r_27')
// (9, 5, 'sp4_h_r_38')
// (10, 5, 'sp4_h_l_38')

reg n666 = 0;
// (4, 2, 'neigh_op_tnr_1')
// (4, 3, 'neigh_op_rgt_1')
// (4, 4, 'local_g0_1')
// (4, 4, 'lutff_3/in_0')
// (4, 4, 'neigh_op_bnr_1')
// (5, 2, 'local_g1_1')
// (5, 2, 'lutff_0/in_0')
// (5, 2, 'neigh_op_top_1')
// (5, 3, 'lutff_1/out')
// (5, 4, 'local_g1_1')
// (5, 4, 'lutff_2/in_2')
// (5, 4, 'neigh_op_bot_1')
// (6, 2, 'neigh_op_tnl_1')
// (6, 3, 'neigh_op_lft_1')
// (6, 4, 'neigh_op_bnl_1')

wire n667;
// (4, 2, 'neigh_op_tnr_4')
// (4, 3, 'local_g3_4')
// (4, 3, 'lutff_0/in_1')
// (4, 3, 'neigh_op_rgt_4')
// (4, 4, 'neigh_op_bnr_4')
// (5, 2, 'neigh_op_top_4')
// (5, 3, 'lutff_4/out')
// (5, 4, 'neigh_op_bot_4')
// (6, 2, 'neigh_op_tnl_4')
// (6, 3, 'neigh_op_lft_4')
// (6, 4, 'neigh_op_bnl_4')

wire n668;
// (4, 2, 'neigh_op_tnr_5')
// (4, 3, 'local_g3_5')
// (4, 3, 'lutff_3/in_1')
// (4, 3, 'neigh_op_rgt_5')
// (4, 4, 'neigh_op_bnr_5')
// (5, 2, 'neigh_op_top_5')
// (5, 3, 'lutff_5/out')
// (5, 4, 'neigh_op_bot_5')
// (6, 2, 'neigh_op_tnl_5')
// (6, 3, 'neigh_op_lft_5')
// (6, 4, 'neigh_op_bnl_5')

wire n669;
// (4, 2, 'neigh_op_tnr_6')
// (4, 3, 'neigh_op_rgt_6')
// (4, 4, 'neigh_op_bnr_6')
// (5, 2, 'neigh_op_top_6')
// (5, 3, 'local_g3_6')
// (5, 3, 'lutff_2/in_1')
// (5, 3, 'lutff_6/out')
// (5, 4, 'neigh_op_bot_6')
// (6, 2, 'neigh_op_tnl_6')
// (6, 3, 'neigh_op_lft_6')
// (6, 4, 'neigh_op_bnl_6')

wire n670;
// (4, 2, 'neigh_op_tnr_7')
// (4, 3, 'neigh_op_rgt_7')
// (4, 4, 'local_g1_7')
// (4, 4, 'lutff_7/in_1')
// (4, 4, 'neigh_op_bnr_7')
// (5, 2, 'neigh_op_top_7')
// (5, 3, 'lutff_7/out')
// (5, 4, 'neigh_op_bot_7')
// (6, 2, 'neigh_op_tnl_7')
// (6, 3, 'neigh_op_lft_7')
// (6, 4, 'neigh_op_bnl_7')

wire n671;
// (4, 3, 'local_g1_5')
// (4, 3, 'lutff_4/in_0')
// (4, 3, 'sp4_h_r_5')
// (5, 3, 'sp4_h_r_16')
// (6, 2, 'neigh_op_tnr_4')
// (6, 3, 'neigh_op_rgt_4')
// (6, 3, 'sp4_h_r_29')
// (6, 4, 'neigh_op_bnr_4')
// (7, 2, 'neigh_op_top_4')
// (7, 3, 'lutff_4/out')
// (7, 3, 'sp4_h_r_40')
// (7, 4, 'neigh_op_bot_4')
// (8, 2, 'neigh_op_tnl_4')
// (8, 3, 'neigh_op_lft_4')
// (8, 3, 'sp4_h_l_40')
// (8, 4, 'neigh_op_bnl_4')

wire n672;
// (4, 3, 'neigh_op_tnr_0')
// (4, 4, 'neigh_op_rgt_0')
// (4, 5, 'neigh_op_bnr_0')
// (5, 3, 'local_g0_0')
// (5, 3, 'lutff_6/in_0')
// (5, 3, 'neigh_op_top_0')
// (5, 4, 'lutff_0/out')
// (5, 5, 'neigh_op_bot_0')
// (6, 3, 'neigh_op_tnl_0')
// (6, 4, 'neigh_op_lft_0')
// (6, 5, 'neigh_op_bnl_0')

wire n673;
// (4, 3, 'neigh_op_tnr_1')
// (4, 4, 'neigh_op_rgt_1')
// (4, 5, 'local_g1_1')
// (4, 5, 'lutff_2/in_0')
// (4, 5, 'neigh_op_bnr_1')
// (5, 3, 'neigh_op_top_1')
// (5, 4, 'lutff_1/out')
// (5, 5, 'neigh_op_bot_1')
// (6, 3, 'neigh_op_tnl_1')
// (6, 4, 'neigh_op_lft_1')
// (6, 5, 'neigh_op_bnl_1')

wire n674;
// (4, 3, 'neigh_op_tnr_2')
// (4, 4, 'neigh_op_rgt_2')
// (4, 5, 'neigh_op_bnr_2')
// (5, 2, 'sp4_r_v_b_45')
// (5, 3, 'neigh_op_top_2')
// (5, 3, 'sp4_r_v_b_32')
// (5, 4, 'lutff_2/out')
// (5, 4, 'sp4_r_v_b_21')
// (5, 5, 'neigh_op_bot_2')
// (5, 5, 'sp4_r_v_b_8')
// (6, 1, 'sp4_v_t_45')
// (6, 2, 'sp4_v_b_45')
// (6, 3, 'neigh_op_tnl_2')
// (6, 3, 'sp4_v_b_32')
// (6, 4, 'neigh_op_lft_2')
// (6, 4, 'sp4_v_b_21')
// (6, 5, 'neigh_op_bnl_2')
// (6, 5, 'sp4_h_r_8')
// (6, 5, 'sp4_v_b_8')
// (7, 5, 'sp4_h_r_21')
// (8, 5, 'local_g3_0')
// (8, 5, 'lutff_4/in_1')
// (8, 5, 'sp4_h_r_32')
// (9, 5, 'sp4_h_r_45')
// (10, 5, 'sp4_h_l_45')

wire n675;
// (4, 3, 'neigh_op_tnr_4')
// (4, 4, 'local_g2_4')
// (4, 4, 'lutff_2/in_2')
// (4, 4, 'neigh_op_rgt_4')
// (4, 5, 'neigh_op_bnr_4')
// (5, 3, 'neigh_op_top_4')
// (5, 4, 'lutff_4/out')
// (5, 5, 'neigh_op_bot_4')
// (6, 3, 'neigh_op_tnl_4')
// (6, 4, 'neigh_op_lft_4')
// (6, 5, 'neigh_op_bnl_4')

wire n676;
// (4, 3, 'neigh_op_tnr_6')
// (4, 4, 'local_g3_6')
// (4, 4, 'lutff_2/in_1')
// (4, 4, 'neigh_op_rgt_6')
// (4, 5, 'neigh_op_bnr_6')
// (5, 3, 'neigh_op_top_6')
// (5, 4, 'lutff_6/out')
// (5, 5, 'neigh_op_bot_6')
// (6, 3, 'neigh_op_tnl_6')
// (6, 4, 'neigh_op_lft_6')
// (6, 5, 'neigh_op_bnl_6')

wire n677;
// (4, 3, 'neigh_op_tnr_7')
// (4, 4, 'neigh_op_rgt_7')
// (4, 5, 'local_g0_7')
// (4, 5, 'lutff_2/in_3')
// (4, 5, 'neigh_op_bnr_7')
// (5, 3, 'neigh_op_top_7')
// (5, 4, 'lutff_7/out')
// (5, 5, 'neigh_op_bot_7')
// (6, 3, 'neigh_op_tnl_7')
// (6, 4, 'neigh_op_lft_7')
// (6, 5, 'neigh_op_bnl_7')

reg n678 = 0;
// (4, 3, 'sp4_r_v_b_36')
// (4, 4, 'local_g1_1')
// (4, 4, 'lutff_1/in_3')
// (4, 4, 'lutff_3/in_1')
// (4, 4, 'neigh_op_tnr_6')
// (4, 4, 'sp4_r_v_b_25')
// (4, 5, 'neigh_op_rgt_6')
// (4, 5, 'sp4_h_r_1')
// (4, 5, 'sp4_r_v_b_12')
// (4, 6, 'neigh_op_bnr_6')
// (4, 6, 'sp4_r_v_b_1')
// (5, 2, 'sp4_v_t_36')
// (5, 3, 'sp4_v_b_36')
// (5, 4, 'neigh_op_top_6')
// (5, 4, 'sp4_v_b_25')
// (5, 5, 'lutff_6/out')
// (5, 5, 'sp4_h_r_12')
// (5, 5, 'sp4_v_b_12')
// (5, 6, 'neigh_op_bot_6')
// (5, 6, 'sp4_v_b_1')
// (6, 4, 'neigh_op_tnl_6')
// (6, 5, 'neigh_op_lft_6')
// (6, 5, 'sp4_h_r_25')
// (6, 6, 'neigh_op_bnl_6')
// (7, 5, 'local_g2_4')
// (7, 5, 'lutff_2/in_0')
// (7, 5, 'sp4_h_r_36')
// (8, 5, 'sp4_h_l_36')

wire n679;
// (4, 3, 'sp4_r_v_b_39')
// (4, 4, 'sp4_r_v_b_26')
// (4, 5, 'sp4_r_v_b_15')
// (4, 6, 'sp4_r_v_b_2')
// (4, 13, 'sp4_h_r_2')
// (5, 2, 'sp4_v_t_39')
// (5, 3, 'sp4_v_b_39')
// (5, 4, 'local_g2_2')
// (5, 4, 'lutff_2/in_0')
// (5, 4, 'sp4_v_b_26')
// (5, 5, 'sp4_v_b_15')
// (5, 6, 'sp4_h_r_9')
// (5, 6, 'sp4_v_b_2')
// (5, 13, 'local_g0_7')
// (5, 13, 'lutff_5/in_0')
// (5, 13, 'sp4_h_r_15')
// (6, 6, 'sp4_h_r_20')
// (6, 6, 'sp4_h_r_4')
// (6, 13, 'sp4_h_r_26')
// (7, 1, 'local_g2_1')
// (7, 1, 'lutff_5/in_0')
// (7, 1, 'lutff_6/in_3')
// (7, 1, 'sp4_r_v_b_33')
// (7, 2, 'local_g3_4')
// (7, 2, 'lutff_2/in_3')
// (7, 2, 'sp4_r_v_b_20')
// (7, 3, 'local_g2_1')
// (7, 3, 'lutff_7/in_2')
// (7, 3, 'sp4_r_v_b_9')
// (7, 4, 'local_g2_4')
// (7, 4, 'lutff_3/in_3')
// (7, 4, 'lutff_5/in_1')
// (7, 4, 'lutff_7/in_1')
// (7, 4, 'sp4_r_v_b_36')
// (7, 5, 'local_g3_1')
// (7, 5, 'lutff_1/in_1')
// (7, 5, 'lutff_5/in_3')
// (7, 5, 'neigh_op_tnr_6')
// (7, 5, 'sp4_r_v_b_25')
// (7, 5, 'sp4_r_v_b_41')
// (7, 6, 'neigh_op_rgt_6')
// (7, 6, 'sp4_h_r_17')
// (7, 6, 'sp4_h_r_33')
// (7, 6, 'sp4_r_v_b_12')
// (7, 6, 'sp4_r_v_b_28')
// (7, 6, 'sp4_r_v_b_44')
// (7, 7, 'neigh_op_bnr_6')
// (7, 7, 'sp4_r_v_b_1')
// (7, 7, 'sp4_r_v_b_17')
// (7, 7, 'sp4_r_v_b_33')
// (7, 8, 'sp4_r_v_b_20')
// (7, 8, 'sp4_r_v_b_4')
// (7, 9, 'sp4_r_v_b_9')
// (7, 10, 'sp4_r_v_b_37')
// (7, 10, 'sp4_r_v_b_44')
// (7, 11, 'sp4_r_v_b_24')
// (7, 11, 'sp4_r_v_b_33')
// (7, 12, 'sp4_r_v_b_13')
// (7, 12, 'sp4_r_v_b_20')
// (7, 13, 'local_g1_0')
// (7, 13, 'lutff_0/in_1')
// (7, 13, 'lutff_7/in_2')
// (7, 13, 'sp4_h_r_39')
// (7, 13, 'sp4_r_v_b_0')
// (7, 13, 'sp4_r_v_b_9')
// (8, 0, 'span12_vert_23')
// (8, 0, 'span4_vert_33')
// (8, 1, 'sp12_v_b_23')
// (8, 1, 'sp4_v_b_33')
// (8, 2, 'sp12_v_b_20')
// (8, 2, 'sp4_v_b_20')
// (8, 3, 'local_g1_6')
// (8, 3, 'lutff_2/in_3')
// (8, 3, 'lutff_4/in_1')
// (8, 3, 'sp12_v_b_19')
// (8, 3, 'sp4_h_r_6')
// (8, 3, 'sp4_v_b_9')
// (8, 3, 'sp4_v_t_36')
// (8, 4, 'sp12_v_b_16')
// (8, 4, 'sp4_v_b_36')
// (8, 4, 'sp4_v_t_41')
// (8, 5, 'neigh_op_top_6')
// (8, 5, 'sp12_v_b_15')
// (8, 5, 'sp4_v_b_25')
// (8, 5, 'sp4_v_b_41')
// (8, 5, 'sp4_v_t_44')
// (8, 6, 'lutff_6/out')
// (8, 6, 'sp12_v_b_12')
// (8, 6, 'sp4_h_r_28')
// (8, 6, 'sp4_h_r_44')
// (8, 6, 'sp4_r_v_b_45')
// (8, 6, 'sp4_v_b_12')
// (8, 6, 'sp4_v_b_28')
// (8, 6, 'sp4_v_b_44')
// (8, 7, 'neigh_op_bot_6')
// (8, 7, 'sp12_v_b_11')
// (8, 7, 'sp4_r_v_b_32')
// (8, 7, 'sp4_v_b_1')
// (8, 7, 'sp4_v_b_17')
// (8, 7, 'sp4_v_b_33')
// (8, 8, 'sp12_v_b_8')
// (8, 8, 'sp4_r_v_b_21')
// (8, 8, 'sp4_v_b_20')
// (8, 8, 'sp4_v_b_4')
// (8, 9, 'sp12_v_b_7')
// (8, 9, 'sp4_r_v_b_8')
// (8, 9, 'sp4_v_b_9')
// (8, 9, 'sp4_v_t_37')
// (8, 9, 'sp4_v_t_44')
// (8, 10, 'sp12_v_b_4')
// (8, 10, 'sp4_r_v_b_45')
// (8, 10, 'sp4_v_b_37')
// (8, 10, 'sp4_v_b_44')
// (8, 11, 'local_g2_3')
// (8, 11, 'lutff_2/in_1')
// (8, 11, 'lutff_6/in_1')
// (8, 11, 'sp12_v_b_3')
// (8, 11, 'sp4_r_v_b_32')
// (8, 11, 'sp4_v_b_24')
// (8, 11, 'sp4_v_b_33')
// (8, 12, 'sp12_v_b_0')
// (8, 12, 'sp4_r_v_b_21')
// (8, 12, 'sp4_v_b_13')
// (8, 12, 'sp4_v_b_20')
// (8, 13, 'sp4_h_l_39')
// (8, 13, 'sp4_r_v_b_8')
// (8, 13, 'sp4_v_b_0')
// (8, 13, 'sp4_v_b_9')
// (9, 3, 'sp4_h_r_19')
// (9, 5, 'local_g3_6')
// (9, 5, 'lutff_4/in_3')
// (9, 5, 'neigh_op_tnl_6')
// (9, 5, 'sp4_v_t_45')
// (9, 6, 'neigh_op_lft_6')
// (9, 6, 'sp4_h_l_44')
// (9, 6, 'sp4_h_r_41')
// (9, 6, 'sp4_v_b_45')
// (9, 7, 'local_g3_6')
// (9, 7, 'lutff_7/in_0')
// (9, 7, 'neigh_op_bnl_6')
// (9, 7, 'sp4_r_v_b_41')
// (9, 7, 'sp4_v_b_32')
// (9, 8, 'local_g0_5')
// (9, 8, 'lutff_7/in_0')
// (9, 8, 'sp4_r_v_b_28')
// (9, 8, 'sp4_v_b_21')
// (9, 9, 'local_g0_0')
// (9, 9, 'local_g1_0')
// (9, 9, 'lutff_0/in_3')
// (9, 9, 'lutff_7/in_1')
// (9, 9, 'sp4_r_v_b_17')
// (9, 9, 'sp4_v_b_8')
// (9, 9, 'sp4_v_t_45')
// (9, 10, 'sp4_r_v_b_4')
// (9, 10, 'sp4_v_b_45')
// (9, 11, 'sp4_v_b_32')
// (9, 12, 'sp4_v_b_21')
// (9, 13, 'local_g1_0')
// (9, 13, 'lutff_1/in_0')
// (9, 13, 'lutff_4/in_1')
// (9, 13, 'lutff_5/in_0')
// (9, 13, 'lutff_6/in_1')
// (9, 13, 'sp4_v_b_8')
// (10, 3, 'sp4_h_r_30')
// (10, 6, 'sp4_h_l_41')
// (10, 6, 'sp4_v_t_41')
// (10, 7, 'sp4_v_b_41')
// (10, 8, 'sp4_v_b_28')
// (10, 9, 'sp4_v_b_17')
// (10, 10, 'local_g0_4')
// (10, 10, 'lutff_4/in_0')
// (10, 10, 'sp4_v_b_4')
// (11, 3, 'sp4_h_r_43')
// (12, 3, 'sp4_h_l_43')

reg n680 = 0;
// (4, 4, 'local_g2_7')
// (4, 4, 'lutff_1/in_0')
// (4, 4, 'neigh_op_tnr_7')
// (4, 5, 'neigh_op_rgt_7')
// (4, 5, 'sp4_h_r_3')
// (4, 6, 'neigh_op_bnr_7')
// (5, 4, 'local_g1_7')
// (5, 4, 'lutff_7/in_3')
// (5, 4, 'neigh_op_top_7')
// (5, 5, 'lutff_7/out')
// (5, 5, 'sp4_h_r_14')
// (5, 6, 'neigh_op_bot_7')
// (6, 4, 'neigh_op_tnl_7')
// (6, 5, 'neigh_op_lft_7')
// (6, 5, 'sp4_h_r_27')
// (6, 6, 'neigh_op_bnl_7')
// (7, 5, 'local_g2_6')
// (7, 5, 'lutff_3/in_1')
// (7, 5, 'sp4_h_r_38')
// (8, 5, 'sp4_h_l_38')

wire n681;
// (4, 4, 'neigh_op_tnr_0')
// (4, 5, 'neigh_op_rgt_0')
// (4, 6, 'neigh_op_bnr_0')
// (5, 4, 'local_g0_0')
// (5, 4, 'lutff_0/in_2')
// (5, 4, 'neigh_op_top_0')
// (5, 5, 'lutff_0/out')
// (5, 6, 'neigh_op_bot_0')
// (6, 4, 'neigh_op_tnl_0')
// (6, 5, 'neigh_op_lft_0')
// (6, 6, 'neigh_op_bnl_0')

wire n682;
// (4, 4, 'neigh_op_tnr_1')
// (4, 5, 'local_g3_1')
// (4, 5, 'lutff_2/in_2')
// (4, 5, 'neigh_op_rgt_1')
// (4, 6, 'neigh_op_bnr_1')
// (5, 4, 'neigh_op_top_1')
// (5, 5, 'lutff_1/out')
// (5, 6, 'neigh_op_bot_1')
// (6, 4, 'neigh_op_tnl_1')
// (6, 5, 'neigh_op_lft_1')
// (6, 6, 'neigh_op_bnl_1')

reg n683 = 0;
// (4, 4, 'neigh_op_tnr_2')
// (4, 5, 'local_g2_2')
// (4, 5, 'lutff_6/in_0')
// (4, 5, 'neigh_op_rgt_2')
// (4, 6, 'neigh_op_bnr_2')
// (5, 4, 'neigh_op_top_2')
// (5, 5, 'local_g1_2')
// (5, 5, 'lutff_1/in_2')
// (5, 5, 'lutff_2/out')
// (5, 6, 'local_g0_2')
// (5, 6, 'lutff_6/in_0')
// (5, 6, 'neigh_op_bot_2')
// (6, 4, 'neigh_op_tnl_2')
// (6, 5, 'neigh_op_lft_2')
// (6, 6, 'neigh_op_bnl_2')

reg n684 = 0;
// (4, 4, 'neigh_op_tnr_3')
// (4, 5, 'local_g3_3')
// (4, 5, 'lutff_6/in_2')
// (4, 5, 'neigh_op_rgt_3')
// (4, 6, 'neigh_op_bnr_3')
// (5, 4, 'neigh_op_top_3')
// (5, 5, 'local_g3_3')
// (5, 5, 'lutff_1/in_3')
// (5, 5, 'lutff_3/out')
// (5, 5, 'sp4_h_r_6')
// (5, 6, 'neigh_op_bot_3')
// (6, 4, 'neigh_op_tnl_3')
// (6, 5, 'neigh_op_lft_3')
// (6, 5, 'sp4_h_r_19')
// (6, 6, 'neigh_op_bnl_3')
// (7, 5, 'local_g3_6')
// (7, 5, 'lutff_4/in_3')
// (7, 5, 'sp4_h_r_30')
// (8, 5, 'sp4_h_r_43')
// (9, 5, 'sp4_h_l_43')

wire n685;
// (4, 4, 'neigh_op_tnr_5')
// (4, 5, 'neigh_op_rgt_5')
// (4, 6, 'local_g0_5')
// (4, 6, 'lutff_2/in_1')
// (4, 6, 'neigh_op_bnr_5')
// (5, 4, 'neigh_op_top_5')
// (5, 5, 'lutff_5/out')
// (5, 6, 'neigh_op_bot_5')
// (6, 4, 'neigh_op_tnl_5')
// (6, 5, 'neigh_op_lft_5')
// (6, 6, 'neigh_op_bnl_5')

wire n686;
// (4, 5, 'neigh_op_tnr_1')
// (4, 6, 'local_g2_1')
// (4, 6, 'lutff_6/in_3')
// (4, 6, 'neigh_op_rgt_1')
// (4, 7, 'neigh_op_bnr_1')
// (5, 5, 'neigh_op_top_1')
// (5, 6, 'lutff_1/out')
// (5, 7, 'neigh_op_bot_1')
// (6, 5, 'neigh_op_tnl_1')
// (6, 6, 'neigh_op_lft_1')
// (6, 7, 'neigh_op_bnl_1')

wire n687;
// (4, 5, 'neigh_op_tnr_2')
// (4, 6, 'neigh_op_rgt_2')
// (4, 7, 'local_g1_2')
// (4, 7, 'lutff_5/in_0')
// (4, 7, 'neigh_op_bnr_2')
// (5, 5, 'neigh_op_top_2')
// (5, 6, 'lutff_2/out')
// (5, 7, 'neigh_op_bot_2')
// (6, 5, 'neigh_op_tnl_2')
// (6, 6, 'neigh_op_lft_2')
// (6, 7, 'neigh_op_bnl_2')

reg n688 = 0;
// (4, 5, 'neigh_op_tnr_3')
// (4, 6, 'neigh_op_rgt_3')
// (4, 6, 'sp4_r_v_b_38')
// (4, 7, 'neigh_op_bnr_3')
// (4, 7, 'sp4_r_v_b_27')
// (4, 8, 'sp4_r_v_b_14')
// (4, 9, 'sp4_r_v_b_3')
// (5, 5, 'neigh_op_top_3')
// (5, 5, 'sp4_v_t_38')
// (5, 6, 'lutff_3/out')
// (5, 6, 'sp4_v_b_38')
// (5, 7, 'neigh_op_bot_3')
// (5, 7, 'sp4_v_b_27')
// (5, 8, 'local_g1_6')
// (5, 8, 'lutff_3/in_0')
// (5, 8, 'sp4_v_b_14')
// (5, 9, 'sp4_v_b_3')
// (6, 5, 'neigh_op_tnl_3')
// (6, 6, 'neigh_op_lft_3')
// (6, 7, 'neigh_op_bnl_3')

reg n689 = 0;
// (4, 5, 'neigh_op_tnr_5')
// (4, 6, 'neigh_op_rgt_5')
// (4, 7, 'neigh_op_bnr_5')
// (5, 5, 'neigh_op_top_5')
// (5, 6, 'lutff_5/out')
// (5, 7, 'local_g0_5')
// (5, 7, 'lutff_7/in_0')
// (5, 7, 'neigh_op_bot_5')
// (6, 5, 'neigh_op_tnl_5')
// (6, 6, 'neigh_op_lft_5')
// (6, 7, 'neigh_op_bnl_5')

reg n690 = 0;
// (4, 5, 'neigh_op_tnr_6')
// (4, 6, 'neigh_op_rgt_6')
// (4, 7, 'neigh_op_bnr_6')
// (5, 5, 'neigh_op_top_6')
// (5, 6, 'lutff_6/out')
// (5, 7, 'local_g0_6')
// (5, 7, 'lutff_7/in_3')
// (5, 7, 'neigh_op_bot_6')
// (6, 5, 'neigh_op_tnl_6')
// (6, 6, 'neigh_op_lft_6')
// (6, 7, 'neigh_op_bnl_6')

wire n691;
// (4, 5, 'neigh_op_tnr_7')
// (4, 6, 'local_g2_7')
// (4, 6, 'lutff_4/in_1')
// (4, 6, 'neigh_op_rgt_7')
// (4, 7, 'neigh_op_bnr_7')
// (5, 5, 'neigh_op_top_7')
// (5, 6, 'lutff_7/out')
// (5, 7, 'neigh_op_bot_7')
// (6, 5, 'neigh_op_tnl_7')
// (6, 6, 'neigh_op_lft_7')
// (6, 7, 'neigh_op_bnl_7')

reg n692 = 0;
// (4, 6, 'local_g3_1')
// (4, 6, 'lutff_0/in_0')
// (4, 6, 'neigh_op_tnr_1')
// (4, 7, 'local_g2_1')
// (4, 7, 'lutff_7/in_2')
// (4, 7, 'neigh_op_rgt_1')
// (4, 8, 'neigh_op_bnr_1')
// (5, 6, 'neigh_op_top_1')
// (5, 7, 'lutff_1/out')
// (5, 8, 'local_g0_1')
// (5, 8, 'lutff_7/in_0')
// (5, 8, 'neigh_op_bot_1')
// (6, 6, 'neigh_op_tnl_1')
// (6, 7, 'neigh_op_lft_1')
// (6, 8, 'neigh_op_bnl_1')

reg n693 = 0;
// (4, 6, 'local_g3_4')
// (4, 6, 'lutff_0/in_3')
// (4, 6, 'lutff_6/in_1')
// (4, 6, 'neigh_op_tnr_4')
// (4, 7, 'local_g3_4')
// (4, 7, 'lutff_5/in_2')
// (4, 7, 'lutff_7/in_0')
// (4, 7, 'neigh_op_rgt_4')
// (4, 8, 'neigh_op_bnr_4')
// (5, 6, 'local_g1_4')
// (5, 6, 'lutff_2/in_1')
// (5, 6, 'neigh_op_top_4')
// (5, 7, 'lutff_4/out')
// (5, 7, 'sp4_h_r_8')
// (5, 8, 'neigh_op_bot_4')
// (6, 6, 'neigh_op_tnl_4')
// (6, 7, 'neigh_op_lft_4')
// (6, 7, 'sp4_h_r_21')
// (6, 8, 'neigh_op_bnl_4')
// (7, 7, 'local_g3_0')
// (7, 7, 'lutff_3/in_2')
// (7, 7, 'sp4_h_r_32')
// (8, 7, 'sp4_h_r_45')
// (9, 7, 'sp4_h_l_45')

wire n694;
// (4, 6, 'local_g3_5')
// (4, 6, 'lutff_4/in_0')
// (4, 6, 'neigh_op_tnr_5')
// (4, 7, 'local_g2_5')
// (4, 7, 'lutff_6/in_1')
// (4, 7, 'neigh_op_rgt_5')
// (4, 8, 'neigh_op_bnr_5')
// (5, 6, 'neigh_op_top_5')
// (5, 7, 'lutff_5/out')
// (5, 8, 'neigh_op_bot_5')
// (6, 6, 'neigh_op_tnl_5')
// (6, 7, 'neigh_op_lft_5')
// (6, 8, 'neigh_op_bnl_5')

reg n695 = 0;
// (4, 6, 'neigh_op_tnr_0')
// (4, 7, 'neigh_op_rgt_0')
// (4, 8, 'neigh_op_bnr_0')
// (5, 6, 'local_g1_0')
// (5, 6, 'lutff_5/in_0')
// (5, 6, 'neigh_op_top_0')
// (5, 7, 'local_g1_0')
// (5, 7, 'lutff_0/out')
// (5, 7, 'lutff_5/in_0')
// (5, 8, 'neigh_op_bot_0')
// (6, 6, 'neigh_op_tnl_0')
// (6, 7, 'neigh_op_lft_0')
// (6, 8, 'neigh_op_bnl_0')

wire n696;
// (4, 6, 'neigh_op_tnr_6')
// (4, 7, 'local_g3_6')
// (4, 7, 'lutff_1/in_2')
// (4, 7, 'neigh_op_rgt_6')
// (4, 8, 'neigh_op_bnr_6')
// (5, 6, 'neigh_op_top_6')
// (5, 7, 'lutff_6/out')
// (5, 8, 'neigh_op_bot_6')
// (6, 6, 'neigh_op_tnl_6')
// (6, 7, 'neigh_op_lft_6')
// (6, 8, 'neigh_op_bnl_6')

wire n697;
// (4, 6, 'neigh_op_tnr_7')
// (4, 7, 'neigh_op_rgt_7')
// (4, 8, 'neigh_op_bnr_7')
// (5, 6, 'neigh_op_top_7')
// (5, 7, 'lutff_7/out')
// (5, 7, 'sp4_r_v_b_47')
// (5, 8, 'neigh_op_bot_7')
// (5, 8, 'sp4_r_v_b_34')
// (5, 9, 'sp4_r_v_b_23')
// (5, 10, 'sp4_r_v_b_10')
// (6, 6, 'neigh_op_tnl_7')
// (6, 6, 'sp4_h_r_3')
// (6, 6, 'sp4_v_t_47')
// (6, 7, 'neigh_op_lft_7')
// (6, 7, 'sp4_v_b_47')
// (6, 8, 'neigh_op_bnl_7')
// (6, 8, 'sp4_v_b_34')
// (6, 9, 'sp4_v_b_23')
// (6, 10, 'sp4_v_b_10')
// (7, 6, 'sp4_h_r_14')
// (8, 6, 'sp4_h_r_27')
// (9, 6, 'local_g3_6')
// (9, 6, 'lutff_3/in_2')
// (9, 6, 'sp4_h_r_38')
// (10, 6, 'sp4_h_l_38')

wire n698;
// (4, 6, 'sp4_h_r_3')
// (4, 6, 'sp4_h_r_5')
// (4, 12, 'sp4_h_r_11')
// (5, 6, 'local_g0_0')
// (5, 6, 'local_g1_6')
// (5, 6, 'lutff_3/in_1')
// (5, 6, 'lutff_6/in_1')
// (5, 6, 'sp4_h_r_14')
// (5, 6, 'sp4_h_r_16')
// (5, 7, 'sp4_r_v_b_45')
// (5, 8, 'sp4_r_v_b_32')
// (5, 9, 'sp4_r_v_b_21')
// (5, 10, 'sp4_r_v_b_8')
// (5, 11, 'sp4_r_v_b_45')
// (5, 12, 'local_g1_6')
// (5, 12, 'lutff_0/in_3')
// (5, 12, 'sp4_h_r_22')
// (5, 12, 'sp4_r_v_b_32')
// (5, 13, 'sp4_r_v_b_21')
// (5, 14, 'local_g2_0')
// (5, 14, 'lutff_7/in_1')
// (5, 14, 'sp4_r_v_b_8')
// (6, 6, 'sp4_h_r_27')
// (6, 6, 'sp4_h_r_29')
// (6, 6, 'sp4_h_r_8')
// (6, 6, 'sp4_v_t_45')
// (6, 7, 'sp4_v_b_45')
// (6, 8, 'sp4_v_b_32')
// (6, 9, 'sp4_v_b_21')
// (6, 10, 'sp4_v_b_8')
// (6, 10, 'sp4_v_t_45')
// (6, 11, 'sp4_v_b_45')
// (6, 12, 'sp4_h_r_35')
// (6, 12, 'sp4_v_b_32')
// (6, 13, 'sp4_v_b_21')
// (6, 14, 'sp4_v_b_8')
// (7, 3, 'sp4_r_v_b_37')
// (7, 4, 'sp4_r_v_b_24')
// (7, 5, 'local_g2_0')
// (7, 5, 'local_g3_0')
// (7, 5, 'lutff_2/in_3')
// (7, 5, 'lutff_3/in_2')
// (7, 5, 'lutff_4/in_1')
// (7, 5, 'lutff_6/in_0')
// (7, 5, 'neigh_op_tnr_0')
// (7, 5, 'sp4_r_v_b_13')
// (7, 5, 'sp4_r_v_b_45')
// (7, 6, 'local_g3_0')
// (7, 6, 'lutff_2/in_3')
// (7, 6, 'lutff_4/in_3')
// (7, 6, 'lutff_7/in_2')
// (7, 6, 'neigh_op_rgt_0')
// (7, 6, 'sp4_h_r_21')
// (7, 6, 'sp4_h_r_38')
// (7, 6, 'sp4_h_r_40')
// (7, 6, 'sp4_r_v_b_0')
// (7, 6, 'sp4_r_v_b_32')
// (7, 7, 'neigh_op_bnr_0')
// (7, 7, 'sp4_r_v_b_21')
// (7, 7, 'sp4_r_v_b_43')
// (7, 8, 'sp4_r_v_b_30')
// (7, 8, 'sp4_r_v_b_8')
// (7, 9, 'sp4_r_v_b_19')
// (7, 9, 'sp4_r_v_b_46')
// (7, 10, 'sp4_r_v_b_35')
// (7, 10, 'sp4_r_v_b_6')
// (7, 11, 'local_g3_6')
// (7, 11, 'lutff_0/in_3')
// (7, 11, 'sp4_r_v_b_22')
// (7, 11, 'sp4_r_v_b_39')
// (7, 11, 'sp4_r_v_b_43')
// (7, 12, 'sp4_h_r_46')
// (7, 12, 'sp4_r_v_b_11')
// (7, 12, 'sp4_r_v_b_26')
// (7, 12, 'sp4_r_v_b_30')
// (7, 13, 'local_g2_7')
// (7, 13, 'local_g3_3')
// (7, 13, 'lutff_1/in_1')
// (7, 13, 'lutff_3/in_2')
// (7, 13, 'lutff_6/in_2')
// (7, 13, 'sp4_r_v_b_15')
// (7, 13, 'sp4_r_v_b_19')
// (7, 14, 'sp4_r_v_b_2')
// (7, 14, 'sp4_r_v_b_6')
// (8, 2, 'sp4_v_t_37')
// (8, 3, 'sp4_v_b_37')
// (8, 4, 'sp4_r_v_b_41')
// (8, 4, 'sp4_v_b_24')
// (8, 4, 'sp4_v_t_45')
// (8, 5, 'neigh_op_top_0')
// (8, 5, 'sp4_r_v_b_28')
// (8, 5, 'sp4_v_b_13')
// (8, 5, 'sp4_v_b_45')
// (8, 6, 'lutff_0/out')
// (8, 6, 'sp4_h_l_38')
// (8, 6, 'sp4_h_l_40')
// (8, 6, 'sp4_h_r_0')
// (8, 6, 'sp4_h_r_32')
// (8, 6, 'sp4_r_v_b_17')
// (8, 6, 'sp4_v_b_0')
// (8, 6, 'sp4_v_b_32')
// (8, 6, 'sp4_v_t_43')
// (8, 7, 'neigh_op_bot_0')
// (8, 7, 'sp4_r_v_b_4')
// (8, 7, 'sp4_v_b_21')
// (8, 7, 'sp4_v_b_43')
// (8, 8, 'sp4_r_v_b_37')
// (8, 8, 'sp4_r_v_b_42')
// (8, 8, 'sp4_v_b_30')
// (8, 8, 'sp4_v_b_8')
// (8, 8, 'sp4_v_t_46')
// (8, 9, 'sp4_r_v_b_24')
// (8, 9, 'sp4_r_v_b_31')
// (8, 9, 'sp4_v_b_19')
// (8, 9, 'sp4_v_b_46')
// (8, 10, 'local_g0_6')
// (8, 10, 'lutff_0/in_0')
// (8, 10, 'lutff_1/in_1')
// (8, 10, 'lutff_3/in_3')
// (8, 10, 'lutff_4/in_2')
// (8, 10, 'sp4_r_v_b_13')
// (8, 10, 'sp4_r_v_b_18')
// (8, 10, 'sp4_v_b_35')
// (8, 10, 'sp4_v_b_6')
// (8, 10, 'sp4_v_t_39')
// (8, 10, 'sp4_v_t_43')
// (8, 11, 'local_g0_6')
// (8, 11, 'lutff_0/in_2')
// (8, 11, 'lutff_3/in_1')
// (8, 11, 'sp4_r_v_b_0')
// (8, 11, 'sp4_r_v_b_7')
// (8, 11, 'sp4_v_b_22')
// (8, 11, 'sp4_v_b_39')
// (8, 11, 'sp4_v_b_43')
// (8, 12, 'sp4_h_l_46')
// (8, 12, 'sp4_v_b_11')
// (8, 12, 'sp4_v_b_26')
// (8, 12, 'sp4_v_b_30')
// (8, 13, 'sp4_v_b_15')
// (8, 13, 'sp4_v_b_19')
// (8, 14, 'sp4_v_b_2')
// (8, 14, 'sp4_v_b_6')
// (9, 3, 'sp4_v_t_41')
// (9, 4, 'sp4_v_b_41')
// (9, 5, 'neigh_op_tnl_0')
// (9, 5, 'sp4_v_b_28')
// (9, 6, 'neigh_op_lft_0')
// (9, 6, 'sp4_h_r_13')
// (9, 6, 'sp4_h_r_45')
// (9, 6, 'sp4_v_b_17')
// (9, 7, 'neigh_op_bnl_0')
// (9, 7, 'sp4_r_v_b_36')
// (9, 7, 'sp4_v_b_4')
// (9, 7, 'sp4_v_t_37')
// (9, 7, 'sp4_v_t_42')
// (9, 8, 'sp4_r_v_b_25')
// (9, 8, 'sp4_v_b_37')
// (9, 8, 'sp4_v_b_42')
// (9, 9, 'sp4_r_v_b_12')
// (9, 9, 'sp4_v_b_24')
// (9, 9, 'sp4_v_b_31')
// (9, 10, 'local_g0_5')
// (9, 10, 'lutff_1/in_2')
// (9, 10, 'lutff_3/in_2')
// (9, 10, 'sp4_r_v_b_1')
// (9, 10, 'sp4_v_b_13')
// (9, 10, 'sp4_v_b_18')
// (9, 11, 'local_g1_7')
// (9, 11, 'lutff_2/in_0')
// (9, 11, 'sp4_r_v_b_44')
// (9, 11, 'sp4_v_b_0')
// (9, 11, 'sp4_v_b_7')
// (9, 12, 'sp4_r_v_b_33')
// (9, 13, 'local_g3_4')
// (9, 13, 'lutff_0/in_3')
// (9, 13, 'lutff_7/in_2')
// (9, 13, 'sp4_r_v_b_20')
// (9, 14, 'sp4_r_v_b_9')
// (10, 6, 'sp4_h_l_45')
// (10, 6, 'sp4_h_r_24')
// (10, 6, 'sp4_v_t_36')
// (10, 7, 'sp4_v_b_36')
// (10, 8, 'sp4_v_b_25')
// (10, 9, 'sp4_v_b_12')
// (10, 10, 'sp4_v_b_1')
// (10, 10, 'sp4_v_t_44')
// (10, 11, 'sp4_v_b_44')
// (10, 12, 'sp4_v_b_33')
// (10, 13, 'sp4_v_b_20')
// (10, 14, 'sp4_v_b_9')
// (11, 6, 'sp4_h_r_37')
// (12, 6, 'sp4_h_l_37')

wire n699;
// (4, 6, 'sp4_h_r_4')
// (5, 6, 'local_g1_1')
// (5, 6, 'lutff_3/in_3')
// (5, 6, 'sp4_h_r_17')
// (6, 4, 'neigh_op_tnr_0')
// (6, 5, 'neigh_op_rgt_0')
// (6, 6, 'neigh_op_bnr_0')
// (6, 6, 'sp4_h_r_28')
// (7, 3, 'sp4_r_v_b_41')
// (7, 4, 'neigh_op_top_0')
// (7, 4, 'sp4_r_v_b_28')
// (7, 5, 'lutff_0/out')
// (7, 5, 'sp4_r_v_b_17')
// (7, 6, 'neigh_op_bot_0')
// (7, 6, 'sp4_h_r_41')
// (7, 6, 'sp4_r_v_b_4')
// (8, 2, 'sp4_v_t_41')
// (8, 3, 'sp4_v_b_41')
// (8, 4, 'neigh_op_tnl_0')
// (8, 4, 'sp4_v_b_28')
// (8, 5, 'neigh_op_lft_0')
// (8, 5, 'sp4_v_b_17')
// (8, 6, 'neigh_op_bnl_0')
// (8, 6, 'sp4_h_l_41')
// (8, 6, 'sp4_v_b_4')

reg n700 = 0;
// (4, 6, 'sp4_r_v_b_37')
// (4, 7, 'sp4_r_v_b_24')
// (4, 8, 'sp4_r_v_b_13')
// (4, 9, 'sp4_r_v_b_0')
// (5, 5, 'sp4_h_r_0')
// (5, 5, 'sp4_v_t_37')
// (5, 6, 'sp4_v_b_37')
// (5, 7, 'sp4_v_b_24')
// (5, 8, 'sp4_v_b_13')
// (5, 9, 'local_g0_0')
// (5, 9, 'lutff_6/in_2')
// (5, 9, 'sp4_v_b_0')
// (6, 4, 'neigh_op_tnr_4')
// (6, 5, 'neigh_op_rgt_4')
// (6, 5, 'sp4_h_r_13')
// (6, 6, 'neigh_op_bnr_4')
// (7, 4, 'neigh_op_top_4')
// (7, 5, 'lutff_4/out')
// (7, 5, 'sp4_h_r_24')
// (7, 6, 'neigh_op_bot_4')
// (8, 4, 'neigh_op_tnl_4')
// (8, 5, 'neigh_op_lft_4')
// (8, 5, 'sp4_h_r_37')
// (8, 6, 'neigh_op_bnl_4')
// (9, 5, 'sp4_h_l_37')

reg n701 = 0;
// (4, 6, 'sp4_r_v_b_47')
// (4, 7, 'sp4_r_v_b_34')
// (4, 8, 'sp4_r_v_b_23')
// (4, 9, 'sp4_r_v_b_10')
// (5, 5, 'sp4_h_r_4')
// (5, 5, 'sp4_v_t_47')
// (5, 6, 'sp4_v_b_47')
// (5, 7, 'sp4_v_b_34')
// (5, 8, 'local_g1_7')
// (5, 8, 'lutff_6/in_0')
// (5, 8, 'sp4_v_b_23')
// (5, 9, 'sp4_v_b_10')
// (6, 4, 'neigh_op_tnr_6')
// (6, 5, 'neigh_op_rgt_6')
// (6, 5, 'sp4_h_r_17')
// (6, 6, 'neigh_op_bnr_6')
// (7, 4, 'neigh_op_top_6')
// (7, 5, 'lutff_6/out')
// (7, 5, 'sp4_h_r_28')
// (7, 6, 'neigh_op_bot_6')
// (8, 4, 'neigh_op_tnl_6')
// (8, 5, 'neigh_op_lft_6')
// (8, 5, 'sp4_h_r_41')
// (8, 6, 'neigh_op_bnl_6')
// (9, 5, 'sp4_h_l_41')

reg n702 = 0;
// (4, 7, 'neigh_op_tnr_0')
// (4, 8, 'neigh_op_rgt_0')
// (4, 9, 'neigh_op_bnr_0')
// (5, 7, 'local_g0_0')
// (5, 7, 'lutff_7/in_1')
// (5, 7, 'neigh_op_top_0')
// (5, 8, 'lutff_0/out')
// (5, 9, 'neigh_op_bot_0')
// (6, 7, 'neigh_op_tnl_0')
// (6, 8, 'neigh_op_lft_0')
// (6, 9, 'neigh_op_bnl_0')

reg n703 = 0;
// (4, 7, 'neigh_op_tnr_1')
// (4, 8, 'neigh_op_rgt_1')
// (4, 9, 'neigh_op_bnr_1')
// (5, 7, 'neigh_op_top_1')
// (5, 8, 'local_g2_1')
// (5, 8, 'lutff_1/out')
// (5, 8, 'lutff_6/in_1')
// (5, 9, 'neigh_op_bot_1')
// (6, 7, 'neigh_op_tnl_1')
// (6, 8, 'neigh_op_lft_1')
// (6, 9, 'neigh_op_bnl_1')

reg n704 = 0;
// (4, 7, 'neigh_op_tnr_2')
// (4, 8, 'neigh_op_rgt_2')
// (4, 9, 'neigh_op_bnr_2')
// (5, 7, 'neigh_op_top_2')
// (5, 8, 'local_g2_2')
// (5, 8, 'lutff_2/out')
// (5, 8, 'lutff_5/in_1')
// (5, 9, 'neigh_op_bot_2')
// (6, 7, 'neigh_op_tnl_2')
// (6, 8, 'neigh_op_lft_2')
// (6, 9, 'neigh_op_bnl_2')

wire n705;
// (4, 7, 'neigh_op_tnr_3')
// (4, 8, 'neigh_op_rgt_3')
// (4, 8, 'sp4_h_r_11')
// (4, 9, 'neigh_op_bnr_3')
// (5, 7, 'neigh_op_top_3')
// (5, 8, 'lutff_3/out')
// (5, 8, 'sp4_h_r_22')
// (5, 9, 'neigh_op_bot_3')
// (6, 7, 'neigh_op_tnl_3')
// (6, 8, 'neigh_op_lft_3')
// (6, 8, 'sp4_h_r_35')
// (6, 9, 'neigh_op_bnl_3')
// (7, 8, 'sp4_h_r_46')
// (8, 8, 'sp4_h_l_46')
// (8, 8, 'sp4_h_r_7')
// (9, 8, 'sp4_h_r_18')
// (10, 8, 'local_g3_7')
// (10, 8, 'lutff_7/in_1')
// (10, 8, 'sp4_h_r_31')
// (11, 8, 'sp4_h_r_42')
// (12, 8, 'sp4_h_l_42')

reg n706 = 0;
// (4, 7, 'neigh_op_tnr_4')
// (4, 8, 'neigh_op_rgt_4')
// (4, 9, 'neigh_op_bnr_4')
// (5, 7, 'neigh_op_top_4')
// (5, 8, 'local_g3_4')
// (5, 8, 'lutff_3/in_2')
// (5, 8, 'lutff_4/out')
// (5, 9, 'neigh_op_bot_4')
// (6, 7, 'neigh_op_tnl_4')
// (6, 8, 'neigh_op_lft_4')
// (6, 9, 'neigh_op_bnl_4')

wire n707;
// (4, 7, 'neigh_op_tnr_5')
// (4, 8, 'neigh_op_rgt_5')
// (4, 9, 'neigh_op_bnr_5')
// (5, 7, 'neigh_op_top_5')
// (5, 8, 'lutff_5/out')
// (5, 8, 'sp4_h_r_10')
// (5, 9, 'neigh_op_bot_5')
// (6, 7, 'neigh_op_tnl_5')
// (6, 8, 'neigh_op_lft_5')
// (6, 8, 'sp4_h_r_23')
// (6, 9, 'neigh_op_bnl_5')
// (7, 8, 'sp4_h_r_34')
// (8, 8, 'sp4_h_r_47')
// (9, 8, 'local_g1_6')
// (9, 8, 'lutff_5/in_0')
// (9, 8, 'sp4_h_l_47')
// (9, 8, 'sp4_h_r_6')
// (10, 8, 'sp4_h_r_19')
// (11, 8, 'sp4_h_r_30')
// (12, 8, 'sp4_h_r_43')
// (13, 8, 'sp4_h_l_43')

wire n708;
// (4, 7, 'neigh_op_tnr_6')
// (4, 8, 'neigh_op_rgt_6')
// (4, 8, 'sp4_h_r_1')
// (4, 9, 'neigh_op_bnr_6')
// (5, 7, 'neigh_op_top_6')
// (5, 8, 'lutff_6/out')
// (5, 8, 'sp4_h_r_12')
// (5, 9, 'neigh_op_bot_6')
// (6, 7, 'neigh_op_tnl_6')
// (6, 8, 'neigh_op_lft_6')
// (6, 8, 'sp4_h_r_25')
// (6, 9, 'neigh_op_bnl_6')
// (7, 8, 'sp4_h_r_36')
// (8, 8, 'sp4_h_l_36')
// (8, 8, 'sp4_h_r_1')
// (9, 8, 'sp4_h_r_12')
// (10, 8, 'local_g3_1')
// (10, 8, 'lutff_1/in_1')
// (10, 8, 'sp4_h_r_25')
// (11, 8, 'sp4_h_r_36')
// (12, 8, 'sp4_h_l_36')

reg n709 = 0;
// (4, 7, 'neigh_op_tnr_7')
// (4, 8, 'neigh_op_rgt_7')
// (4, 9, 'neigh_op_bnr_7')
// (5, 7, 'neigh_op_top_7')
// (5, 8, 'local_g2_7')
// (5, 8, 'lutff_5/in_0')
// (5, 8, 'lutff_7/out')
// (5, 9, 'neigh_op_bot_7')
// (6, 7, 'neigh_op_tnl_7')
// (6, 8, 'neigh_op_lft_7')
// (6, 9, 'neigh_op_bnl_7')

reg n710 = 0;
// (4, 7, 'sp4_h_r_1')
// (5, 7, 'local_g1_4')
// (5, 7, 'lutff_7/in_2')
// (5, 7, 'sp4_h_r_12')
// (6, 5, 'neigh_op_tnr_2')
// (6, 6, 'neigh_op_rgt_2')
// (6, 7, 'neigh_op_bnr_2')
// (6, 7, 'sp4_h_r_25')
// (7, 4, 'sp4_r_v_b_45')
// (7, 5, 'neigh_op_top_2')
// (7, 5, 'sp4_r_v_b_32')
// (7, 6, 'lutff_2/out')
// (7, 6, 'sp4_r_v_b_21')
// (7, 7, 'neigh_op_bot_2')
// (7, 7, 'sp4_h_r_36')
// (7, 7, 'sp4_r_v_b_8')
// (8, 3, 'sp4_v_t_45')
// (8, 4, 'sp4_v_b_45')
// (8, 5, 'neigh_op_tnl_2')
// (8, 5, 'sp4_v_b_32')
// (8, 6, 'neigh_op_lft_2')
// (8, 6, 'sp4_v_b_21')
// (8, 7, 'neigh_op_bnl_2')
// (8, 7, 'sp4_h_l_36')
// (8, 7, 'sp4_v_b_8')

wire n711;
// (4, 7, 'sp4_r_v_b_36')
// (4, 7, 'sp4_r_v_b_43')
// (4, 8, 'local_g0_6')
// (4, 8, 'lutff_3/in_1')
// (4, 8, 'lutff_4/in_2')
// (4, 8, 'sp4_r_v_b_25')
// (4, 8, 'sp4_r_v_b_30')
// (4, 9, 'local_g3_3')
// (4, 9, 'lutff_1/in_1')
// (4, 9, 'lutff_2/in_2')
// (4, 9, 'lutff_4/in_0')
// (4, 9, 'lutff_5/in_3')
// (4, 9, 'lutff_6/in_0')
// (4, 9, 'sp4_r_v_b_12')
// (4, 9, 'sp4_r_v_b_19')
// (4, 10, 'sp4_r_v_b_1')
// (4, 10, 'sp4_r_v_b_6')
// (5, 6, 'sp4_v_t_36')
// (5, 6, 'sp4_v_t_43')
// (5, 7, 'sp4_v_b_36')
// (5, 7, 'sp4_v_b_43')
// (5, 8, 'local_g2_6')
// (5, 8, 'lutff_0/in_2')
// (5, 8, 'lutff_2/in_2')
// (5, 8, 'sp4_v_b_25')
// (5, 8, 'sp4_v_b_30')
// (5, 9, 'local_g0_4')
// (5, 9, 'lutff_2/in_2')
// (5, 9, 'lutff_5/in_3')
// (5, 9, 'sp4_v_b_12')
// (5, 9, 'sp4_v_b_19')
// (5, 10, 'local_g1_1')
// (5, 10, 'lutff_0/in_2')
// (5, 10, 'lutff_1/in_1')
// (5, 10, 'lutff_2/in_2')
// (5, 10, 'lutff_3/in_1')
// (5, 10, 'lutff_7/in_3')
// (5, 10, 'sp4_h_r_1')
// (5, 10, 'sp4_v_b_1')
// (5, 10, 'sp4_v_b_6')
// (6, 10, 'sp4_h_r_12')
// (7, 9, 'neigh_op_tnr_2')
// (7, 10, 'local_g3_2')
// (7, 10, 'lutff_1/in_2')
// (7, 10, 'neigh_op_rgt_2')
// (7, 10, 'sp4_h_r_25')
// (7, 10, 'sp4_r_v_b_36')
// (7, 11, 'local_g0_2')
// (7, 11, 'lutff_1/in_3')
// (7, 11, 'lutff_2/in_0')
// (7, 11, 'lutff_5/in_3')
// (7, 11, 'neigh_op_bnr_2')
// (7, 11, 'sp4_r_v_b_25')
// (7, 12, 'sp4_r_v_b_12')
// (7, 13, 'local_g1_1')
// (7, 13, 'lutff_2/in_0')
// (7, 13, 'lutff_5/in_3')
// (7, 13, 'sp4_r_v_b_1')
// (8, 7, 'sp4_r_v_b_40')
// (8, 8, 'sp4_r_v_b_29')
// (8, 9, 'neigh_op_top_2')
// (8, 9, 'sp4_r_v_b_16')
// (8, 9, 'sp4_v_t_36')
// (8, 10, 'local_g1_2')
// (8, 10, 'lutff_0/in_1')
// (8, 10, 'lutff_1/in_0')
// (8, 10, 'lutff_2/out')
// (8, 10, 'lutff_3/in_2')
// (8, 10, 'lutff_7/in_0')
// (8, 10, 'sp4_h_r_36')
// (8, 10, 'sp4_r_v_b_5')
// (8, 10, 'sp4_v_b_36')
// (8, 11, 'local_g0_2')
// (8, 11, 'lutff_1/in_1')
// (8, 11, 'neigh_op_bot_2')
// (8, 11, 'sp4_v_b_25')
// (8, 12, 'sp4_v_b_12')
// (8, 13, 'sp4_v_b_1')
// (9, 6, 'sp4_v_t_40')
// (9, 7, 'sp4_v_b_40')
// (9, 8, 'local_g3_5')
// (9, 8, 'lutff_1/in_1')
// (9, 8, 'sp4_v_b_29')
// (9, 9, 'local_g2_2')
// (9, 9, 'lutff_4/in_2')
// (9, 9, 'neigh_op_tnl_2')
// (9, 9, 'sp4_v_b_16')
// (9, 10, 'local_g0_2')
// (9, 10, 'lutff_0/in_0')
// (9, 10, 'neigh_op_lft_2')
// (9, 10, 'sp4_h_l_36')
// (9, 10, 'sp4_v_b_5')
// (9, 11, 'local_g2_2')
// (9, 11, 'lutff_1/in_3')
// (9, 11, 'lutff_4/in_0')
// (9, 11, 'neigh_op_bnl_2')

wire n712;
// (4, 7, 'sp4_r_v_b_40')
// (4, 8, 'sp4_h_r_5')
// (4, 8, 'sp4_r_v_b_29')
// (4, 9, 'local_g3_0')
// (4, 9, 'lutff_3/in_0')
// (4, 9, 'sp4_r_v_b_16')
// (4, 10, 'sp4_r_v_b_5')
// (5, 6, 'local_g1_5')
// (5, 6, 'lutff_5/in_1')
// (5, 6, 'sp4_h_r_5')
// (5, 6, 'sp4_v_t_40')
// (5, 7, 'sp4_r_v_b_43')
// (5, 7, 'sp4_v_b_40')
// (5, 8, 'local_g1_0')
// (5, 8, 'lutff_1/in_0')
// (5, 8, 'lutff_4/in_3')
// (5, 8, 'lutff_7/in_2')
// (5, 8, 'sp4_h_r_16')
// (5, 8, 'sp4_r_v_b_30')
// (5, 8, 'sp4_v_b_29')
// (5, 9, 'local_g3_3')
// (5, 9, 'lutff_0/in_0')
// (5, 9, 'lutff_1/in_1')
// (5, 9, 'lutff_3/in_3')
// (5, 9, 'sp4_r_v_b_19')
// (5, 9, 'sp4_v_b_16')
// (5, 10, 'sp4_r_v_b_6')
// (5, 10, 'sp4_v_b_5')
// (6, 6, 'sp4_h_r_0')
// (6, 6, 'sp4_h_r_16')
// (6, 6, 'sp4_v_t_43')
// (6, 7, 'sp4_v_b_43')
// (6, 8, 'sp4_h_r_29')
// (6, 8, 'sp4_v_b_30')
// (6, 9, 'sp4_v_b_19')
// (6, 10, 'sp4_v_b_6')
// (7, 5, 'neigh_op_tnr_4')
// (7, 5, 'sp4_r_v_b_37')
// (7, 6, 'neigh_op_rgt_4')
// (7, 6, 'sp4_h_r_13')
// (7, 6, 'sp4_h_r_29')
// (7, 6, 'sp4_r_v_b_24')
// (7, 7, 'local_g1_4')
// (7, 7, 'lutff_3/in_0')
// (7, 7, 'neigh_op_bnr_4')
// (7, 7, 'sp4_r_v_b_13')
// (7, 8, 'sp4_h_r_40')
// (7, 8, 'sp4_r_v_b_0')
// (8, 4, 'sp4_v_t_37')
// (8, 5, 'neigh_op_top_4')
// (8, 5, 'sp4_v_b_37')
// (8, 6, 'lutff_4/out')
// (8, 6, 'sp4_h_r_24')
// (8, 6, 'sp4_h_r_40')
// (8, 6, 'sp4_v_b_24')
// (8, 7, 'neigh_op_bot_4')
// (8, 7, 'sp4_v_b_13')
// (8, 8, 'sp4_h_l_40')
// (8, 8, 'sp4_v_b_0')
// (9, 5, 'neigh_op_tnl_4')
// (9, 6, 'neigh_op_lft_4')
// (9, 6, 'sp4_h_l_40')
// (9, 6, 'sp4_h_r_37')
// (9, 7, 'neigh_op_bnl_4')
// (10, 6, 'sp4_h_l_37')

wire n713;
// (4, 8, 'lutff_1/cout')
// (4, 8, 'lutff_2/in_3')

reg n714 = 0;
// (4, 8, 'neigh_op_tnr_0')
// (4, 9, 'neigh_op_rgt_0')
// (4, 10, 'neigh_op_bnr_0')
// (5, 8, 'neigh_op_top_0')
// (5, 9, 'local_g2_0')
// (5, 9, 'lutff_0/out')
// (5, 9, 'lutff_7/in_3')
// (5, 10, 'neigh_op_bot_0')
// (6, 8, 'neigh_op_tnl_0')
// (6, 9, 'neigh_op_lft_0')
// (6, 10, 'neigh_op_bnl_0')

reg n715 = 0;
// (4, 8, 'neigh_op_tnr_1')
// (4, 9, 'neigh_op_rgt_1')
// (4, 10, 'neigh_op_bnr_1')
// (5, 8, 'neigh_op_top_1')
// (5, 9, 'local_g3_1')
// (5, 9, 'lutff_1/out')
// (5, 9, 'lutff_6/in_0')
// (5, 10, 'neigh_op_bot_1')
// (6, 8, 'neigh_op_tnl_1')
// (6, 9, 'neigh_op_lft_1')
// (6, 10, 'neigh_op_bnl_1')

reg n716 = 0;
// (4, 8, 'neigh_op_tnr_2')
// (4, 9, 'neigh_op_rgt_2')
// (4, 10, 'neigh_op_bnr_2')
// (5, 8, 'local_g0_2')
// (5, 8, 'lutff_3/in_1')
// (5, 8, 'neigh_op_top_2')
// (5, 9, 'lutff_2/out')
// (5, 10, 'neigh_op_bot_2')
// (6, 8, 'neigh_op_tnl_2')
// (6, 9, 'neigh_op_lft_2')
// (6, 10, 'neigh_op_bnl_2')

reg n717 = 0;
// (4, 8, 'neigh_op_tnr_3')
// (4, 9, 'neigh_op_rgt_3')
// (4, 10, 'neigh_op_bnr_3')
// (5, 8, 'neigh_op_top_3')
// (5, 9, 'local_g2_3')
// (5, 9, 'lutff_3/out')
// (5, 9, 'lutff_4/in_3')
// (5, 10, 'neigh_op_bot_3')
// (6, 8, 'neigh_op_tnl_3')
// (6, 9, 'neigh_op_lft_3')
// (6, 10, 'neigh_op_bnl_3')

wire n718;
// (4, 8, 'neigh_op_tnr_4')
// (4, 9, 'neigh_op_rgt_4')
// (4, 10, 'neigh_op_bnr_4')
// (5, 8, 'neigh_op_top_4')
// (5, 9, 'lutff_4/out')
// (5, 9, 'sp4_h_r_8')
// (5, 10, 'neigh_op_bot_4')
// (6, 8, 'neigh_op_tnl_4')
// (6, 9, 'neigh_op_lft_4')
// (6, 9, 'sp4_h_r_21')
// (6, 10, 'neigh_op_bnl_4')
// (7, 9, 'sp4_h_r_32')
// (8, 9, 'sp4_h_r_45')
// (9, 9, 'sp4_h_l_45')
// (9, 9, 'sp4_h_r_11')
// (10, 9, 'sp4_h_r_22')
// (11, 9, 'local_g3_3')
// (11, 9, 'lutff_3/in_1')
// (11, 9, 'sp4_h_r_35')
// (12, 9, 'sp4_h_r_46')
// (13, 9, 'sp4_h_l_46')

reg n719 = 0;
// (4, 8, 'neigh_op_tnr_5')
// (4, 9, 'neigh_op_rgt_5')
// (4, 10, 'neigh_op_bnr_5')
// (5, 8, 'local_g0_5')
// (5, 8, 'lutff_6/in_3')
// (5, 8, 'neigh_op_top_5')
// (5, 9, 'lutff_5/out')
// (5, 10, 'neigh_op_bot_5')
// (6, 8, 'neigh_op_tnl_5')
// (6, 9, 'neigh_op_lft_5')
// (6, 10, 'neigh_op_bnl_5')

wire n720;
// (4, 8, 'neigh_op_tnr_6')
// (4, 9, 'neigh_op_rgt_6')
// (4, 9, 'sp4_h_r_1')
// (4, 10, 'neigh_op_bnr_6')
// (5, 8, 'neigh_op_top_6')
// (5, 9, 'lutff_6/out')
// (5, 9, 'sp4_h_r_12')
// (5, 10, 'neigh_op_bot_6')
// (6, 8, 'neigh_op_tnl_6')
// (6, 9, 'neigh_op_lft_6')
// (6, 9, 'sp4_h_r_25')
// (6, 10, 'neigh_op_bnl_6')
// (7, 9, 'sp4_h_r_36')
// (8, 9, 'sp4_h_l_36')
// (8, 9, 'sp4_h_r_1')
// (9, 9, 'sp4_h_r_12')
// (10, 9, 'local_g3_1')
// (10, 9, 'lutff_2/in_0')
// (10, 9, 'sp4_h_r_25')
// (11, 9, 'sp4_h_r_36')
// (12, 9, 'sp4_h_l_36')

wire n721;
// (4, 8, 'neigh_op_tnr_7')
// (4, 9, 'neigh_op_rgt_7')
// (4, 9, 'sp4_h_r_3')
// (4, 10, 'neigh_op_bnr_7')
// (5, 8, 'neigh_op_top_7')
// (5, 9, 'lutff_7/out')
// (5, 9, 'sp4_h_r_14')
// (5, 10, 'neigh_op_bot_7')
// (6, 8, 'neigh_op_tnl_7')
// (6, 9, 'neigh_op_lft_7')
// (6, 9, 'sp4_h_r_27')
// (6, 10, 'neigh_op_bnl_7')
// (7, 9, 'sp4_h_r_38')
// (8, 9, 'sp4_h_l_38')
// (8, 9, 'sp4_h_r_11')
// (9, 9, 'sp4_h_r_22')
// (10, 9, 'local_g3_3')
// (10, 9, 'lutff_7/in_3')
// (10, 9, 'sp4_h_r_35')
// (11, 9, 'sp4_h_r_46')
// (12, 9, 'sp4_h_l_46')

reg n722 = 0;
// (4, 8, 'sp4_h_r_0')
// (5, 8, 'local_g1_5')
// (5, 8, 'lutff_5/in_3')
// (5, 8, 'sp4_h_r_13')
// (6, 5, 'neigh_op_tnr_7')
// (6, 6, 'neigh_op_rgt_7')
// (6, 7, 'neigh_op_bnr_7')
// (6, 8, 'sp4_h_r_24')
// (7, 5, 'neigh_op_top_7')
// (7, 5, 'sp4_r_v_b_42')
// (7, 6, 'lutff_7/out')
// (7, 6, 'sp4_r_v_b_31')
// (7, 7, 'neigh_op_bot_7')
// (7, 7, 'sp4_r_v_b_18')
// (7, 8, 'sp4_h_r_37')
// (7, 8, 'sp4_r_v_b_7')
// (8, 4, 'sp4_v_t_42')
// (8, 5, 'neigh_op_tnl_7')
// (8, 5, 'sp4_v_b_42')
// (8, 6, 'neigh_op_lft_7')
// (8, 6, 'sp4_v_b_31')
// (8, 7, 'neigh_op_bnl_7')
// (8, 7, 'sp4_v_b_18')
// (8, 8, 'sp4_h_l_37')
// (8, 8, 'sp4_v_b_7')

reg n723 = 0;
// (4, 9, 'neigh_op_tnr_0')
// (4, 10, 'neigh_op_rgt_0')
// (4, 11, 'neigh_op_bnr_0')
// (5, 9, 'local_g1_0')
// (5, 9, 'lutff_6/in_1')
// (5, 9, 'neigh_op_top_0')
// (5, 10, 'lutff_0/out')
// (5, 11, 'neigh_op_bot_0')
// (6, 9, 'neigh_op_tnl_0')
// (6, 10, 'neigh_op_lft_0')
// (6, 11, 'neigh_op_bnl_0')

reg n724 = 0;
// (4, 9, 'neigh_op_tnr_1')
// (4, 10, 'neigh_op_rgt_1')
// (4, 11, 'neigh_op_bnr_1')
// (5, 9, 'local_g0_1')
// (5, 9, 'lutff_7/in_0')
// (5, 9, 'neigh_op_top_1')
// (5, 10, 'lutff_1/out')
// (5, 11, 'neigh_op_bot_1')
// (6, 9, 'neigh_op_tnl_1')
// (6, 10, 'neigh_op_lft_1')
// (6, 11, 'neigh_op_bnl_1')

reg n725 = 0;
// (4, 9, 'neigh_op_tnr_2')
// (4, 10, 'neigh_op_rgt_2')
// (4, 11, 'neigh_op_bnr_2')
// (5, 9, 'local_g0_2')
// (5, 9, 'lutff_4/in_0')
// (5, 9, 'neigh_op_top_2')
// (5, 10, 'lutff_2/out')
// (5, 11, 'neigh_op_bot_2')
// (6, 9, 'neigh_op_tnl_2')
// (6, 10, 'neigh_op_lft_2')
// (6, 11, 'neigh_op_bnl_2')

wire n726;
// (4, 9, 'neigh_op_tnr_3')
// (4, 10, 'neigh_op_rgt_3')
// (4, 11, 'neigh_op_bnr_3')
// (5, 9, 'neigh_op_top_3')
// (5, 10, 'local_g2_3')
// (5, 10, 'lutff_0/in_3')
// (5, 10, 'lutff_3/out')
// (5, 10, 'sp4_h_r_6')
// (5, 11, 'neigh_op_bot_3')
// (6, 9, 'neigh_op_tnl_3')
// (6, 10, 'neigh_op_lft_3')
// (6, 10, 'sp4_h_r_19')
// (6, 11, 'neigh_op_bnl_3')
// (7, 10, 'local_g2_6')
// (7, 10, 'lutff_3/in_3')
// (7, 10, 'sp4_h_r_30')
// (8, 10, 'sp4_h_r_43')
// (9, 10, 'sp4_h_l_43')

reg n727 = 0;
// (4, 9, 'neigh_op_tnr_4')
// (4, 10, 'neigh_op_rgt_4')
// (4, 11, 'neigh_op_bnr_4')
// (5, 9, 'neigh_op_top_4')
// (5, 10, 'lutff_4/out')
// (5, 10, 'sp4_h_r_8')
// (5, 11, 'neigh_op_bot_4')
// (6, 9, 'neigh_op_tnl_4')
// (6, 10, 'neigh_op_lft_4')
// (6, 10, 'sp4_h_r_21')
// (6, 11, 'neigh_op_bnl_4')
// (7, 10, 'sp4_h_r_32')
// (8, 10, 'sp4_h_r_45')
// (9, 10, 'local_g0_0')
// (9, 10, 'lutff_4/in_0')
// (9, 10, 'sp4_h_l_45')
// (9, 10, 'sp4_h_r_8')
// (10, 10, 'sp4_h_r_21')
// (11, 10, 'sp4_h_r_32')
// (12, 10, 'sp4_h_r_45')
// (13, 10, 'sp4_h_l_45')

wire n728;
// (4, 9, 'neigh_op_tnr_7')
// (4, 10, 'neigh_op_rgt_7')
// (4, 11, 'neigh_op_bnr_7')
// (5, 9, 'neigh_op_top_7')
// (5, 10, 'local_g0_7')
// (5, 10, 'lutff_1/in_2')
// (5, 10, 'lutff_4/in_3')
// (5, 10, 'lutff_7/out')
// (5, 11, 'neigh_op_bot_7')
// (6, 9, 'neigh_op_tnl_7')
// (6, 10, 'neigh_op_lft_7')
// (6, 11, 'neigh_op_bnl_7')

wire n729;
// (4, 9, 'sp4_r_v_b_42')
// (4, 10, 'sp4_r_v_b_31')
// (4, 11, 'local_g3_2')
// (4, 11, 'lutff_4/in_1')
// (4, 11, 'lutff_5/in_2')
// (4, 11, 'sp4_r_v_b_18')
// (4, 12, 'sp4_r_v_b_7')
// (5, 8, 'sp4_v_t_42')
// (5, 9, 'sp4_v_b_42')
// (5, 10, 'sp4_v_b_31')
// (5, 11, 'sp4_v_b_18')
// (5, 12, 'sp4_h_r_2')
// (5, 12, 'sp4_v_b_7')
// (6, 12, 'sp4_h_r_15')
// (7, 12, 'sp4_h_r_26')
// (8, 12, 'sp4_h_r_39')
// (9, 12, 'sp4_h_l_39')
// (9, 12, 'sp4_h_r_2')
// (10, 11, 'neigh_op_tnr_5')
// (10, 12, 'neigh_op_rgt_5')
// (10, 12, 'sp4_h_r_15')
// (10, 13, 'neigh_op_bnr_5')
// (11, 11, 'neigh_op_top_5')
// (11, 12, 'lutff_5/out')
// (11, 12, 'sp4_h_r_26')
// (11, 13, 'neigh_op_bot_5')
// (12, 11, 'neigh_op_tnl_5')
// (12, 12, 'neigh_op_lft_5')
// (12, 12, 'sp4_h_r_39')
// (12, 13, 'neigh_op_bnl_5')
// (13, 12, 'sp4_h_l_39')

reg n730 = 0;
// (4, 9, 'sp4_r_v_b_44')
// (4, 10, 'neigh_op_tnr_2')
// (4, 10, 'sp4_r_v_b_33')
// (4, 11, 'neigh_op_rgt_2')
// (4, 11, 'sp4_r_v_b_20')
// (4, 12, 'neigh_op_bnr_2')
// (4, 12, 'sp4_r_v_b_9')
// (5, 8, 'sp4_v_t_44')
// (5, 9, 'sp4_v_b_44')
// (5, 10, 'neigh_op_top_2')
// (5, 10, 'sp4_v_b_33')
// (5, 11, 'local_g2_2')
// (5, 11, 'lutff_2/in_2')
// (5, 11, 'lutff_2/out')
// (5, 11, 'sp4_v_b_20')
// (5, 12, 'neigh_op_bot_2')
// (5, 12, 'sp4_h_r_3')
// (5, 12, 'sp4_v_b_9')
// (6, 10, 'neigh_op_tnl_2')
// (6, 11, 'neigh_op_lft_2')
// (6, 12, 'neigh_op_bnl_2')
// (6, 12, 'sp4_h_r_14')
// (7, 12, 'local_g2_3')
// (7, 12, 'lutff_1/in_2')
// (7, 12, 'sp4_h_r_27')
// (8, 12, 'sp4_h_r_38')
// (9, 12, 'sp4_h_l_38')

reg n731 = 0;
// (4, 10, 'neigh_op_tnr_1')
// (4, 11, 'neigh_op_rgt_1')
// (4, 12, 'neigh_op_bnr_1')
// (5, 9, 'sp4_r_v_b_43')
// (5, 10, 'neigh_op_top_1')
// (5, 10, 'sp4_r_v_b_30')
// (5, 11, 'local_g3_1')
// (5, 11, 'lutff_1/in_1')
// (5, 11, 'lutff_1/out')
// (5, 11, 'sp4_r_v_b_19')
// (5, 12, 'neigh_op_bot_1')
// (5, 12, 'sp4_r_v_b_6')
// (6, 8, 'sp4_v_t_43')
// (6, 9, 'sp4_v_b_43')
// (6, 10, 'neigh_op_tnl_1')
// (6, 10, 'sp4_v_b_30')
// (6, 11, 'neigh_op_lft_1')
// (6, 11, 'sp4_v_b_19')
// (6, 12, 'neigh_op_bnl_1')
// (6, 12, 'sp4_h_r_0')
// (6, 12, 'sp4_v_b_6')
// (7, 12, 'local_g0_5')
// (7, 12, 'lutff_3/in_0')
// (7, 12, 'sp4_h_r_13')
// (8, 12, 'sp4_h_r_24')
// (9, 12, 'sp4_h_r_37')
// (10, 12, 'sp4_h_l_37')

reg n732 = 0;
// (4, 10, 'neigh_op_tnr_3')
// (4, 11, 'neigh_op_rgt_3')
// (4, 12, 'neigh_op_bnr_3')
// (5, 9, 'sp4_r_v_b_47')
// (5, 10, 'neigh_op_top_3')
// (5, 10, 'sp4_r_v_b_34')
// (5, 11, 'local_g1_3')
// (5, 11, 'lutff_3/in_1')
// (5, 11, 'lutff_3/out')
// (5, 11, 'sp4_r_v_b_23')
// (5, 12, 'neigh_op_bot_3')
// (5, 12, 'sp4_r_v_b_10')
// (6, 8, 'sp4_v_t_47')
// (6, 9, 'sp4_v_b_47')
// (6, 10, 'neigh_op_tnl_3')
// (6, 10, 'sp4_v_b_34')
// (6, 11, 'neigh_op_lft_3')
// (6, 11, 'sp4_v_b_23')
// (6, 12, 'neigh_op_bnl_3')
// (6, 12, 'sp4_h_r_4')
// (6, 12, 'sp4_v_b_10')
// (7, 12, 'local_g1_1')
// (7, 12, 'lutff_5/in_3')
// (7, 12, 'sp4_h_r_17')
// (8, 12, 'sp4_h_r_28')
// (9, 12, 'sp4_h_r_41')
// (10, 12, 'sp4_h_l_41')

reg n733 = 0;
// (4, 10, 'neigh_op_tnr_7')
// (4, 11, 'neigh_op_rgt_7')
// (4, 12, 'neigh_op_bnr_7')
// (5, 9, 'sp4_r_v_b_39')
// (5, 10, 'neigh_op_top_7')
// (5, 10, 'sp4_r_v_b_26')
// (5, 11, 'local_g0_7')
// (5, 11, 'local_g3_7')
// (5, 11, 'lutff_0/in_1')
// (5, 11, 'lutff_1/in_3')
// (5, 11, 'lutff_7/in_2')
// (5, 11, 'lutff_7/out')
// (5, 11, 'sp4_r_v_b_15')
// (5, 12, 'neigh_op_bot_7')
// (5, 12, 'sp4_r_v_b_2')
// (6, 8, 'sp4_v_t_39')
// (6, 9, 'sp4_v_b_39')
// (6, 10, 'neigh_op_tnl_7')
// (6, 10, 'sp4_v_b_26')
// (6, 11, 'neigh_op_lft_7')
// (6, 11, 'sp4_v_b_15')
// (6, 12, 'neigh_op_bnl_7')
// (6, 12, 'sp4_h_r_2')
// (6, 12, 'sp4_v_b_2')
// (7, 12, 'sp4_h_r_15')
// (8, 12, 'sp4_h_r_26')
// (9, 12, 'local_g3_7')
// (9, 12, 'lutff_4/in_0')
// (9, 12, 'sp4_h_r_39')
// (10, 12, 'sp4_h_l_39')

wire n734;
// (4, 10, 'sp4_r_v_b_36')
// (4, 11, 'neigh_op_tnr_6')
// (4, 11, 'sp4_r_v_b_25')
// (4, 12, 'neigh_op_rgt_6')
// (4, 12, 'sp4_r_v_b_12')
// (4, 13, 'neigh_op_bnr_6')
// (4, 13, 'sp4_r_v_b_1')
// (5, 9, 'sp4_h_r_6')
// (5, 9, 'sp4_v_t_36')
// (5, 10, 'sp4_v_b_36')
// (5, 11, 'neigh_op_top_6')
// (5, 11, 'sp4_r_v_b_40')
// (5, 11, 'sp4_v_b_25')
// (5, 12, 'lutff_6/out')
// (5, 12, 'sp4_r_v_b_29')
// (5, 12, 'sp4_r_v_b_45')
// (5, 12, 'sp4_v_b_12')
// (5, 13, 'neigh_op_bot_6')
// (5, 13, 'sp4_r_v_b_16')
// (5, 13, 'sp4_r_v_b_32')
// (5, 13, 'sp4_v_b_1')
// (5, 14, 'sp4_r_v_b_21')
// (5, 14, 'sp4_r_v_b_5')
// (5, 15, 'sp4_r_v_b_8')
// (6, 9, 'sp4_h_r_19')
// (6, 10, 'sp4_h_r_10')
// (6, 10, 'sp4_v_t_40')
// (6, 11, 'neigh_op_tnl_6')
// (6, 11, 'sp4_h_r_8')
// (6, 11, 'sp4_v_b_40')
// (6, 11, 'sp4_v_t_45')
// (6, 12, 'neigh_op_lft_6')
// (6, 12, 'sp4_v_b_29')
// (6, 12, 'sp4_v_b_45')
// (6, 13, 'neigh_op_bnl_6')
// (6, 13, 'sp4_v_b_16')
// (6, 13, 'sp4_v_b_32')
// (6, 14, 'sp4_v_b_21')
// (6, 14, 'sp4_v_b_5')
// (6, 15, 'sp4_v_b_8')
// (7, 9, 'sp4_h_r_30')
// (7, 10, 'sp4_h_r_23')
// (7, 11, 'sp4_h_r_21')
// (8, 9, 'sp4_h_r_43')
// (8, 10, 'sp4_h_r_34')
// (8, 11, 'sp4_h_r_32')
// (9, 9, 'sp4_h_l_43')
// (9, 9, 'sp4_h_r_2')
// (9, 10, 'sp4_h_r_47')
// (9, 11, 'sp4_h_r_45')
// (10, 9, 'sp4_h_r_15')
// (10, 10, 'sp4_h_l_47')
// (10, 10, 'sp4_h_r_6')
// (10, 11, 'sp4_h_l_45')
// (10, 11, 'sp4_h_r_11')
// (10, 11, 'sp4_h_r_4')
// (11, 9, 'sp4_h_r_26')
// (11, 10, 'sp4_h_r_19')
// (11, 11, 'sp4_h_r_17')
// (11, 11, 'sp4_h_r_22')
// (12, 9, 'sp4_h_r_39')
// (12, 10, 'sp4_h_r_30')
// (12, 11, 'local_g3_3')
// (12, 11, 'lutff_global/cen')
// (12, 11, 'sp4_h_r_28')
// (12, 11, 'sp4_h_r_35')
// (13, 8, 'sp4_r_v_b_47')
// (13, 9, 'local_g0_2')
// (13, 9, 'lutff_global/cen')
// (13, 9, 'sp4_h_l_39')
// (13, 9, 'sp4_h_r_10')
// (13, 9, 'sp4_r_v_b_34')
// (13, 10, 'local_g3_3')
// (13, 10, 'lutff_global/cen')
// (13, 10, 'sp4_h_r_43')
// (13, 10, 'sp4_r_v_b_23')
// (13, 11, 'local_g2_2')
// (13, 11, 'lutff_global/cen')
// (13, 11, 'sp4_h_r_41')
// (13, 11, 'sp4_h_r_46')
// (13, 11, 'sp4_r_v_b_10')
// (14, 7, 'sp4_v_t_47')
// (14, 8, 'sp4_v_b_47')
// (14, 9, 'sp4_h_r_23')
// (14, 9, 'sp4_v_b_34')
// (14, 10, 'local_g0_2')
// (14, 10, 'lutff_global/cen')
// (14, 10, 'sp4_h_l_43')
// (14, 10, 'sp4_h_r_2')
// (14, 10, 'sp4_v_b_23')
// (14, 11, 'local_g0_2')
// (14, 11, 'lutff_global/cen')
// (14, 11, 'sp4_h_l_41')
// (14, 11, 'sp4_h_l_46')
// (14, 11, 'sp4_v_b_10')
// (15, 9, 'sp4_h_r_34')
// (15, 10, 'sp4_h_r_15')
// (16, 9, 'sp4_h_r_47')
// (16, 10, 'sp4_h_r_26')
// (17, 9, 'sp4_h_l_47')
// (17, 10, 'sp4_h_r_39')
// (18, 10, 'sp4_h_l_39')

wire n735;
// (4, 10, 'sp4_r_v_b_42')
// (4, 11, 'neigh_op_tnr_1')
// (4, 11, 'sp4_r_v_b_31')
// (4, 12, 'neigh_op_rgt_1')
// (4, 12, 'sp4_h_r_7')
// (4, 12, 'sp4_r_v_b_18')
// (4, 13, 'neigh_op_bnr_1')
// (4, 13, 'sp4_r_v_b_7')
// (5, 9, 'sp4_v_t_42')
// (5, 10, 'sp4_r_v_b_43')
// (5, 10, 'sp4_v_b_42')
// (5, 11, 'neigh_op_top_1')
// (5, 11, 'sp4_r_v_b_30')
// (5, 11, 'sp4_v_b_31')
// (5, 12, 'local_g0_1')
// (5, 12, 'lutff_1/out')
// (5, 12, 'lutff_5/in_2')
// (5, 12, 'sp4_h_r_18')
// (5, 12, 'sp4_r_v_b_19')
// (5, 12, 'sp4_v_b_18')
// (5, 13, 'neigh_op_bot_1')
// (5, 13, 'sp4_h_r_7')
// (5, 13, 'sp4_r_v_b_6')
// (5, 13, 'sp4_v_b_7')
// (6, 9, 'sp4_v_t_43')
// (6, 10, 'sp4_v_b_43')
// (6, 11, 'neigh_op_tnl_1')
// (6, 11, 'sp4_v_b_30')
// (6, 12, 'neigh_op_lft_1')
// (6, 12, 'sp4_h_r_31')
// (6, 12, 'sp4_v_b_19')
// (6, 13, 'neigh_op_bnl_1')
// (6, 13, 'sp4_h_r_18')
// (6, 13, 'sp4_h_r_6')
// (6, 13, 'sp4_v_b_6')
// (7, 12, 'sp4_h_r_42')
// (7, 13, 'sp4_h_r_19')
// (7, 13, 'sp4_h_r_31')
// (8, 12, 'sp4_h_l_42')
// (8, 12, 'sp4_h_r_7')
// (8, 13, 'sp4_h_r_30')
// (8, 13, 'sp4_h_r_42')
// (9, 12, 'sp4_h_r_18')
// (9, 13, 'sp4_h_l_42')
// (9, 13, 'sp4_h_r_43')
// (9, 13, 'sp4_h_r_7')
// (10, 12, 'sp4_h_r_31')
// (10, 13, 'sp4_h_l_43')
// (10, 13, 'sp4_h_r_18')
// (10, 13, 'sp4_h_r_2')
// (11, 12, 'sp4_h_r_42')
// (11, 13, 'sp4_h_r_15')
// (11, 13, 'sp4_h_r_31')
// (12, 12, 'sp4_h_l_42')
// (12, 12, 'sp4_h_r_7')
// (12, 13, 'sp4_h_r_26')
// (12, 13, 'sp4_h_r_42')
// (13, 12, 'sp4_h_r_18')
// (13, 13, 'sp4_h_l_42')
// (13, 13, 'sp4_h_r_3')
// (13, 13, 'sp4_h_r_39')
// (14, 12, 'sp4_h_r_31')
// (14, 13, 'local_g0_2')
// (14, 13, 'lutff_global/cen')
// (14, 13, 'sp4_h_l_39')
// (14, 13, 'sp4_h_r_14')
// (14, 13, 'sp4_h_r_2')
// (15, 12, 'local_g2_2')
// (15, 12, 'lutff_global/cen')
// (15, 12, 'sp4_h_r_42')
// (15, 13, 'local_g3_3')
// (15, 13, 'lutff_global/cen')
// (15, 13, 'sp4_h_r_15')
// (15, 13, 'sp4_h_r_27')
// (16, 12, 'sp4_h_l_42')
// (16, 13, 'local_g2_2')
// (16, 13, 'lutff_global/cen')
// (16, 13, 'sp4_h_r_26')
// (16, 13, 'sp4_h_r_38')
// (17, 13, 'sp4_h_l_38')
// (17, 13, 'sp4_h_r_39')
// (18, 13, 'sp4_h_l_39')

wire n736;
// (4, 11, 'local_g3_3')
// (4, 11, 'lutff_4/in_2')
// (4, 11, 'neigh_op_tnr_3')
// (4, 12, 'neigh_op_rgt_3')
// (4, 13, 'neigh_op_bnr_3')
// (5, 11, 'neigh_op_top_3')
// (5, 12, 'lutff_3/out')
// (5, 13, 'neigh_op_bot_3')
// (6, 11, 'neigh_op_tnl_3')
// (6, 12, 'neigh_op_lft_3')
// (6, 13, 'neigh_op_bnl_3')

wire n737;
// (4, 11, 'local_g3_5')
// (4, 11, 'lutff_0/in_0')
// (4, 11, 'lutff_4/in_0')
// (4, 11, 'neigh_op_tnr_5')
// (4, 12, 'neigh_op_rgt_5')
// (4, 13, 'neigh_op_bnr_5')
// (5, 11, 'neigh_op_top_5')
// (5, 12, 'lutff_5/out')
// (5, 13, 'neigh_op_bot_5')
// (6, 11, 'neigh_op_tnl_5')
// (6, 12, 'neigh_op_lft_5')
// (6, 13, 'neigh_op_bnl_5')

reg n738 = 0;
// (4, 11, 'neigh_op_tnr_0')
// (4, 12, 'neigh_op_rgt_0')
// (4, 13, 'neigh_op_bnr_0')
// (5, 11, 'neigh_op_top_0')
// (5, 12, 'lutff_0/out')
// (5, 12, 'sp4_h_r_0')
// (5, 13, 'neigh_op_bot_0')
// (6, 11, 'neigh_op_tnl_0')
// (6, 12, 'neigh_op_lft_0')
// (6, 12, 'sp4_h_r_13')
// (6, 13, 'neigh_op_bnl_0')
// (7, 12, 'local_g3_0')
// (7, 12, 'lutff_2/in_1')
// (7, 12, 'sp4_h_r_24')
// (8, 12, 'sp4_h_r_37')
// (9, 12, 'sp4_h_l_37')

wire n739;
// (4, 11, 'neigh_op_tnr_2')
// (4, 12, 'neigh_op_rgt_2')
// (4, 12, 'sp4_r_v_b_36')
// (4, 13, 'neigh_op_bnr_2')
// (4, 13, 'sp4_r_v_b_25')
// (4, 14, 'sp4_r_v_b_12')
// (4, 15, 'sp4_r_v_b_1')
// (5, 11, 'neigh_op_top_2')
// (5, 11, 'sp4_h_r_1')
// (5, 11, 'sp4_v_t_36')
// (5, 12, 'lutff_2/out')
// (5, 12, 'sp4_v_b_36')
// (5, 13, 'neigh_op_bot_2')
// (5, 13, 'sp4_v_b_25')
// (5, 14, 'sp4_v_b_12')
// (5, 15, 'sp4_v_b_1')
// (6, 11, 'neigh_op_tnl_2')
// (6, 11, 'sp4_h_r_12')
// (6, 12, 'neigh_op_lft_2')
// (6, 13, 'neigh_op_bnl_2')
// (7, 11, 'sp4_h_r_25')
// (8, 11, 'sp4_h_r_36')
// (9, 11, 'sp4_h_l_36')
// (9, 11, 'sp4_h_r_4')
// (10, 11, 'local_g1_1')
// (10, 11, 'lutff_0/in_0')
// (10, 11, 'sp4_h_r_17')
// (11, 11, 'sp4_h_r_28')
// (12, 11, 'sp4_h_r_41')
// (13, 11, 'sp4_h_l_41')

wire n740;
// (4, 12, 'lutff_1/cout')
// (4, 12, 'lutff_2/in_3')

wire n741;
// (4, 12, 'lutff_2/cout')
// (4, 12, 'lutff_3/in_3')

wire n742;
// (4, 12, 'lutff_3/cout')
// (4, 12, 'lutff_4/in_3')

wire n743;
// (4, 12, 'lutff_4/cout')
// (4, 12, 'lutff_5/in_3')

wire n744;
// (4, 12, 'neigh_op_tnr_3')
// (4, 13, 'local_g2_3')
// (4, 13, 'lutff_5/in_0')
// (4, 13, 'neigh_op_rgt_3')
// (4, 14, 'neigh_op_bnr_3')
// (5, 12, 'neigh_op_top_3')
// (5, 13, 'lutff_3/out')
// (5, 14, 'neigh_op_bot_3')
// (6, 12, 'neigh_op_tnl_3')
// (6, 13, 'neigh_op_lft_3')
// (6, 14, 'neigh_op_bnl_3')

wire n745;
// (4, 12, 'neigh_op_tnr_4')
// (4, 13, 'neigh_op_rgt_4')
// (4, 14, 'neigh_op_bnr_4')
// (5, 12, 'neigh_op_top_4')
// (5, 13, 'local_g0_4')
// (5, 13, 'lutff_0/in_0')
// (5, 13, 'lutff_4/out')
// (5, 14, 'neigh_op_bot_4')
// (6, 12, 'neigh_op_tnl_4')
// (6, 13, 'neigh_op_lft_4')
// (6, 14, 'neigh_op_bnl_4')

reg n746 = 0;
// (4, 12, 'neigh_op_tnr_5')
// (4, 13, 'neigh_op_rgt_5')
// (4, 14, 'neigh_op_bnr_5')
// (5, 12, 'neigh_op_top_5')
// (5, 13, 'lutff_5/out')
// (5, 13, 'sp4_h_r_10')
// (5, 14, 'neigh_op_bot_5')
// (6, 12, 'neigh_op_tnl_5')
// (6, 13, 'neigh_op_lft_5')
// (6, 13, 'sp4_h_r_23')
// (6, 14, 'neigh_op_bnl_5')
// (7, 13, 'sp4_h_r_34')
// (8, 13, 'local_g2_7')
// (8, 13, 'lutff_7/in_2')
// (8, 13, 'sp4_h_r_47')
// (9, 13, 'sp4_h_l_47')

wire n747;
// (4, 12, 'neigh_op_tnr_6')
// (4, 13, 'neigh_op_rgt_6')
// (4, 14, 'neigh_op_bnr_6')
// (5, 12, 'neigh_op_top_6')
// (5, 13, 'local_g0_6')
// (5, 13, 'lutff_6/out')
// (5, 13, 'lutff_7/in_1')
// (5, 14, 'neigh_op_bot_6')
// (6, 12, 'neigh_op_tnl_6')
// (6, 13, 'neigh_op_lft_6')
// (6, 14, 'neigh_op_bnl_6')

wire n748;
// (4, 12, 'neigh_op_tnr_7')
// (4, 13, 'neigh_op_rgt_7')
// (4, 14, 'neigh_op_bnr_7')
// (5, 12, 'neigh_op_top_7')
// (5, 13, 'lutff_7/out')
// (5, 14, 'local_g0_7')
// (5, 14, 'local_g1_7')
// (5, 14, 'lutff_2/in_3')
// (5, 14, 'lutff_5/in_3')
// (5, 14, 'neigh_op_bot_7')
// (6, 12, 'neigh_op_tnl_7')
// (6, 13, 'neigh_op_lft_7')
// (6, 14, 'neigh_op_bnl_7')

wire n749;
// (4, 12, 'sp4_h_r_9')
// (5, 12, 'local_g1_4')
// (5, 12, 'lutff_3/in_2')
// (5, 12, 'sp4_h_r_20')
// (6, 11, 'neigh_op_tnr_6')
// (6, 12, 'neigh_op_rgt_6')
// (6, 12, 'sp4_h_r_33')
// (6, 13, 'neigh_op_bnr_6')
// (7, 11, 'neigh_op_top_6')
// (7, 12, 'lutff_6/out')
// (7, 12, 'sp4_h_r_44')
// (7, 13, 'neigh_op_bot_6')
// (8, 11, 'neigh_op_tnl_6')
// (8, 12, 'neigh_op_lft_6')
// (8, 12, 'sp4_h_l_44')
// (8, 13, 'neigh_op_bnl_6')

reg n750 = 0;
// (4, 12, 'sp4_r_v_b_47')
// (4, 13, 'sp4_r_v_b_34')
// (4, 14, 'neigh_op_tnr_5')
// (4, 14, 'sp4_r_v_b_23')
// (4, 15, 'neigh_op_rgt_5')
// (4, 15, 'sp4_r_v_b_10')
// (4, 16, 'neigh_op_bnr_5')
// (5, 11, 'sp4_h_r_3')
// (5, 11, 'sp4_v_t_47')
// (5, 12, 'sp4_v_b_47')
// (5, 13, 'sp4_v_b_34')
// (5, 14, 'neigh_op_top_5')
// (5, 14, 'sp4_v_b_23')
// (5, 15, 'lutff_5/out')
// (5, 15, 'sp4_v_b_10')
// (5, 16, 'neigh_op_bot_5')
// (6, 11, 'sp4_h_r_14')
// (6, 14, 'neigh_op_tnl_5')
// (6, 15, 'neigh_op_lft_5')
// (6, 16, 'neigh_op_bnl_5')
// (7, 11, 'sp4_h_r_27')
// (8, 8, 'sp4_r_v_b_38')
// (8, 9, 'sp4_r_v_b_27')
// (8, 10, 'local_g2_6')
// (8, 10, 'lutff_1/in_3')
// (8, 10, 'sp4_r_v_b_14')
// (8, 11, 'sp4_h_r_38')
// (8, 11, 'sp4_r_v_b_3')
// (9, 7, 'sp4_v_t_38')
// (9, 8, 'sp4_v_b_38')
// (9, 9, 'sp4_v_b_27')
// (9, 10, 'sp4_v_b_14')
// (9, 11, 'sp4_h_l_38')
// (9, 11, 'sp4_v_b_3')

wire n751;
// (4, 13, 'lutff_4/cout')
// (4, 13, 'lutff_5/in_3')

reg n752 = 0;
// (4, 13, 'neigh_op_tnr_0')
// (4, 14, 'local_g2_0')
// (4, 14, 'lutff_6/in_0')
// (4, 14, 'neigh_op_rgt_0')
// (4, 15, 'local_g0_0')
// (4, 15, 'lutff_0/in_0')
// (4, 15, 'neigh_op_bnr_0')
// (5, 13, 'neigh_op_top_0')
// (5, 14, 'local_g3_0')
// (5, 14, 'lutff_0/in_3')
// (5, 14, 'lutff_0/out')
// (5, 14, 'lutff_3/in_2')
// (5, 15, 'local_g1_0')
// (5, 15, 'lutff_1/in_2')
// (5, 15, 'neigh_op_bot_0')
// (6, 13, 'neigh_op_tnl_0')
// (6, 14, 'neigh_op_lft_0')
// (6, 15, 'neigh_op_bnl_0')

reg n753 = 0;
// (4, 13, 'neigh_op_tnr_1')
// (4, 14, 'neigh_op_rgt_1')
// (4, 15, 'neigh_op_bnr_1')
// (5, 13, 'neigh_op_top_1')
// (5, 14, 'local_g0_1')
// (5, 14, 'lutff_1/in_2')
// (5, 14, 'lutff_1/out')
// (5, 14, 'sp4_h_r_2')
// (5, 15, 'local_g0_1')
// (5, 15, 'lutff_6/in_1')
// (5, 15, 'neigh_op_bot_1')
// (6, 13, 'neigh_op_tnl_1')
// (6, 14, 'neigh_op_lft_1')
// (6, 14, 'sp4_h_r_15')
// (6, 15, 'neigh_op_bnl_1')
// (7, 14, 'sp4_h_r_26')
// (8, 14, 'sp4_h_r_39')
// (8, 15, 'sp4_r_v_b_42')
// (8, 16, 'sp4_r_v_b_31')
// (8, 17, 'sp4_r_v_b_18')
// (8, 18, 'sp4_r_v_b_7')
// (9, 14, 'sp4_h_l_39')
// (9, 14, 'sp4_v_t_42')
// (9, 15, 'local_g2_2')
// (9, 15, 'lutff_6/in_2')
// (9, 15, 'sp4_v_b_42')
// (9, 16, 'sp4_v_b_31')
// (9, 17, 'sp4_v_b_18')
// (9, 18, 'sp4_v_b_7')

wire n754;
// (4, 13, 'neigh_op_tnr_3')
// (4, 14, 'neigh_op_rgt_3')
// (4, 15, 'neigh_op_bnr_3')
// (5, 13, 'local_g0_3')
// (5, 13, 'lutff_2/in_3')
// (5, 13, 'neigh_op_top_3')
// (5, 14, 'lutff_3/out')
// (5, 14, 'sp4_h_r_6')
// (5, 15, 'neigh_op_bot_3')
// (6, 13, 'neigh_op_tnl_3')
// (6, 14, 'neigh_op_lft_3')
// (6, 14, 'sp4_h_r_19')
// (6, 15, 'neigh_op_bnl_3')
// (7, 14, 'sp4_h_r_30')
// (8, 14, 'local_g3_3')
// (8, 14, 'lutff_global/cen')
// (8, 14, 'sp4_h_r_43')
// (9, 14, 'sp4_h_l_43')

wire n755;
// (4, 13, 'neigh_op_tnr_4')
// (4, 14, 'local_g3_4')
// (4, 14, 'lutff_5/in_0')
// (4, 14, 'neigh_op_rgt_4')
// (4, 15, 'neigh_op_bnr_4')
// (5, 13, 'neigh_op_top_4')
// (5, 13, 'sp4_r_v_b_36')
// (5, 14, 'lutff_4/out')
// (5, 14, 'sp4_r_v_b_25')
// (5, 15, 'neigh_op_bot_4')
// (5, 15, 'sp4_r_v_b_12')
// (5, 16, 'sp4_r_v_b_1')
// (6, 12, 'sp4_h_r_6')
// (6, 12, 'sp4_v_t_36')
// (6, 13, 'neigh_op_tnl_4')
// (6, 13, 'sp4_v_b_36')
// (6, 14, 'neigh_op_lft_4')
// (6, 14, 'sp4_v_b_25')
// (6, 15, 'neigh_op_bnl_4')
// (6, 15, 'sp4_v_b_12')
// (6, 16, 'sp4_v_b_1')
// (7, 12, 'sp4_h_r_19')
// (8, 12, 'sp4_h_r_30')
// (9, 12, 'sp4_h_r_43')
// (10, 12, 'sp4_h_l_43')
// (10, 12, 'sp4_h_r_6')
// (11, 12, 'sp4_h_r_19')
// (12, 12, 'sp4_h_r_30')
// (13, 12, 'local_g3_3')
// (13, 12, 'lutff_global/cen')
// (13, 12, 'sp4_h_r_43')
// (14, 12, 'sp4_h_l_43')

wire n756;
// (4, 13, 'neigh_op_tnr_7')
// (4, 14, 'neigh_op_rgt_7')
// (4, 15, 'local_g1_7')
// (4, 15, 'lutff_3/in_1')
// (4, 15, 'lutff_4/in_2')
// (4, 15, 'lutff_5/in_1')
// (4, 15, 'lutff_6/in_2')
// (4, 15, 'neigh_op_bnr_7')
// (5, 13, 'neigh_op_top_7')
// (5, 14, 'local_g2_7')
// (5, 14, 'lutff_1/in_0')
// (5, 14, 'lutff_7/out')
// (5, 15, 'local_g0_7')
// (5, 15, 'lutff_0/in_3')
// (5, 15, 'lutff_2/in_1')
// (5, 15, 'lutff_4/in_1')
// (5, 15, 'lutff_6/in_3')
// (5, 15, 'neigh_op_bot_7')
// (6, 13, 'neigh_op_tnl_7')
// (6, 14, 'neigh_op_lft_7')
// (6, 15, 'neigh_op_bnl_7')

reg n757 = 0;
// (4, 13, 'sp4_r_v_b_40')
// (4, 14, 'neigh_op_tnr_0')
// (4, 14, 'sp4_r_v_b_29')
// (4, 15, 'neigh_op_rgt_0')
// (4, 15, 'sp4_r_v_b_16')
// (4, 16, 'neigh_op_bnr_0')
// (4, 16, 'sp4_r_v_b_5')
// (5, 12, 'sp4_h_r_10')
// (5, 12, 'sp4_v_t_40')
// (5, 13, 'sp4_v_b_40')
// (5, 14, 'neigh_op_top_0')
// (5, 14, 'sp4_v_b_29')
// (5, 15, 'lutff_0/out')
// (5, 15, 'sp4_v_b_16')
// (5, 16, 'neigh_op_bot_0')
// (5, 16, 'sp4_v_b_5')
// (6, 12, 'sp4_h_r_23')
// (6, 14, 'neigh_op_tnl_0')
// (6, 15, 'neigh_op_lft_0')
// (6, 16, 'neigh_op_bnl_0')
// (7, 12, 'sp4_h_r_34')
// (8, 9, 'sp4_r_v_b_47')
// (8, 10, 'local_g2_2')
// (8, 10, 'lutff_0/in_2')
// (8, 10, 'sp4_r_v_b_34')
// (8, 11, 'sp4_r_v_b_23')
// (8, 12, 'sp4_h_r_47')
// (8, 12, 'sp4_r_v_b_10')
// (9, 8, 'sp4_v_t_47')
// (9, 9, 'sp4_v_b_47')
// (9, 10, 'sp4_v_b_34')
// (9, 11, 'sp4_v_b_23')
// (9, 12, 'sp4_h_l_47')
// (9, 12, 'sp4_v_b_10')

wire n758;
// (4, 14, 'neigh_op_tnr_1')
// (4, 15, 'local_g3_1')
// (4, 15, 'lutff_4/in_0')
// (4, 15, 'neigh_op_rgt_1')
// (4, 16, 'local_g1_1')
// (4, 16, 'lutff_4/in_2')
// (4, 16, 'neigh_op_bnr_1')
// (5, 14, 'neigh_op_top_1')
// (5, 15, 'lutff_1/out')
// (5, 16, 'local_g0_1')
// (5, 16, 'lutff_5/in_0')
// (5, 16, 'neigh_op_bot_1')
// (6, 14, 'neigh_op_tnl_1')
// (6, 15, 'neigh_op_lft_1')
// (6, 16, 'neigh_op_bnl_1')

reg n759 = 0;
// (4, 14, 'neigh_op_tnr_2')
// (4, 15, 'neigh_op_rgt_2')
// (4, 15, 'sp4_h_r_9')
// (4, 16, 'neigh_op_bnr_2')
// (5, 14, 'neigh_op_top_2')
// (5, 15, 'lutff_2/out')
// (5, 15, 'sp4_h_r_20')
// (5, 16, 'neigh_op_bot_2')
// (6, 14, 'neigh_op_tnl_2')
// (6, 15, 'neigh_op_lft_2')
// (6, 15, 'sp4_h_r_33')
// (6, 16, 'neigh_op_bnl_2')
// (7, 12, 'sp4_r_v_b_38')
// (7, 13, 'local_g1_3')
// (7, 13, 'lutff_3/in_3')
// (7, 13, 'sp4_r_v_b_27')
// (7, 14, 'sp4_r_v_b_14')
// (7, 15, 'sp4_h_r_44')
// (7, 15, 'sp4_r_v_b_3')
// (8, 11, 'sp4_v_t_38')
// (8, 12, 'sp4_v_b_38')
// (8, 13, 'sp4_v_b_27')
// (8, 14, 'sp4_v_b_14')
// (8, 15, 'sp4_h_l_44')
// (8, 15, 'sp4_v_b_3')

wire n760;
// (4, 14, 'neigh_op_tnr_3')
// (4, 15, 'neigh_op_rgt_3')
// (4, 16, 'neigh_op_bnr_3')
// (5, 14, 'neigh_op_top_3')
// (5, 15, 'lutff_3/out')
// (5, 16, 'local_g0_3')
// (5, 16, 'lutff_0/in_1')
// (5, 16, 'neigh_op_bot_3')
// (6, 14, 'neigh_op_tnl_3')
// (6, 15, 'neigh_op_lft_3')
// (6, 16, 'neigh_op_bnl_3')

reg n761 = 0;
// (4, 14, 'neigh_op_tnr_7')
// (4, 15, 'neigh_op_rgt_7')
// (4, 16, 'neigh_op_bnr_7')
// (5, 11, 'sp4_r_v_b_36')
// (5, 12, 'sp4_r_v_b_25')
// (5, 13, 'sp4_r_v_b_12')
// (5, 14, 'neigh_op_top_7')
// (5, 14, 'sp4_r_v_b_1')
// (5, 15, 'lutff_7/out')
// (5, 15, 'sp4_r_v_b_47')
// (5, 16, 'neigh_op_bot_7')
// (5, 16, 'sp4_r_v_b_34')
// (5, 17, 'sp4_r_v_b_23')
// (5, 18, 'sp4_r_v_b_10')
// (6, 10, 'sp4_h_r_1')
// (6, 10, 'sp4_v_t_36')
// (6, 11, 'sp4_v_b_36')
// (6, 12, 'sp4_v_b_25')
// (6, 13, 'sp4_v_b_12')
// (6, 14, 'neigh_op_tnl_7')
// (6, 14, 'sp4_v_b_1')
// (6, 14, 'sp4_v_t_47')
// (6, 15, 'neigh_op_lft_7')
// (6, 15, 'sp4_v_b_47')
// (6, 16, 'neigh_op_bnl_7')
// (6, 16, 'sp4_v_b_34')
// (6, 17, 'sp4_v_b_23')
// (6, 18, 'sp4_v_b_10')
// (7, 10, 'sp4_h_r_12')
// (8, 10, 'local_g3_1')
// (8, 10, 'lutff_3/in_1')
// (8, 10, 'sp4_h_r_25')
// (9, 10, 'sp4_h_r_36')
// (10, 10, 'sp4_h_l_36')

wire n762;
// (4, 14, 'sp4_h_r_4')
// (5, 14, 'sp4_h_r_17')
// (6, 14, 'sp4_h_r_28')
// (7, 14, 'sp4_h_r_41')
// (8, 14, 'sp4_h_l_41')
// (8, 14, 'sp4_h_r_1')
// (8, 14, 'sp4_h_r_7')
// (9, 14, 'local_g0_2')
// (9, 14, 'lutff_global/cen')
// (9, 14, 'sp4_h_r_12')
// (9, 14, 'sp4_h_r_18')
// (10, 11, 'sp4_r_v_b_41')
// (10, 12, 'sp4_r_v_b_28')
// (10, 13, 'neigh_op_tnr_2')
// (10, 13, 'sp4_r_v_b_17')
// (10, 14, 'neigh_op_rgt_2')
// (10, 14, 'sp4_h_r_25')
// (10, 14, 'sp4_h_r_31')
// (10, 14, 'sp4_r_v_b_4')
// (10, 15, 'neigh_op_bnr_2')
// (10, 15, 'sp4_r_v_b_42')
// (10, 16, 'sp4_r_v_b_31')
// (10, 17, 'sp4_r_v_b_18')
// (10, 18, 'sp4_r_v_b_7')
// (11, 10, 'sp4_v_t_41')
// (11, 11, 'sp4_v_b_41')
// (11, 12, 'sp4_v_b_28')
// (11, 13, 'neigh_op_top_2')
// (11, 13, 'sp4_v_b_17')
// (11, 14, 'lutff_2/out')
// (11, 14, 'sp4_h_r_36')
// (11, 14, 'sp4_h_r_42')
// (11, 14, 'sp4_v_b_4')
// (11, 14, 'sp4_v_t_42')
// (11, 15, 'neigh_op_bot_2')
// (11, 15, 'sp4_v_b_42')
// (11, 16, 'sp4_v_b_31')
// (11, 17, 'local_g0_2')
// (11, 17, 'lutff_global/cen')
// (11, 17, 'sp4_v_b_18')
// (11, 18, 'sp4_v_b_7')
// (12, 13, 'neigh_op_tnl_2')
// (12, 14, 'neigh_op_lft_2')
// (12, 14, 'sp4_h_l_36')
// (12, 14, 'sp4_h_l_42')
// (12, 15, 'neigh_op_bnl_2')

wire n763;
// (4, 15, 'neigh_op_tnr_2')
// (4, 16, 'neigh_op_rgt_2')
// (4, 17, 'neigh_op_bnr_2')
// (5, 15, 'neigh_op_top_2')
// (5, 16, 'lutff_2/out')
// (5, 17, 'local_g0_2')
// (5, 17, 'lutff_4/in_2')
// (5, 17, 'neigh_op_bot_2')
// (6, 15, 'neigh_op_tnl_2')
// (6, 16, 'neigh_op_lft_2')
// (6, 17, 'neigh_op_bnl_2')

reg n764 = 0;
// (4, 15, 'neigh_op_tnr_3')
// (4, 16, 'neigh_op_rgt_3')
// (4, 17, 'neigh_op_bnr_3')
// (5, 9, 'sp4_r_v_b_38')
// (5, 9, 'sp4_r_v_b_42')
// (5, 10, 'sp4_r_v_b_27')
// (5, 10, 'sp4_r_v_b_31')
// (5, 11, 'local_g2_6')
// (5, 11, 'local_g3_2')
// (5, 11, 'lutff_1/in_0')
// (5, 11, 'lutff_2/in_0')
// (5, 11, 'lutff_3/in_0')
// (5, 11, 'lutff_4/in_1')
// (5, 11, 'lutff_7/in_3')
// (5, 11, 'sp4_r_v_b_14')
// (5, 11, 'sp4_r_v_b_18')
// (5, 12, 'sp4_r_v_b_3')
// (5, 12, 'sp4_r_v_b_7')
// (5, 13, 'sp4_r_v_b_42')
// (5, 14, 'sp4_r_v_b_31')
// (5, 15, 'neigh_op_top_3')
// (5, 15, 'sp4_r_v_b_18')
// (5, 16, 'lutff_3/out')
// (5, 16, 'sp4_r_v_b_7')
// (5, 17, 'neigh_op_bot_3')
// (6, 8, 'sp4_v_t_38')
// (6, 8, 'sp4_v_t_42')
// (6, 9, 'sp4_v_b_38')
// (6, 9, 'sp4_v_b_42')
// (6, 10, 'sp4_v_b_27')
// (6, 10, 'sp4_v_b_31')
// (6, 11, 'sp4_v_b_14')
// (6, 11, 'sp4_v_b_18')
// (6, 12, 'sp4_v_b_3')
// (6, 12, 'sp4_v_b_7')
// (6, 12, 'sp4_v_t_42')
// (6, 13, 'sp4_v_b_42')
// (6, 14, 'sp4_v_b_31')
// (6, 15, 'neigh_op_tnl_3')
// (6, 15, 'sp4_v_b_18')
// (6, 16, 'neigh_op_lft_3')
// (6, 16, 'sp4_v_b_7')
// (6, 17, 'neigh_op_bnl_3')

wire n765;
// (4, 15, 'neigh_op_tnr_4')
// (4, 16, 'neigh_op_rgt_4')
// (4, 17, 'neigh_op_bnr_4')
// (5, 15, 'neigh_op_top_4')
// (5, 16, 'lutff_4/out')
// (5, 16, 'sp4_r_v_b_41')
// (5, 17, 'neigh_op_bot_4')
// (5, 17, 'sp4_r_v_b_28')
// (5, 18, 'sp4_r_v_b_17')
// (5, 19, 'local_g1_4')
// (5, 19, 'lutff_3/in_0')
// (5, 19, 'sp4_r_v_b_4')
// (6, 15, 'neigh_op_tnl_4')
// (6, 15, 'sp4_v_t_41')
// (6, 16, 'neigh_op_lft_4')
// (6, 16, 'sp4_v_b_41')
// (6, 17, 'neigh_op_bnl_4')
// (6, 17, 'sp4_v_b_28')
// (6, 18, 'sp4_v_b_17')
// (6, 19, 'sp4_v_b_4')

wire n766;
// (4, 15, 'neigh_op_tnr_5')
// (4, 16, 'neigh_op_rgt_5')
// (4, 17, 'neigh_op_bnr_5')
// (5, 15, 'neigh_op_top_5')
// (5, 16, 'local_g2_5')
// (5, 16, 'lutff_3/in_2')
// (5, 16, 'lutff_5/out')
// (5, 16, 'lutff_6/in_1')
// (5, 17, 'neigh_op_bot_5')
// (6, 15, 'neigh_op_tnl_5')
// (6, 16, 'neigh_op_lft_5')
// (6, 17, 'neigh_op_bnl_5')

wire n767;
// (4, 15, 'neigh_op_tnr_7')
// (4, 16, 'neigh_op_rgt_7')
// (4, 17, 'neigh_op_bnr_7')
// (5, 15, 'neigh_op_top_7')
// (5, 16, 'local_g1_7')
// (5, 16, 'lutff_2/in_2')
// (5, 16, 'lutff_7/out')
// (5, 17, 'local_g0_7')
// (5, 17, 'lutff_7/in_2')
// (5, 17, 'neigh_op_bot_7')
// (6, 15, 'neigh_op_tnl_7')
// (6, 16, 'neigh_op_lft_7')
// (6, 17, 'neigh_op_bnl_7')

wire n768;
// (4, 16, 'neigh_op_tnr_0')
// (4, 17, 'neigh_op_rgt_0')
// (4, 18, 'neigh_op_bnr_0')
// (5, 16, 'neigh_op_top_0')
// (5, 17, 'lutff_0/out')
// (5, 17, 'sp4_h_r_0')
// (5, 18, 'neigh_op_bot_0')
// (6, 16, 'neigh_op_tnl_0')
// (6, 17, 'neigh_op_lft_0')
// (6, 17, 'sp4_h_r_13')
// (6, 18, 'neigh_op_bnl_0')
// (7, 17, 'sp4_h_r_24')
// (8, 17, 'sp4_h_r_37')
// (8, 18, 'sp4_r_v_b_40')
// (8, 19, 'sp4_r_v_b_29')
// (8, 20, 'sp4_r_v_b_16')
// (8, 21, 'local_g1_5')
// (8, 21, 'lutff_4/in_2')
// (8, 21, 'sp4_r_v_b_5')
// (9, 17, 'sp4_h_l_37')
// (9, 17, 'sp4_v_t_40')
// (9, 18, 'sp4_v_b_40')
// (9, 19, 'sp4_v_b_29')
// (9, 20, 'sp4_v_b_16')
// (9, 21, 'sp4_v_b_5')

reg n769 = 0;
// (4, 16, 'neigh_op_tnr_1')
// (4, 17, 'neigh_op_rgt_1')
// (4, 18, 'neigh_op_bnr_1')
// (5, 16, 'neigh_op_top_1')
// (5, 17, 'lutff_1/out')
// (5, 17, 'sp4_h_r_2')
// (5, 18, 'neigh_op_bot_1')
// (6, 16, 'neigh_op_tnl_1')
// (6, 17, 'neigh_op_lft_1')
// (6, 17, 'sp4_h_r_15')
// (6, 18, 'neigh_op_bnl_1')
// (7, 17, 'local_g3_2')
// (7, 17, 'lutff_5/in_2')
// (7, 17, 'sp4_h_r_26')
// (8, 17, 'sp4_h_r_39')
// (9, 17, 'sp4_h_l_39')

wire n770;
// (4, 16, 'neigh_op_tnr_3')
// (4, 17, 'neigh_op_rgt_3')
// (4, 18, 'neigh_op_bnr_3')
// (5, 16, 'neigh_op_top_3')
// (5, 17, 'local_g3_3')
// (5, 17, 'lutff_3/out')
// (5, 17, 'lutff_5/in_1')
// (5, 18, 'neigh_op_bot_3')
// (6, 16, 'neigh_op_tnl_3')
// (6, 17, 'neigh_op_lft_3')
// (6, 18, 'neigh_op_bnl_3')

wire n771;
// (4, 16, 'neigh_op_tnr_4')
// (4, 17, 'neigh_op_rgt_4')
// (4, 18, 'neigh_op_bnr_4')
// (5, 16, 'neigh_op_top_4')
// (5, 17, 'lutff_4/out')
// (5, 17, 'sp4_h_r_8')
// (5, 18, 'neigh_op_bot_4')
// (6, 16, 'neigh_op_tnl_4')
// (6, 17, 'neigh_op_lft_4')
// (6, 17, 'sp4_h_r_21')
// (6, 18, 'neigh_op_bnl_4')
// (7, 17, 'sp4_h_r_32')
// (8, 17, 'sp4_h_r_45')
// (8, 18, 'sp4_r_v_b_45')
// (8, 19, 'sp4_r_v_b_32')
// (8, 20, 'sp4_r_v_b_21')
// (8, 21, 'local_g2_0')
// (8, 21, 'lutff_3/in_1')
// (8, 21, 'sp4_r_v_b_8')
// (9, 17, 'sp4_h_l_45')
// (9, 17, 'sp4_v_t_45')
// (9, 18, 'sp4_v_b_45')
// (9, 19, 'sp4_v_b_32')
// (9, 20, 'sp4_v_b_21')
// (9, 21, 'sp4_v_b_8')

reg n772 = 0;
// (4, 16, 'neigh_op_tnr_5')
// (4, 17, 'local_g2_5')
// (4, 17, 'lutff_2/in_1')
// (4, 17, 'neigh_op_rgt_5')
// (4, 18, 'neigh_op_bnr_5')
// (5, 16, 'neigh_op_top_5')
// (5, 17, 'local_g1_5')
// (5, 17, 'local_g2_5')
// (5, 17, 'lutff_3/in_3')
// (5, 17, 'lutff_5/out')
// (5, 17, 'lutff_7/in_0')
// (5, 18, 'neigh_op_bot_5')
// (6, 16, 'neigh_op_tnl_5')
// (6, 17, 'neigh_op_lft_5')
// (6, 18, 'neigh_op_bnl_5')

reg n773 = 0;
// (4, 16, 'neigh_op_tnr_7')
// (4, 17, 'neigh_op_rgt_7')
// (4, 18, 'neigh_op_bnr_7')
// (5, 16, 'neigh_op_top_7')
// (5, 17, 'local_g1_7')
// (5, 17, 'lutff_3/in_1')
// (5, 17, 'lutff_7/in_1')
// (5, 17, 'lutff_7/out')
// (5, 18, 'neigh_op_bot_7')
// (6, 16, 'neigh_op_tnl_7')
// (6, 17, 'neigh_op_lft_7')
// (6, 18, 'neigh_op_bnl_7')

wire n774;
// (4, 17, 'neigh_op_tnr_1')
// (4, 18, 'neigh_op_rgt_1')
// (4, 19, 'neigh_op_bnr_1')
// (5, 17, 'neigh_op_top_1')
// (5, 18, 'local_g1_1')
// (5, 18, 'lutff_0/in_0')
// (5, 18, 'lutff_1/out')
// (5, 19, 'neigh_op_bot_1')
// (6, 17, 'neigh_op_tnl_1')
// (6, 18, 'neigh_op_lft_1')
// (6, 19, 'neigh_op_bnl_1')

wire n775;
// (4, 17, 'neigh_op_tnr_3')
// (4, 18, 'neigh_op_rgt_3')
// (4, 19, 'neigh_op_bnr_3')
// (5, 17, 'neigh_op_top_3')
// (5, 18, 'local_g2_3')
// (5, 18, 'lutff_3/out')
// (5, 18, 'lutff_6/in_3')
// (5, 19, 'neigh_op_bot_3')
// (6, 17, 'neigh_op_tnl_3')
// (6, 18, 'neigh_op_lft_3')
// (6, 19, 'neigh_op_bnl_3')

wire n776;
// (4, 17, 'neigh_op_tnr_4')
// (4, 18, 'neigh_op_rgt_4')
// (4, 19, 'neigh_op_bnr_4')
// (5, 17, 'neigh_op_top_4')
// (5, 18, 'lutff_4/out')
// (5, 19, 'local_g0_4')
// (5, 19, 'lutff_2/in_2')
// (5, 19, 'neigh_op_bot_4')
// (6, 17, 'neigh_op_tnl_4')
// (6, 18, 'neigh_op_lft_4')
// (6, 19, 'neigh_op_bnl_4')

reg n777 = 0;
// (4, 18, 'local_g2_2')
// (4, 18, 'lutff_3/in_1')
// (4, 18, 'neigh_op_tnr_2')
// (4, 19, 'neigh_op_rgt_2')
// (4, 19, 'sp4_h_r_9')
// (4, 19, 'sp4_r_v_b_36')
// (4, 20, 'neigh_op_bnr_2')
// (4, 20, 'sp4_r_v_b_25')
// (4, 21, 'local_g2_4')
// (4, 21, 'lutff_2/in_2')
// (4, 21, 'sp4_r_v_b_12')
// (4, 22, 'sp4_r_v_b_1')
// (5, 12, 'sp4_r_v_b_40')
// (5, 13, 'sp4_r_v_b_29')
// (5, 14, 'sp4_r_v_b_16')
// (5, 15, 'sp4_r_v_b_5')
// (5, 16, 'sp4_r_v_b_40')
// (5, 17, 'sp4_r_v_b_29')
// (5, 18, 'local_g0_2')
// (5, 18, 'lutff_4/in_0')
// (5, 18, 'neigh_op_top_2')
// (5, 18, 'sp4_r_v_b_16')
// (5, 18, 'sp4_v_t_36')
// (5, 19, 'lutff_2/out')
// (5, 19, 'sp4_h_r_20')
// (5, 19, 'sp4_h_r_4')
// (5, 19, 'sp4_r_v_b_5')
// (5, 19, 'sp4_v_b_36')
// (5, 20, 'neigh_op_bot_2')
// (5, 20, 'sp4_v_b_25')
// (5, 21, 'sp4_v_b_12')
// (5, 22, 'sp4_v_b_1')
// (6, 11, 'sp4_h_r_10')
// (6, 11, 'sp4_v_t_40')
// (6, 12, 'sp4_v_b_40')
// (6, 13, 'sp4_v_b_29')
// (6, 14, 'sp4_v_b_16')
// (6, 15, 'sp4_v_b_5')
// (6, 15, 'sp4_v_t_40')
// (6, 16, 'sp4_v_b_40')
// (6, 17, 'sp4_v_b_29')
// (6, 18, 'neigh_op_tnl_2')
// (6, 18, 'sp4_v_b_16')
// (6, 19, 'neigh_op_lft_2')
// (6, 19, 'sp4_h_r_17')
// (6, 19, 'sp4_h_r_33')
// (6, 19, 'sp4_v_b_5')
// (6, 20, 'neigh_op_bnl_2')
// (7, 11, 'sp4_h_r_23')
// (7, 16, 'sp4_r_v_b_38')
// (7, 17, 'local_g1_3')
// (7, 17, 'lutff_0/in_2')
// (7, 17, 'sp4_r_v_b_27')
// (7, 18, 'sp4_r_v_b_14')
// (7, 19, 'sp4_h_r_28')
// (7, 19, 'sp4_h_r_44')
// (7, 19, 'sp4_r_v_b_3')
// (8, 11, 'local_g2_2')
// (8, 11, 'lutff_2/in_0')
// (8, 11, 'sp4_h_r_34')
// (8, 12, 'sp4_r_v_b_42')
// (8, 13, 'sp4_r_v_b_31')
// (8, 14, 'local_g3_2')
// (8, 14, 'lutff_3/in_0')
// (8, 14, 'sp4_r_v_b_18')
// (8, 15, 'sp4_r_v_b_7')
// (8, 15, 'sp4_v_t_38')
// (8, 16, 'sp4_r_v_b_41')
// (8, 16, 'sp4_v_b_38')
// (8, 17, 'sp4_r_v_b_28')
// (8, 17, 'sp4_v_b_27')
// (8, 18, 'local_g3_1')
// (8, 18, 'lutff_7/in_3')
// (8, 18, 'sp4_r_v_b_17')
// (8, 18, 'sp4_v_b_14')
// (8, 19, 'sp4_h_l_44')
// (8, 19, 'sp4_h_r_41')
// (8, 19, 'sp4_r_v_b_4')
// (8, 19, 'sp4_v_b_3')
// (9, 11, 'sp4_h_r_47')
// (9, 11, 'sp4_v_t_42')
// (9, 12, 'sp4_v_b_42')
// (9, 13, 'sp4_v_b_31')
// (9, 14, 'sp4_v_b_18')
// (9, 15, 'sp4_v_b_7')
// (9, 15, 'sp4_v_t_41')
// (9, 16, 'sp4_v_b_41')
// (9, 17, 'sp4_v_b_28')
// (9, 18, 'sp4_v_b_17')
// (9, 19, 'sp4_h_l_41')
// (9, 19, 'sp4_v_b_4')
// (10, 11, 'sp4_h_l_47')

wire n778;
// (4, 18, 'lutff_1/cout')
// (4, 18, 'lutff_2/in_3')

wire n779;
// (4, 18, 'lutff_3/cout')
// (4, 18, 'lutff_4/in_3')

wire n780;
// (4, 18, 'lutff_5/cout')
// (4, 18, 'lutff_6/in_3')

wire n781;
// (4, 18, 'lutff_7/cout')
// (4, 19, 'carry_in')
// (4, 19, 'carry_in_mux')
// (4, 19, 'lutff_0/in_3')

wire n782;
// (4, 18, 'neigh_op_tnr_0')
// (4, 19, 'neigh_op_rgt_0')
// (4, 20, 'neigh_op_bnr_0')
// (5, 18, 'neigh_op_top_0')
// (5, 19, 'local_g1_0')
// (5, 19, 'lutff_0/out')
// (5, 19, 'lutff_7/in_0')
// (5, 20, 'neigh_op_bot_0')
// (6, 18, 'neigh_op_tnl_0')
// (6, 19, 'neigh_op_lft_0')
// (6, 20, 'neigh_op_bnl_0')

wire n783;
// (4, 18, 'neigh_op_tnr_1')
// (4, 19, 'local_g2_1')
// (4, 19, 'lutff_5/in_2')
// (4, 19, 'neigh_op_rgt_1')
// (4, 20, 'neigh_op_bnr_1')
// (5, 18, 'neigh_op_top_1')
// (5, 19, 'lutff_1/out')
// (5, 20, 'neigh_op_bot_1')
// (6, 18, 'neigh_op_tnl_1')
// (6, 19, 'neigh_op_lft_1')
// (6, 20, 'neigh_op_bnl_1')

wire n784;
// (4, 18, 'neigh_op_tnr_3')
// (4, 19, 'local_g3_3')
// (4, 19, 'lutff_7/in_3')
// (4, 19, 'neigh_op_rgt_3')
// (4, 20, 'neigh_op_bnr_3')
// (5, 18, 'neigh_op_top_3')
// (5, 19, 'local_g3_3')
// (5, 19, 'lutff_3/out')
// (5, 19, 'lutff_5/in_1')
// (5, 20, 'neigh_op_bot_3')
// (6, 18, 'neigh_op_tnl_3')
// (6, 19, 'neigh_op_lft_3')
// (6, 20, 'neigh_op_bnl_3')

wire n785;
// (4, 18, 'neigh_op_tnr_4')
// (4, 19, 'local_g2_4')
// (4, 19, 'lutff_7/in_1')
// (4, 19, 'neigh_op_rgt_4')
// (4, 20, 'local_g1_4')
// (4, 20, 'lutff_0/in_1')
// (4, 20, 'lutff_1/in_0')
// (4, 20, 'lutff_3/in_0')
// (4, 20, 'lutff_6/in_3')
// (4, 20, 'neigh_op_bnr_4')
// (5, 18, 'local_g0_4')
// (5, 18, 'lutff_1/in_1')
// (5, 18, 'neigh_op_top_4')
// (5, 19, 'local_g2_4')
// (5, 19, 'local_g3_4')
// (5, 19, 'lutff_4/out')
// (5, 19, 'lutff_5/in_2')
// (5, 19, 'lutff_7/in_3')
// (5, 20, 'local_g1_4')
// (5, 20, 'lutff_0/in_1')
// (5, 20, 'lutff_3/in_0')
// (5, 20, 'lutff_6/in_3')
// (5, 20, 'neigh_op_bot_4')
// (6, 18, 'neigh_op_tnl_4')
// (6, 19, 'neigh_op_lft_4')
// (6, 20, 'neigh_op_bnl_4')

wire n786;
// (4, 18, 'neigh_op_tnr_6')
// (4, 19, 'local_g3_6')
// (4, 19, 'lutff_7/in_0')
// (4, 19, 'neigh_op_rgt_6')
// (4, 20, 'neigh_op_bnr_6')
// (5, 18, 'local_g1_6')
// (5, 18, 'lutff_0/in_3')
// (5, 18, 'neigh_op_top_6')
// (5, 19, 'local_g3_6')
// (5, 19, 'lutff_5/in_0')
// (5, 19, 'lutff_6/out')
// (5, 20, 'neigh_op_bot_6')
// (6, 18, 'neigh_op_tnl_6')
// (6, 19, 'neigh_op_lft_6')
// (6, 20, 'neigh_op_bnl_6')

wire n787;
// (4, 18, 'neigh_op_tnr_7')
// (4, 19, 'neigh_op_rgt_7')
// (4, 20, 'neigh_op_bnr_7')
// (5, 18, 'local_g1_7')
// (5, 18, 'lutff_6/in_2')
// (5, 18, 'neigh_op_top_7')
// (5, 19, 'lutff_7/out')
// (5, 20, 'neigh_op_bot_7')
// (6, 18, 'neigh_op_tnl_7')
// (6, 19, 'neigh_op_lft_7')
// (6, 20, 'neigh_op_bnl_7')

wire n788;
// (4, 19, 'lutff_0/cout')
// (4, 19, 'lutff_1/in_3')

wire n789;
// (4, 19, 'lutff_1/cout')
// (4, 19, 'lutff_2/in_3')

wire n790;
// (4, 19, 'lutff_3/cout')
// (4, 19, 'lutff_4/in_3')

wire n791;
// (4, 19, 'neigh_op_tnr_1')
// (4, 20, 'neigh_op_rgt_1')
// (4, 21, 'neigh_op_bnr_1')
// (5, 19, 'neigh_op_top_1')
// (5, 20, 'local_g1_1')
// (5, 20, 'lutff_0/in_2')
// (5, 20, 'lutff_1/out')
// (5, 21, 'neigh_op_bot_1')
// (6, 19, 'neigh_op_tnl_1')
// (6, 20, 'neigh_op_lft_1')
// (6, 21, 'neigh_op_bnl_1')

wire n792;
// (4, 19, 'neigh_op_tnr_2')
// (4, 20, 'neigh_op_rgt_2')
// (4, 21, 'neigh_op_bnr_2')
// (5, 19, 'neigh_op_top_2')
// (5, 20, 'local_g3_2')
// (5, 20, 'lutff_2/out')
// (5, 20, 'lutff_6/in_1')
// (5, 21, 'neigh_op_bot_2')
// (6, 19, 'neigh_op_tnl_2')
// (6, 20, 'neigh_op_lft_2')
// (6, 21, 'neigh_op_bnl_2')

wire n793;
// (4, 19, 'neigh_op_tnr_3')
// (4, 20, 'neigh_op_rgt_3')
// (4, 21, 'neigh_op_bnr_3')
// (5, 19, 'local_g0_3')
// (5, 19, 'lutff_2/in_1')
// (5, 19, 'neigh_op_top_3')
// (5, 20, 'lutff_3/out')
// (5, 21, 'neigh_op_bot_3')
// (6, 19, 'neigh_op_tnl_3')
// (6, 20, 'neigh_op_lft_3')
// (6, 21, 'neigh_op_bnl_3')

wire n794;
// (4, 19, 'neigh_op_tnr_4')
// (4, 20, 'neigh_op_rgt_4')
// (4, 21, 'neigh_op_bnr_4')
// (5, 19, 'neigh_op_top_4')
// (5, 20, 'local_g3_4')
// (5, 20, 'lutff_0/in_3')
// (5, 20, 'lutff_4/out')
// (5, 21, 'neigh_op_bot_4')
// (6, 19, 'neigh_op_tnl_4')
// (6, 20, 'neigh_op_lft_4')
// (6, 21, 'neigh_op_bnl_4')

wire n795;
// (4, 19, 'neigh_op_tnr_5')
// (4, 20, 'neigh_op_rgt_5')
// (4, 21, 'neigh_op_bnr_5')
// (5, 19, 'neigh_op_top_5')
// (5, 20, 'local_g1_5')
// (5, 20, 'lutff_5/out')
// (5, 20, 'lutff_6/in_0')
// (5, 21, 'neigh_op_bot_5')
// (6, 19, 'neigh_op_tnl_5')
// (6, 20, 'neigh_op_lft_5')
// (6, 21, 'neigh_op_bnl_5')

wire n796;
// (4, 19, 'neigh_op_tnr_7')
// (4, 20, 'neigh_op_rgt_7')
// (4, 21, 'neigh_op_bnr_7')
// (5, 19, 'neigh_op_top_7')
// (5, 20, 'local_g3_7')
// (5, 20, 'lutff_0/in_0')
// (5, 20, 'lutff_7/out')
// (5, 21, 'neigh_op_bot_7')
// (6, 19, 'neigh_op_tnl_7')
// (6, 20, 'neigh_op_lft_7')
// (6, 21, 'neigh_op_bnl_7')

wire n797;
// (4, 19, 'sp4_h_r_10')
// (5, 19, 'local_g1_7')
// (5, 19, 'lutff_3/in_1')
// (5, 19, 'sp4_h_r_23')
// (6, 19, 'sp4_h_r_34')
// (7, 19, 'sp4_h_r_47')
// (8, 18, 'neigh_op_tnr_1')
// (8, 19, 'neigh_op_rgt_1')
// (8, 19, 'sp4_h_l_47')
// (8, 19, 'sp4_h_r_7')
// (8, 20, 'local_g1_1')
// (8, 20, 'lutff_1/in_1')
// (8, 20, 'neigh_op_bnr_1')
// (9, 18, 'neigh_op_top_1')
// (9, 19, 'lutff_1/out')
// (9, 19, 'sp4_h_r_18')
// (9, 20, 'neigh_op_bot_1')
// (10, 18, 'neigh_op_tnl_1')
// (10, 19, 'neigh_op_lft_1')
// (10, 19, 'sp4_h_r_31')
// (10, 20, 'neigh_op_bnl_1')
// (11, 19, 'sp4_h_r_42')
// (12, 19, 'sp4_h_l_42')

wire n798;
// (4, 21, 'lutff_1/cout')
// (4, 21, 'lutff_2/in_3')

wire n799;
// (4, 21, 'lutff_2/cout')
// (4, 21, 'lutff_3/in_3')

wire n800;
// (4, 21, 'lutff_4/cout')
// (4, 21, 'lutff_5/in_3')

wire n801;
// (4, 21, 'lutff_5/cout')
// (4, 21, 'lutff_6/in_3')

wire n802;
// (4, 21, 'lutff_6/cout')
// (4, 21, 'lutff_7/in_3')

wire n803;
// (4, 21, 'lutff_7/cout')
// (4, 22, 'carry_in')
// (4, 22, 'carry_in_mux')
// (4, 22, 'lutff_0/in_3')

wire n804;
// (4, 22, 'lutff_0/cout')
// (4, 22, 'lutff_1/in_3')

wire n805;
// (5, 2, 'local_g0_0')
// (5, 2, 'lutff_5/in_1')
// (5, 2, 'sp4_h_r_0')
// (6, 1, 'neigh_op_tnr_4')
// (6, 2, 'neigh_op_rgt_4')
// (6, 2, 'sp4_h_r_13')
// (6, 3, 'neigh_op_bnr_4')
// (7, 1, 'neigh_op_top_4')
// (7, 2, 'lutff_4/out')
// (7, 2, 'sp4_h_r_24')
// (7, 3, 'neigh_op_bot_4')
// (8, 1, 'neigh_op_tnl_4')
// (8, 2, 'neigh_op_lft_4')
// (8, 2, 'sp4_h_r_37')
// (8, 3, 'neigh_op_bnl_4')
// (9, 2, 'sp4_h_l_37')

wire n806;
// (5, 2, 'sp4_h_r_2')
// (6, 2, 'sp4_h_r_15')
// (6, 3, 'sp4_r_v_b_40')
// (6, 4, 'sp4_r_v_b_29')
// (6, 5, 'sp4_r_v_b_16')
// (6, 6, 'sp4_r_v_b_5')
// (6, 7, 'sp4_r_v_b_43')
// (6, 8, 'sp4_r_v_b_30')
// (6, 9, 'sp4_r_v_b_19')
// (6, 10, 'sp4_r_v_b_6')
// (6, 11, 'sp4_r_v_b_39')
// (6, 12, 'sp4_r_v_b_26')
// (6, 13, 'sp4_r_v_b_15')
// (6, 14, 'sp4_r_v_b_2')
// (7, 2, 'local_g3_2')
// (7, 2, 'lutff_2/in_1')
// (7, 2, 'sp4_h_r_26')
// (7, 2, 'sp4_v_t_40')
// (7, 3, 'sp4_v_b_40')
// (7, 4, 'local_g2_5')
// (7, 4, 'lutff_5/in_0')
// (7, 4, 'lutff_7/in_0')
// (7, 4, 'sp4_v_b_29')
// (7, 5, 'sp4_v_b_16')
// (7, 6, 'sp4_h_r_0')
// (7, 6, 'sp4_v_b_5')
// (7, 6, 'sp4_v_t_43')
// (7, 7, 'sp4_v_b_43')
// (7, 8, 'sp4_v_b_30')
// (7, 9, 'sp4_v_b_19')
// (7, 10, 'sp4_v_b_6')
// (7, 10, 'sp4_v_t_39')
// (7, 11, 'sp4_v_b_39')
// (7, 12, 'sp4_v_b_26')
// (7, 13, 'local_g1_7')
// (7, 13, 'lutff_0/in_0')
// (7, 13, 'sp4_v_b_15')
// (7, 14, 'sp4_v_b_2')
// (8, 2, 'sp4_h_r_39')
// (8, 3, 'local_g3_5')
// (8, 3, 'lutff_4/in_2')
// (8, 3, 'sp4_r_v_b_45')
// (8, 4, 'sp4_r_v_b_32')
// (8, 5, 'local_g2_4')
// (8, 5, 'lutff_7/in_1')
// (8, 5, 'neigh_op_tnr_4')
// (8, 5, 'sp4_r_v_b_21')
// (8, 5, 'sp4_r_v_b_37')
// (8, 6, 'neigh_op_rgt_4')
// (8, 6, 'sp4_h_r_13')
// (8, 6, 'sp4_r_v_b_24')
// (8, 6, 'sp4_r_v_b_40')
// (8, 6, 'sp4_r_v_b_8')
// (8, 7, 'neigh_op_bnr_4')
// (8, 7, 'sp4_r_v_b_13')
// (8, 7, 'sp4_r_v_b_29')
// (8, 8, 'sp4_r_v_b_0')
// (8, 8, 'sp4_r_v_b_16')
// (8, 9, 'sp4_r_v_b_38')
// (8, 9, 'sp4_r_v_b_5')
// (8, 10, 'sp4_r_v_b_27')
// (8, 10, 'sp4_r_v_b_40')
// (8, 11, 'local_g2_6')
// (8, 11, 'lutff_6/in_0')
// (8, 11, 'sp4_r_v_b_14')
// (8, 11, 'sp4_r_v_b_29')
// (8, 12, 'sp4_r_v_b_16')
// (8, 12, 'sp4_r_v_b_3')
// (8, 13, 'sp4_r_v_b_5')
// (9, 2, 'sp4_h_l_39')
// (9, 2, 'sp4_v_t_45')
// (9, 3, 'sp4_v_b_45')
// (9, 4, 'local_g2_0')
// (9, 4, 'lutff_1/in_1')
// (9, 4, 'lutff_2/in_2')
// (9, 4, 'sp4_v_b_32')
// (9, 4, 'sp4_v_t_37')
// (9, 5, 'local_g0_4')
// (9, 5, 'lutff_2/in_0')
// (9, 5, 'lutff_4/in_0')
// (9, 5, 'neigh_op_top_4')
// (9, 5, 'sp4_r_v_b_36')
// (9, 5, 'sp4_v_b_21')
// (9, 5, 'sp4_v_b_37')
// (9, 5, 'sp4_v_t_40')
// (9, 6, 'lutff_4/out')
// (9, 6, 'sp4_h_r_24')
// (9, 6, 'sp4_r_v_b_25')
// (9, 6, 'sp4_v_b_24')
// (9, 6, 'sp4_v_b_40')
// (9, 6, 'sp4_v_b_8')
// (9, 7, 'neigh_op_bot_4')
// (9, 7, 'sp4_r_v_b_12')
// (9, 7, 'sp4_v_b_13')
// (9, 7, 'sp4_v_b_29')
// (9, 8, 'sp4_r_v_b_1')
// (9, 8, 'sp4_v_b_0')
// (9, 8, 'sp4_v_b_16')
// (9, 8, 'sp4_v_t_38')
// (9, 9, 'local_g1_5')
// (9, 9, 'lutff_0/in_0')
// (9, 9, 'sp4_r_v_b_36')
// (9, 9, 'sp4_v_b_38')
// (9, 9, 'sp4_v_b_5')
// (9, 9, 'sp4_v_t_40')
// (9, 10, 'sp4_r_v_b_25')
// (9, 10, 'sp4_v_b_27')
// (9, 10, 'sp4_v_b_40')
// (9, 11, 'sp4_r_v_b_12')
// (9, 11, 'sp4_v_b_14')
// (9, 11, 'sp4_v_b_29')
// (9, 12, 'local_g0_3')
// (9, 12, 'lutff_6/in_3')
// (9, 12, 'sp4_r_v_b_1')
// (9, 12, 'sp4_v_b_16')
// (9, 12, 'sp4_v_b_3')
// (9, 13, 'local_g1_5')
// (9, 13, 'lutff_1/in_1')
// (9, 13, 'lutff_3/in_3')
// (9, 13, 'lutff_4/in_2')
// (9, 13, 'sp4_v_b_5')
// (10, 4, 'sp4_v_t_36')
// (10, 5, 'neigh_op_tnl_4')
// (10, 5, 'sp4_v_b_36')
// (10, 6, 'neigh_op_lft_4')
// (10, 6, 'sp4_h_r_37')
// (10, 6, 'sp4_v_b_25')
// (10, 7, 'neigh_op_bnl_4')
// (10, 7, 'sp4_v_b_12')
// (10, 8, 'sp4_v_b_1')
// (10, 8, 'sp4_v_t_36')
// (10, 9, 'sp4_v_b_36')
// (10, 10, 'local_g3_1')
// (10, 10, 'lutff_6/in_0')
// (10, 10, 'sp4_v_b_25')
// (10, 11, 'sp4_v_b_12')
// (10, 12, 'sp4_v_b_1')
// (11, 6, 'sp4_h_l_37')

wire n807;
// (5, 5, 'sp12_h_r_1')
// (6, 5, 'sp12_h_r_2')
// (7, 5, 'sp12_h_r_5')
// (8, 5, 'local_g0_6')
// (8, 5, 'lutff_5/in_1')
// (8, 5, 'sp12_h_r_6')
// (9, 5, 'local_g0_1')
// (9, 5, 'lutff_1/in_2')
// (9, 5, 'sp12_h_r_9')
// (10, 5, 'sp12_h_r_10')
// (11, 2, 'sp4_r_v_b_42')
// (11, 3, 'sp4_r_v_b_31')
// (11, 4, 'sp4_r_v_b_18')
// (11, 5, 'sp12_h_r_13')
// (11, 5, 'sp4_r_v_b_7')
// (12, 1, 'sp4_v_t_42')
// (12, 2, 'sp4_v_b_42')
// (12, 3, 'local_g2_7')
// (12, 3, 'lutff_7/in_2')
// (12, 3, 'sp4_v_b_31')
// (12, 4, 'sp4_v_b_18')
// (12, 5, 'sp12_h_r_14')
// (12, 5, 'sp4_h_r_2')
// (12, 5, 'sp4_v_b_7')
// (13, 2, 'sp4_r_v_b_47')
// (13, 3, 'sp4_r_v_b_34')
// (13, 4, 'neigh_op_tnr_5')
// (13, 4, 'sp4_r_v_b_23')
// (13, 5, 'neigh_op_rgt_5')
// (13, 5, 'sp12_h_r_17')
// (13, 5, 'sp4_h_r_15')
// (13, 5, 'sp4_r_v_b_10')
// (13, 6, 'neigh_op_bnr_5')
// (14, 1, 'sp4_v_t_47')
// (14, 2, 'sp4_v_b_47')
// (14, 3, 'local_g3_2')
// (14, 3, 'lutff_7/in_2')
// (14, 3, 'sp4_v_b_34')
// (14, 4, 'neigh_op_top_5')
// (14, 4, 'sp4_v_b_23')
// (14, 5, 'lutff_5/out')
// (14, 5, 'sp12_h_r_18')
// (14, 5, 'sp4_h_r_26')
// (14, 5, 'sp4_v_b_10')
// (14, 6, 'neigh_op_bot_5')
// (15, 4, 'neigh_op_tnl_5')
// (15, 5, 'neigh_op_lft_5')
// (15, 5, 'sp12_h_r_21')
// (15, 5, 'sp4_h_r_39')
// (15, 6, 'neigh_op_bnl_5')
// (16, 5, 'sp12_h_r_22')
// (16, 5, 'sp4_h_l_39')
// (17, 5, 'sp12_h_l_22')

wire n808;
// (5, 5, 'sp4_h_r_9')
// (6, 5, 'sp4_h_r_20')
// (7, 4, 'neigh_op_tnr_6')
// (7, 5, 'local_g2_1')
// (7, 5, 'lutff_1/in_0')
// (7, 5, 'neigh_op_rgt_6')
// (7, 5, 'sp4_h_r_33')
// (7, 6, 'neigh_op_bnr_6')
// (8, 4, 'neigh_op_top_6')
// (8, 5, 'lutff_6/out')
// (8, 5, 'sp4_h_r_44')
// (8, 6, 'neigh_op_bot_6')
// (9, 4, 'neigh_op_tnl_6')
// (9, 5, 'neigh_op_lft_6')
// (9, 5, 'sp4_h_l_44')
// (9, 6, 'neigh_op_bnl_6')

wire n809;
// (5, 6, 'lutff_1/cout')
// (5, 6, 'lutff_2/in_3')

reg n810 = 0;
// (5, 6, 'sp4_r_v_b_38')
// (5, 7, 'sp4_r_v_b_27')
// (5, 8, 'sp4_r_v_b_14')
// (5, 9, 'local_g1_3')
// (5, 9, 'lutff_4/in_2')
// (5, 9, 'sp4_r_v_b_3')
// (6, 4, 'neigh_op_tnr_2')
// (6, 5, 'neigh_op_rgt_2')
// (6, 5, 'sp4_h_r_9')
// (6, 5, 'sp4_v_t_38')
// (6, 6, 'neigh_op_bnr_2')
// (6, 6, 'sp4_v_b_38')
// (6, 7, 'sp4_v_b_27')
// (6, 8, 'sp4_v_b_14')
// (6, 9, 'sp4_v_b_3')
// (7, 4, 'neigh_op_top_2')
// (7, 5, 'lutff_2/out')
// (7, 5, 'sp4_h_r_20')
// (7, 6, 'neigh_op_bot_2')
// (8, 4, 'neigh_op_tnl_2')
// (8, 5, 'neigh_op_lft_2')
// (8, 5, 'sp4_h_r_33')
// (8, 6, 'neigh_op_bnl_2')
// (9, 5, 'sp4_h_r_44')
// (10, 5, 'sp4_h_l_44')

wire n811;
// (5, 8, 'local_g1_2')
// (5, 8, 'lutff_2/in_3')
// (5, 8, 'sp4_h_r_2')
// (5, 8, 'sp4_r_v_b_42')
// (5, 9, 'local_g0_7')
// (5, 9, 'lutff_2/in_3')
// (5, 9, 'lutff_5/in_0')
// (5, 9, 'sp4_r_v_b_31')
// (5, 10, 'local_g3_2')
// (5, 10, 'lutff_2/in_3')
// (5, 10, 'lutff_3/in_0')
// (5, 10, 'lutff_7/in_0')
// (5, 10, 'sp4_r_v_b_18')
// (5, 11, 'sp4_r_v_b_7')
// (6, 7, 'sp4_h_r_1')
// (6, 7, 'sp4_v_t_42')
// (6, 8, 'sp4_h_r_15')
// (6, 8, 'sp4_v_b_42')
// (6, 9, 'sp4_v_b_31')
// (6, 10, 'sp4_h_r_0')
// (6, 10, 'sp4_v_b_18')
// (6, 11, 'sp4_v_b_7')
// (7, 7, 'sp4_h_r_12')
// (7, 8, 'sp4_h_r_26')
// (7, 8, 'sp4_r_v_b_38')
// (7, 9, 'sp4_r_v_b_27')
// (7, 10, 'local_g1_5')
// (7, 10, 'lutff_1/in_1')
// (7, 10, 'sp4_h_r_13')
// (7, 10, 'sp4_r_v_b_14')
// (7, 11, 'local_g1_3')
// (7, 11, 'lutff_2/in_2')
// (7, 11, 'sp4_r_v_b_3')
// (8, 5, 'sp4_r_v_b_44')
// (8, 6, 'neigh_op_tnr_2')
// (8, 6, 'sp4_r_v_b_33')
// (8, 7, 'neigh_op_rgt_2')
// (8, 7, 'sp4_h_r_25')
// (8, 7, 'sp4_h_r_9')
// (8, 7, 'sp4_r_v_b_20')
// (8, 7, 'sp4_r_v_b_36')
// (8, 7, 'sp4_v_t_38')
// (8, 8, 'neigh_op_bnr_2')
// (8, 8, 'sp4_h_r_39')
// (8, 8, 'sp4_r_v_b_25')
// (8, 8, 'sp4_r_v_b_9')
// (8, 8, 'sp4_v_b_38')
// (8, 9, 'sp4_r_v_b_12')
// (8, 9, 'sp4_v_b_27')
// (8, 10, 'local_g1_1')
// (8, 10, 'lutff_7/in_3')
// (8, 10, 'sp4_h_r_24')
// (8, 10, 'sp4_r_v_b_1')
// (8, 10, 'sp4_v_b_14')
// (8, 11, 'local_g0_3')
// (8, 11, 'lutff_1/in_2')
// (8, 11, 'sp4_v_b_3')
// (9, 4, 'sp4_v_t_44')
// (9, 5, 'sp12_v_t_23')
// (9, 5, 'sp4_v_b_44')
// (9, 6, 'neigh_op_top_2')
// (9, 6, 'sp12_v_b_23')
// (9, 6, 'sp4_v_b_33')
// (9, 6, 'sp4_v_t_36')
// (9, 7, 'local_g3_2')
// (9, 7, 'lutff_0/in_1')
// (9, 7, 'lutff_2/out')
// (9, 7, 'sp12_v_b_20')
// (9, 7, 'sp4_h_r_20')
// (9, 7, 'sp4_h_r_36')
// (9, 7, 'sp4_r_v_b_37')
// (9, 7, 'sp4_v_b_20')
// (9, 7, 'sp4_v_b_36')
// (9, 8, 'local_g1_2')
// (9, 8, 'lutff_0/in_3')
// (9, 8, 'lutff_1/in_0')
// (9, 8, 'lutff_3/in_2')
// (9, 8, 'lutff_6/in_1')
// (9, 8, 'neigh_op_bot_2')
// (9, 8, 'sp12_v_b_19')
// (9, 8, 'sp4_h_l_39')
// (9, 8, 'sp4_r_v_b_24')
// (9, 8, 'sp4_v_b_25')
// (9, 8, 'sp4_v_b_9')
// (9, 9, 'local_g0_4')
// (9, 9, 'lutff_1/in_3')
// (9, 9, 'lutff_3/in_3')
// (9, 9, 'lutff_6/in_2')
// (9, 9, 'sp12_v_b_16')
// (9, 9, 'sp4_r_v_b_13')
// (9, 9, 'sp4_v_b_12')
// (9, 10, 'local_g1_0')
// (9, 10, 'lutff_0/in_3')
// (9, 10, 'lutff_5/in_0')
// (9, 10, 'sp12_v_b_15')
// (9, 10, 'sp4_h_r_37')
// (9, 10, 'sp4_r_v_b_0')
// (9, 10, 'sp4_v_b_1')
// (9, 11, 'local_g3_4')
// (9, 11, 'lutff_1/in_0')
// (9, 11, 'sp12_v_b_12')
// (9, 12, 'sp12_v_b_11')
// (9, 13, 'sp12_v_b_8')
// (9, 14, 'sp12_v_b_7')
// (9, 15, 'sp12_v_b_4')
// (9, 16, 'sp12_v_b_3')
// (9, 17, 'sp12_v_b_0')
// (10, 6, 'neigh_op_tnl_2')
// (10, 6, 'sp4_v_t_37')
// (10, 7, 'local_g0_2')
// (10, 7, 'lutff_0/in_2')
// (10, 7, 'neigh_op_lft_2')
// (10, 7, 'sp4_h_l_36')
// (10, 7, 'sp4_h_r_33')
// (10, 7, 'sp4_v_b_37')
// (10, 8, 'local_g3_2')
// (10, 8, 'lutff_2/in_1')
// (10, 8, 'neigh_op_bnl_2')
// (10, 8, 'sp4_v_b_24')
// (10, 9, 'local_g0_5')
// (10, 9, 'lutff_4/in_3')
// (10, 9, 'lutff_5/in_2')
// (10, 9, 'lutff_6/in_1')
// (10, 9, 'sp4_v_b_13')
// (10, 10, 'local_g1_0')
// (10, 10, 'lutff_1/in_2')
// (10, 10, 'lutff_2/in_3')
// (10, 10, 'sp4_h_l_37')
// (10, 10, 'sp4_v_b_0')
// (11, 7, 'sp4_h_r_44')
// (12, 7, 'sp4_h_l_44')

reg n812 = 0;
// (5, 8, 'sp4_h_r_1')
// (6, 8, 'sp4_h_r_12')
// (7, 7, 'local_g3_2')
// (7, 7, 'lutff_4/in_3')
// (7, 7, 'neigh_op_tnr_2')
// (7, 8, 'neigh_op_rgt_2')
// (7, 8, 'sp4_h_r_25')
// (7, 8, 'sp4_h_r_9')
// (7, 9, 'local_g1_2')
// (7, 9, 'lutff_6/in_1')
// (7, 9, 'neigh_op_bnr_2')
// (8, 7, 'local_g0_2')
// (8, 7, 'lutff_0/in_2')
// (8, 7, 'neigh_op_top_2')
// (8, 8, 'lutff_2/out')
// (8, 8, 'sp4_h_r_20')
// (8, 8, 'sp4_h_r_36')
// (8, 9, 'local_g0_2')
// (8, 9, 'local_g1_2')
// (8, 9, 'lutff_0/in_1')
// (8, 9, 'lutff_1/in_3')
// (8, 9, 'neigh_op_bot_2')
// (9, 7, 'neigh_op_tnl_2')
// (9, 8, 'neigh_op_lft_2')
// (9, 8, 'sp4_h_l_36')
// (9, 8, 'sp4_h_r_33')
// (9, 8, 'sp4_h_r_4')
// (9, 9, 'neigh_op_bnl_2')
// (10, 8, 'local_g1_1')
// (10, 8, 'lutff_2/in_2')
// (10, 8, 'sp4_h_r_17')
// (10, 8, 'sp4_h_r_44')
// (10, 9, 'sp4_r_v_b_44')
// (10, 10, 'local_g0_2')
// (10, 10, 'lutff_1/in_3')
// (10, 10, 'sp4_r_v_b_33')
// (10, 11, 'sp4_r_v_b_20')
// (10, 12, 'sp4_r_v_b_9')
// (11, 8, 'sp4_h_l_44')
// (11, 8, 'sp4_h_r_28')
// (11, 8, 'sp4_v_t_44')
// (11, 9, 'sp4_v_b_44')
// (11, 10, 'sp4_v_b_33')
// (11, 11, 'sp4_v_b_20')
// (11, 12, 'sp4_v_b_9')
// (12, 8, 'sp4_h_r_41')
// (13, 8, 'sp4_h_l_41')

wire n813;
// (5, 11, 'lutff_1/cout')
// (5, 11, 'lutff_2/in_3')

wire n814;
// (5, 11, 'lutff_2/cout')
// (5, 11, 'lutff_3/in_3')

wire n815;
// (5, 11, 'lutff_3/cout')
// (5, 11, 'lutff_4/in_3')

wire n816;
// (5, 11, 'sp4_r_v_b_37')
// (5, 12, 'sp4_r_v_b_24')
// (5, 13, 'sp4_r_v_b_13')
// (5, 14, 'local_g1_0')
// (5, 14, 'lutff_7/in_0')
// (5, 14, 'sp4_r_v_b_0')
// (6, 10, 'sp4_h_r_6')
// (6, 10, 'sp4_v_t_37')
// (6, 11, 'sp4_v_b_37')
// (6, 12, 'sp4_v_b_24')
// (6, 13, 'sp4_v_b_13')
// (6, 14, 'sp4_h_r_4')
// (6, 14, 'sp4_v_b_0')
// (7, 3, 'sp4_r_v_b_36')
// (7, 4, 'sp4_r_v_b_25')
// (7, 5, 'sp4_r_v_b_12')
// (7, 6, 'sp4_r_v_b_1')
// (7, 10, 'sp4_h_r_19')
// (7, 14, 'local_g1_1')
// (7, 14, 'lutff_1/in_1')
// (7, 14, 'sp4_h_r_17')
// (8, 2, 'sp4_v_t_36')
// (8, 3, 'sp4_v_b_36')
// (8, 4, 'sp4_v_b_25')
// (8, 5, 'local_g0_4')
// (8, 5, 'lutff_2/in_2')
// (8, 5, 'sp4_v_b_12')
// (8, 6, 'local_g1_0')
// (8, 6, 'lutff_1/in_2')
// (8, 6, 'lutff_7/in_0')
// (8, 6, 'sp4_h_r_8')
// (8, 6, 'sp4_v_b_1')
// (8, 10, 'sp4_h_r_30')
// (8, 14, 'sp4_h_r_28')
// (9, 6, 'sp4_h_r_21')
// (9, 10, 'sp4_h_r_43')
// (9, 11, 'sp4_r_v_b_41')
// (9, 12, 'sp4_r_v_b_28')
// (9, 13, 'sp4_r_v_b_17')
// (9, 14, 'sp4_h_r_41')
// (9, 14, 'sp4_r_v_b_4')
// (10, 6, 'sp4_h_r_32')
// (10, 10, 'sp4_h_l_43')
// (10, 10, 'sp4_h_r_10')
// (10, 10, 'sp4_v_t_41')
// (10, 11, 'sp4_v_b_41')
// (10, 12, 'sp4_v_b_28')
// (10, 13, 'sp4_v_b_17')
// (10, 14, 'sp4_h_l_41')
// (10, 14, 'sp4_v_b_4')
// (11, 4, 'sp4_r_v_b_42')
// (11, 5, 'local_g1_7')
// (11, 5, 'lutff_6/in_0')
// (11, 5, 'sp4_r_v_b_31')
// (11, 6, 'sp4_h_r_45')
// (11, 6, 'sp4_r_v_b_18')
// (11, 7, 'local_g2_7')
// (11, 7, 'lutff_1/in_2')
// (11, 7, 'sp4_r_v_b_39')
// (11, 7, 'sp4_r_v_b_7')
// (11, 8, 'sp4_r_v_b_26')
// (11, 8, 'sp4_r_v_b_42')
// (11, 9, 'neigh_op_tnr_1')
// (11, 9, 'sp4_r_v_b_15')
// (11, 9, 'sp4_r_v_b_31')
// (11, 10, 'neigh_op_rgt_1')
// (11, 10, 'sp4_h_r_23')
// (11, 10, 'sp4_r_v_b_18')
// (11, 10, 'sp4_r_v_b_2')
// (11, 11, 'local_g1_1')
// (11, 11, 'lutff_6/in_2')
// (11, 11, 'neigh_op_bnr_1')
// (11, 11, 'sp4_r_v_b_7')
// (12, 3, 'sp4_r_v_b_43')
// (12, 3, 'sp4_v_t_42')
// (12, 4, 'sp4_r_v_b_30')
// (12, 4, 'sp4_v_b_42')
// (12, 5, 'local_g3_3')
// (12, 5, 'lutff_7/in_1')
// (12, 5, 'sp4_r_v_b_19')
// (12, 5, 'sp4_v_b_31')
// (12, 6, 'local_g0_2')
// (12, 6, 'lutff_7/in_1')
// (12, 6, 'sp4_h_l_45')
// (12, 6, 'sp4_r_v_b_6')
// (12, 6, 'sp4_v_b_18')
// (12, 6, 'sp4_v_t_39')
// (12, 7, 'sp4_r_v_b_38')
// (12, 7, 'sp4_v_b_39')
// (12, 7, 'sp4_v_b_7')
// (12, 7, 'sp4_v_t_42')
// (12, 8, 'sp4_r_v_b_27')
// (12, 8, 'sp4_v_b_26')
// (12, 8, 'sp4_v_b_42')
// (12, 9, 'neigh_op_top_1')
// (12, 9, 'sp4_r_v_b_14')
// (12, 9, 'sp4_v_b_15')
// (12, 9, 'sp4_v_b_31')
// (12, 10, 'lutff_1/out')
// (12, 10, 'sp4_h_r_34')
// (12, 10, 'sp4_r_v_b_3')
// (12, 10, 'sp4_v_b_18')
// (12, 10, 'sp4_v_b_2')
// (12, 11, 'neigh_op_bot_1')
// (12, 11, 'sp4_v_b_7')
// (13, 2, 'sp4_v_t_43')
// (13, 3, 'local_g3_3')
// (13, 3, 'lutff_5/in_1')
// (13, 3, 'sp4_v_b_43')
// (13, 4, 'sp4_v_b_30')
// (13, 5, 'sp4_v_b_19')
// (13, 6, 'sp4_v_b_6')
// (13, 6, 'sp4_v_t_38')
// (13, 7, 'sp4_v_b_38')
// (13, 8, 'sp4_v_b_27')
// (13, 9, 'neigh_op_tnl_1')
// (13, 9, 'sp4_v_b_14')
// (13, 10, 'neigh_op_lft_1')
// (13, 10, 'sp4_h_r_47')
// (13, 10, 'sp4_v_b_3')
// (13, 11, 'neigh_op_bnl_1')
// (14, 10, 'sp4_h_l_47')

wire n817;
// (5, 12, 'local_g1_7')
// (5, 12, 'lutff_3/in_3')
// (5, 12, 'sp4_h_r_7')
// (6, 12, 'sp4_h_r_18')
// (7, 12, 'sp4_h_r_31')
// (8, 12, 'sp4_h_r_42')
// (9, 12, 'local_g1_3')
// (9, 12, 'lutff_0/in_2')
// (9, 12, 'lutff_1/in_3')
// (9, 12, 'sp4_h_l_42')
// (9, 12, 'sp4_h_r_11')
// (10, 12, 'sp4_h_r_22')
// (11, 11, 'neigh_op_tnr_7')
// (11, 12, 'neigh_op_rgt_7')
// (11, 12, 'sp4_h_r_35')
// (11, 13, 'neigh_op_bnr_7')
// (12, 11, 'neigh_op_top_7')
// (12, 12, 'local_g2_7')
// (12, 12, 'lutff_6/in_3')
// (12, 12, 'lutff_7/out')
// (12, 12, 'sp4_h_r_46')
// (12, 13, 'neigh_op_bot_7')
// (13, 11, 'neigh_op_tnl_7')
// (13, 12, 'neigh_op_lft_7')
// (13, 12, 'sp4_h_l_46')
// (13, 13, 'neigh_op_bnl_7')

wire n818;
// (5, 14, 'sp4_h_r_8')
// (6, 9, 'sp4_r_v_b_46')
// (6, 10, 'sp4_r_v_b_35')
// (6, 11, 'sp4_r_v_b_22')
// (6, 12, 'sp4_r_v_b_11')
// (6, 13, 'neigh_op_tnr_0')
// (6, 13, 'sp4_r_v_b_45')
// (6, 14, 'neigh_op_rgt_0')
// (6, 14, 'sp4_h_r_21')
// (6, 14, 'sp4_r_v_b_32')
// (6, 15, 'neigh_op_bnr_0')
// (6, 15, 'sp4_r_v_b_21')
// (6, 16, 'sp4_r_v_b_8')
// (7, 8, 'sp4_v_t_46')
// (7, 9, 'sp4_v_b_46')
// (7, 10, 'sp4_v_b_35')
// (7, 11, 'sp4_v_b_22')
// (7, 12, 'local_g1_3')
// (7, 12, 'lutff_global/cen')
// (7, 12, 'sp4_v_b_11')
// (7, 12, 'sp4_v_t_45')
// (7, 13, 'neigh_op_top_0')
// (7, 13, 'sp4_v_b_45')
// (7, 14, 'local_g1_0')
// (7, 14, 'lutff_0/out')
// (7, 14, 'lutff_2/in_1')
// (7, 14, 'sp4_h_r_32')
// (7, 14, 'sp4_v_b_32')
// (7, 15, 'neigh_op_bot_0')
// (7, 15, 'sp4_v_b_21')
// (7, 16, 'sp4_v_b_8')
// (8, 11, 'sp4_r_v_b_39')
// (8, 12, 'sp4_r_v_b_26')
// (8, 13, 'neigh_op_tnl_0')
// (8, 13, 'sp4_r_v_b_15')
// (8, 14, 'neigh_op_lft_0')
// (8, 14, 'sp4_h_r_45')
// (8, 14, 'sp4_r_v_b_2')
// (8, 15, 'neigh_op_bnl_0')
// (9, 10, 'sp4_v_t_39')
// (9, 11, 'sp4_v_b_39')
// (9, 12, 'local_g2_2')
// (9, 12, 'lutff_global/cen')
// (9, 12, 'sp4_v_b_26')
// (9, 13, 'sp4_v_b_15')
// (9, 14, 'sp4_h_l_45')
// (9, 14, 'sp4_v_b_2')

reg n819 = 0;
// (5, 14, 'sp4_r_v_b_45')
// (5, 15, 'local_g2_0')
// (5, 15, 'lutff_3/in_1')
// (5, 15, 'sp4_r_v_b_32')
// (5, 16, 'sp4_r_v_b_21')
// (5, 17, 'sp4_r_v_b_8')
// (6, 13, 'sp4_h_r_2')
// (6, 13, 'sp4_v_t_45')
// (6, 14, 'sp4_v_b_45')
// (6, 15, 'sp4_v_b_32')
// (6, 16, 'sp4_v_b_21')
// (6, 17, 'sp4_v_b_8')
// (7, 13, 'sp4_h_r_15')
// (8, 13, 'sp4_h_r_26')
// (9, 13, 'sp4_h_r_39')
// (10, 12, 'neigh_op_tnr_3')
// (10, 13, 'neigh_op_rgt_3')
// (10, 13, 'sp4_h_l_39')
// (10, 13, 'sp4_h_r_11')
// (10, 14, 'local_g0_3')
// (10, 14, 'lutff_0/in_1')
// (10, 14, 'neigh_op_bnr_3')
// (11, 12, 'neigh_op_top_3')
// (11, 13, 'lutff_3/out')
// (11, 13, 'sp4_h_r_22')
// (11, 14, 'neigh_op_bot_3')
// (12, 12, 'neigh_op_tnl_3')
// (12, 13, 'neigh_op_lft_3')
// (12, 13, 'sp4_h_r_35')
// (12, 14, 'neigh_op_bnl_3')
// (13, 13, 'sp4_h_r_46')
// (14, 13, 'sp4_h_l_46')

wire n820;
// (5, 15, 'sp4_h_r_0')
// (6, 15, 'sp4_h_r_13')
// (6, 18, 'sp4_r_v_b_37')
// (6, 19, 'sp4_r_v_b_24')
// (6, 20, 'sp4_r_v_b_13')
// (6, 21, 'sp4_r_v_b_0')
// (7, 15, 'local_g3_0')
// (7, 15, 'lutff_7/in_2')
// (7, 15, 'sp4_h_r_24')
// (7, 17, 'sp4_h_r_6')
// (7, 17, 'sp4_v_t_37')
// (7, 18, 'sp4_v_b_37')
// (7, 19, 'sp4_v_b_24')
// (7, 20, 'local_g1_5')
// (7, 20, 'lutff_7/in_1')
// (7, 20, 'sp4_v_b_13')
// (7, 21, 'sp4_v_b_0')
// (8, 15, 'sp4_h_r_37')
// (8, 16, 'neigh_op_tnr_7')
// (8, 16, 'sp4_r_v_b_43')
// (8, 17, 'neigh_op_rgt_7')
// (8, 17, 'sp4_h_r_19')
// (8, 17, 'sp4_r_v_b_30')
// (8, 18, 'neigh_op_bnr_7')
// (8, 18, 'sp4_r_v_b_19')
// (8, 19, 'local_g1_6')
// (8, 19, 'lutff_7/in_2')
// (8, 19, 'sp4_r_v_b_6')
// (9, 15, 'sp4_h_l_37')
// (9, 15, 'sp4_v_t_43')
// (9, 16, 'local_g1_7')
// (9, 16, 'lutff_7/in_1')
// (9, 16, 'neigh_op_top_7')
// (9, 16, 'sp4_v_b_43')
// (9, 17, 'lutff_7/out')
// (9, 17, 'sp4_h_r_30')
// (9, 17, 'sp4_v_b_30')
// (9, 18, 'neigh_op_bot_7')
// (9, 18, 'sp4_v_b_19')
// (9, 19, 'sp4_v_b_6')
// (10, 16, 'neigh_op_tnl_7')
// (10, 17, 'neigh_op_lft_7')
// (10, 17, 'sp4_h_r_43')
// (10, 18, 'neigh_op_bnl_7')
// (11, 17, 'sp4_h_l_43')

wire n821;
// (5, 16, 'sp4_h_r_6')
// (6, 15, 'neigh_op_tnr_7')
// (6, 16, 'neigh_op_rgt_7')
// (6, 16, 'sp4_h_r_19')
// (6, 17, 'neigh_op_bnr_7')
// (7, 15, 'neigh_op_top_7')
// (7, 15, 'sp4_r_v_b_42')
// (7, 16, 'lutff_7/out')
// (7, 16, 'sp4_h_r_30')
// (7, 16, 'sp4_r_v_b_31')
// (7, 17, 'neigh_op_bot_7')
// (7, 17, 'sp4_r_v_b_18')
// (7, 18, 'local_g1_7')
// (7, 18, 'lutff_7/in_1')
// (7, 18, 'sp4_r_v_b_7')
// (8, 14, 'sp4_v_t_42')
// (8, 15, 'local_g3_2')
// (8, 15, 'lutff_7/in_2')
// (8, 15, 'neigh_op_tnl_7')
// (8, 15, 'sp4_v_b_42')
// (8, 16, 'neigh_op_lft_7')
// (8, 16, 'sp4_h_r_43')
// (8, 16, 'sp4_v_b_31')
// (8, 17, 'local_g2_7')
// (8, 17, 'lutff_7/in_2')
// (8, 17, 'neigh_op_bnl_7')
// (8, 17, 'sp4_r_v_b_43')
// (8, 17, 'sp4_v_b_18')
// (8, 18, 'sp4_r_v_b_30')
// (8, 18, 'sp4_v_b_7')
// (8, 19, 'sp4_r_v_b_19')
// (8, 20, 'sp4_r_v_b_6')
// (9, 16, 'sp4_h_l_43')
// (9, 16, 'sp4_v_t_43')
// (9, 17, 'sp4_v_b_43')
// (9, 18, 'local_g3_6')
// (9, 18, 'lutff_7/in_2')
// (9, 18, 'sp4_v_b_30')
// (9, 19, 'sp4_v_b_19')
// (9, 20, 'sp4_v_b_6')

wire n822;
// (5, 19, 'local_g0_2')
// (5, 19, 'lutff_1/in_3')
// (5, 19, 'sp4_h_r_10')
// (6, 18, 'neigh_op_tnr_1')
// (6, 19, 'neigh_op_rgt_1')
// (6, 19, 'sp4_h_r_23')
// (6, 20, 'neigh_op_bnr_1')
// (7, 18, 'neigh_op_top_1')
// (7, 19, 'lutff_1/out')
// (7, 19, 'sp4_h_r_34')
// (7, 20, 'neigh_op_bot_1')
// (8, 18, 'neigh_op_tnl_1')
// (8, 19, 'neigh_op_lft_1')
// (8, 19, 'sp4_h_r_47')
// (8, 20, 'neigh_op_bnl_1')
// (9, 19, 'sp4_h_l_47')

wire n823;
// (6, 0, 'logic_op_tnr_1')
// (6, 1, 'neigh_op_rgt_1')
// (6, 2, 'neigh_op_bnr_1')
// (7, 0, 'logic_op_top_1')
// (7, 1, 'lutff_1/out')
// (7, 2, 'neigh_op_bot_1')
// (8, 0, 'logic_op_tnl_1')
// (8, 1, 'neigh_op_lft_1')
// (8, 2, 'local_g3_1')
// (8, 2, 'lutff_2/in_2')
// (8, 2, 'neigh_op_bnl_1')

wire n824;
// (6, 0, 'logic_op_tnr_2')
// (6, 1, 'neigh_op_rgt_2')
// (6, 2, 'neigh_op_bnr_2')
// (7, 0, 'logic_op_top_2')
// (7, 1, 'lutff_2/out')
// (7, 2, 'local_g1_2')
// (7, 2, 'lutff_0/in_3')
// (7, 2, 'neigh_op_bot_2')
// (8, 0, 'logic_op_tnl_2')
// (8, 1, 'neigh_op_lft_2')
// (8, 2, 'neigh_op_bnl_2')

reg n825 = 0;
// (6, 0, 'logic_op_tnr_3')
// (6, 1, 'neigh_op_rgt_3')
// (6, 2, 'neigh_op_bnr_3')
// (7, 0, 'logic_op_top_3')
// (7, 1, 'local_g1_3')
// (7, 1, 'lutff_3/out')
// (7, 1, 'lutff_5/in_1')
// (7, 2, 'neigh_op_bot_3')
// (8, 0, 'logic_op_tnl_3')
// (8, 1, 'local_g0_3')
// (8, 1, 'lutff_1/in_0')
// (8, 1, 'neigh_op_lft_3')
// (8, 2, 'neigh_op_bnl_3')

wire n826;
// (6, 0, 'logic_op_tnr_5')
// (6, 1, 'neigh_op_rgt_5')
// (6, 2, 'neigh_op_bnr_5')
// (7, 0, 'logic_op_top_5')
// (7, 1, 'lutff_5/out')
// (7, 1, 'sp4_r_v_b_43')
// (7, 2, 'neigh_op_bot_5')
// (7, 2, 'sp4_r_v_b_30')
// (7, 3, 'sp4_r_v_b_19')
// (7, 4, 'sp4_r_v_b_6')
// (8, 0, 'logic_op_tnl_5')
// (8, 0, 'span4_vert_43')
// (8, 1, 'neigh_op_lft_5')
// (8, 1, 'sp4_v_b_43')
// (8, 2, 'neigh_op_bnl_5')
// (8, 2, 'sp4_v_b_30')
// (8, 3, 'local_g1_3')
// (8, 3, 'lutff_4/in_0')
// (8, 3, 'sp4_v_b_19')
// (8, 4, 'sp4_v_b_6')

wire n827;
// (6, 0, 'logic_op_tnr_6')
// (6, 1, 'neigh_op_rgt_6')
// (6, 1, 'sp4_r_v_b_44')
// (6, 2, 'neigh_op_bnr_6')
// (6, 2, 'sp4_r_v_b_33')
// (6, 3, 'sp4_r_v_b_20')
// (6, 4, 'sp4_r_v_b_9')
// (7, 0, 'logic_op_top_6')
// (7, 0, 'span4_vert_44')
// (7, 1, 'lutff_6/out')
// (7, 1, 'sp4_v_b_44')
// (7, 2, 'neigh_op_bot_6')
// (7, 2, 'sp4_v_b_33')
// (7, 3, 'sp4_v_b_20')
// (7, 4, 'local_g0_1')
// (7, 4, 'lutff_7/in_2')
// (7, 4, 'sp4_v_b_9')
// (8, 0, 'logic_op_tnl_6')
// (8, 1, 'neigh_op_lft_6')
// (8, 2, 'neigh_op_bnl_6')

wire n828;
// (6, 0, 'logic_op_tnr_7')
// (6, 1, 'neigh_op_rgt_7')
// (6, 2, 'neigh_op_bnr_7')
// (7, 0, 'logic_op_top_7')
// (7, 1, 'lutff_7/out')
// (7, 2, 'neigh_op_bot_7')
// (8, 0, 'logic_op_tnl_7')
// (8, 1, 'local_g0_7')
// (8, 1, 'lutff_3/in_2')
// (8, 1, 'neigh_op_lft_7')
// (8, 2, 'neigh_op_bnl_7')

wire n829;
// (6, 1, 'neigh_op_tnr_0')
// (6, 2, 'neigh_op_rgt_0')
// (6, 3, 'neigh_op_bnr_0')
// (7, 1, 'neigh_op_top_0')
// (7, 2, 'local_g1_0')
// (7, 2, 'lutff_0/out')
// (7, 2, 'lutff_6/in_1')
// (7, 3, 'neigh_op_bot_0')
// (8, 1, 'neigh_op_tnl_0')
// (8, 2, 'neigh_op_lft_0')
// (8, 3, 'neigh_op_bnl_0')

wire n830;
// (6, 1, 'neigh_op_tnr_1')
// (6, 2, 'neigh_op_rgt_1')
// (6, 3, 'neigh_op_bnr_1')
// (7, 1, 'neigh_op_top_1')
// (7, 2, 'lutff_1/out')
// (7, 3, 'local_g1_1')
// (7, 3, 'lutff_4/in_0')
// (7, 3, 'neigh_op_bot_1')
// (8, 1, 'neigh_op_tnl_1')
// (8, 2, 'neigh_op_lft_1')
// (8, 3, 'neigh_op_bnl_1')

wire n831;
// (6, 1, 'neigh_op_tnr_2')
// (6, 2, 'neigh_op_rgt_2')
// (6, 2, 'sp4_r_v_b_36')
// (6, 3, 'neigh_op_bnr_2')
// (6, 3, 'sp4_r_v_b_25')
// (6, 4, 'sp4_r_v_b_12')
// (6, 5, 'sp4_r_v_b_1')
// (7, 1, 'neigh_op_top_2')
// (7, 1, 'sp4_v_t_36')
// (7, 2, 'lutff_2/out')
// (7, 2, 'sp4_v_b_36')
// (7, 3, 'neigh_op_bot_2')
// (7, 3, 'sp4_v_b_25')
// (7, 4, 'local_g1_4')
// (7, 4, 'lutff_6/in_1')
// (7, 4, 'sp4_v_b_12')
// (7, 5, 'sp4_v_b_1')
// (8, 1, 'neigh_op_tnl_2')
// (8, 2, 'neigh_op_lft_2')
// (8, 3, 'neigh_op_bnl_2')

wire n832;
// (6, 1, 'neigh_op_tnr_5')
// (6, 2, 'neigh_op_rgt_5')
// (6, 3, 'neigh_op_bnr_5')
// (7, 1, 'neigh_op_top_5')
// (7, 2, 'local_g3_5')
// (7, 2, 'lutff_5/out')
// (7, 2, 'lutff_6/in_0')
// (7, 3, 'neigh_op_bot_5')
// (8, 1, 'neigh_op_tnl_5')
// (8, 2, 'neigh_op_lft_5')
// (8, 3, 'neigh_op_bnl_5')

wire n833;
// (6, 1, 'neigh_op_tnr_6')
// (6, 2, 'neigh_op_rgt_6')
// (6, 3, 'neigh_op_bnr_6')
// (7, 1, 'neigh_op_top_6')
// (7, 2, 'lutff_6/out')
// (7, 3, 'local_g1_6')
// (7, 3, 'lutff_4/in_1')
// (7, 3, 'neigh_op_bot_6')
// (8, 1, 'neigh_op_tnl_6')
// (8, 2, 'neigh_op_lft_6')
// (8, 3, 'neigh_op_bnl_6')

reg n834 = 0;
// (6, 1, 'sp4_r_v_b_24')
// (6, 2, 'neigh_op_tnr_0')
// (6, 2, 'sp4_r_v_b_13')
// (6, 3, 'neigh_op_rgt_0')
// (6, 3, 'sp4_r_v_b_0')
// (6, 4, 'neigh_op_bnr_0')
// (7, 0, 'span4_vert_24')
// (7, 1, 'local_g3_0')
// (7, 1, 'lutff_6/in_1')
// (7, 1, 'sp4_r_v_b_25')
// (7, 1, 'sp4_v_b_24')
// (7, 2, 'neigh_op_top_0')
// (7, 2, 'sp4_r_v_b_12')
// (7, 2, 'sp4_v_b_13')
// (7, 3, 'lutff_0/out')
// (7, 3, 'sp4_r_v_b_1')
// (7, 3, 'sp4_v_b_0')
// (7, 4, 'neigh_op_bot_0')
// (8, 0, 'span4_vert_25')
// (8, 1, 'local_g3_1')
// (8, 1, 'lutff_1/in_3')
// (8, 1, 'sp4_v_b_25')
// (8, 2, 'neigh_op_tnl_0')
// (8, 2, 'sp4_v_b_12')
// (8, 3, 'neigh_op_lft_0')
// (8, 3, 'sp4_v_b_1')
// (8, 4, 'neigh_op_bnl_0')

reg n835 = 0;
// (6, 1, 'sp4_r_v_b_28')
// (6, 2, 'neigh_op_tnr_2')
// (6, 2, 'sp4_r_v_b_17')
// (6, 3, 'neigh_op_rgt_2')
// (6, 3, 'sp4_r_v_b_4')
// (6, 4, 'neigh_op_bnr_2')
// (7, 0, 'span4_vert_28')
// (7, 1, 'local_g3_4')
// (7, 1, 'lutff_1/in_0')
// (7, 1, 'sp4_v_b_28')
// (7, 2, 'neigh_op_top_2')
// (7, 2, 'sp4_v_b_17')
// (7, 3, 'local_g3_2')
// (7, 3, 'lutff_2/out')
// (7, 3, 'lutff_7/in_0')
// (7, 3, 'sp4_v_b_4')
// (7, 4, 'neigh_op_bot_2')
// (8, 2, 'neigh_op_tnl_2')
// (8, 3, 'neigh_op_lft_2')
// (8, 4, 'neigh_op_bnl_2')

reg n836 = 0;
// (6, 1, 'sp4_r_v_b_34')
// (6, 2, 'neigh_op_tnr_5')
// (6, 2, 'sp4_r_v_b_23')
// (6, 3, 'neigh_op_rgt_5')
// (6, 3, 'sp4_r_v_b_10')
// (6, 4, 'neigh_op_bnr_5')
// (7, 0, 'span4_vert_34')
// (7, 1, 'local_g3_2')
// (7, 1, 'lutff_1/in_2')
// (7, 1, 'sp4_v_b_34')
// (7, 2, 'neigh_op_top_5')
// (7, 2, 'sp4_v_b_23')
// (7, 3, 'lutff_5/out')
// (7, 3, 'sp4_v_b_10')
// (7, 4, 'neigh_op_bot_5')
// (8, 2, 'neigh_op_tnl_5')
// (8, 3, 'local_g0_5')
// (8, 3, 'lutff_2/in_1')
// (8, 3, 'neigh_op_lft_5')
// (8, 4, 'neigh_op_bnl_5')

wire n837;
// (6, 2, 'neigh_op_tnr_1')
// (6, 3, 'neigh_op_rgt_1')
// (6, 4, 'neigh_op_bnr_1')
// (7, 2, 'local_g1_1')
// (7, 2, 'lutff_2/in_2')
// (7, 2, 'neigh_op_top_1')
// (7, 3, 'lutff_1/out')
// (7, 4, 'neigh_op_bot_1')
// (8, 2, 'neigh_op_tnl_1')
// (8, 3, 'neigh_op_lft_1')
// (8, 4, 'neigh_op_bnl_1')

wire n838;
// (6, 2, 'neigh_op_tnr_6')
// (6, 3, 'neigh_op_rgt_6')
// (6, 4, 'neigh_op_bnr_6')
// (7, 2, 'local_g1_6')
// (7, 2, 'lutff_1/in_0')
// (7, 2, 'neigh_op_top_6')
// (7, 3, 'lutff_6/out')
// (7, 4, 'neigh_op_bot_6')
// (8, 2, 'neigh_op_tnl_6')
// (8, 3, 'neigh_op_lft_6')
// (8, 4, 'neigh_op_bnl_6')

wire n839;
// (6, 2, 'neigh_op_tnr_7')
// (6, 3, 'neigh_op_rgt_7')
// (6, 4, 'neigh_op_bnr_7')
// (7, 2, 'local_g1_7')
// (7, 2, 'lutff_2/in_0')
// (7, 2, 'neigh_op_top_7')
// (7, 3, 'lutff_7/out')
// (7, 4, 'neigh_op_bot_7')
// (8, 2, 'neigh_op_tnl_7')
// (8, 3, 'neigh_op_lft_7')
// (8, 4, 'neigh_op_bnl_7')

wire n840;
// (6, 2, 'sp4_h_r_3')
// (6, 3, 'sp4_h_r_10')
// (7, 2, 'sp4_h_r_14')
// (7, 3, 'sp4_h_r_23')
// (8, 2, 'local_g3_3')
// (8, 2, 'lutff_global/cen')
// (8, 2, 'sp4_h_r_27')
// (8, 2, 'sp4_r_v_b_42')
// (8, 3, 'local_g2_2')
// (8, 3, 'lutff_global/cen')
// (8, 3, 'sp4_h_r_34')
// (8, 3, 'sp4_r_v_b_31')
// (8, 4, 'sp4_r_v_b_18')
// (8, 5, 'sp4_r_v_b_7')
// (9, 1, 'sp4_v_t_42')
// (9, 2, 'sp4_h_r_38')
// (9, 2, 'sp4_v_b_42')
// (9, 3, 'sp4_h_r_47')
// (9, 3, 'sp4_v_b_31')
// (9, 4, 'local_g0_2')
// (9, 4, 'lutff_global/cen')
// (9, 4, 'sp4_v_b_18')
// (9, 5, 'local_g0_2')
// (9, 5, 'lutff_global/cen')
// (9, 5, 'sp4_h_r_2')
// (9, 5, 'sp4_v_b_7')
// (10, 2, 'sp4_h_l_38')
// (10, 2, 'sp4_h_r_0')
// (10, 3, 'sp4_h_l_47')
// (10, 3, 'sp4_h_r_7')
// (10, 5, 'sp4_h_r_15')
// (11, 2, 'sp4_h_r_13')
// (11, 3, 'sp4_h_r_18')
// (11, 5, 'sp4_h_r_26')
// (12, 2, 'neigh_op_tnr_5')
// (12, 2, 'sp4_h_r_24')
// (12, 2, 'sp4_r_v_b_39')
// (12, 3, 'neigh_op_rgt_5')
// (12, 3, 'sp4_h_r_31')
// (12, 3, 'sp4_r_v_b_26')
// (12, 4, 'neigh_op_bnr_5')
// (12, 4, 'sp4_r_v_b_15')
// (12, 5, 'sp4_h_r_39')
// (12, 5, 'sp4_r_v_b_2')
// (13, 1, 'sp4_v_t_39')
// (13, 2, 'neigh_op_top_5')
// (13, 2, 'sp4_h_r_37')
// (13, 2, 'sp4_v_b_39')
// (13, 3, 'lutff_5/out')
// (13, 3, 'sp4_h_r_42')
// (13, 3, 'sp4_r_v_b_43')
// (13, 3, 'sp4_v_b_26')
// (13, 4, 'neigh_op_bot_5')
// (13, 4, 'sp4_r_v_b_30')
// (13, 4, 'sp4_v_b_15')
// (13, 5, 'sp4_h_l_39')
// (13, 5, 'sp4_r_v_b_19')
// (13, 5, 'sp4_v_b_2')
// (13, 6, 'sp4_r_v_b_6')
// (14, 2, 'neigh_op_tnl_5')
// (14, 2, 'sp4_h_l_37')
// (14, 2, 'sp4_v_t_43')
// (14, 3, 'neigh_op_lft_5')
// (14, 3, 'sp4_h_l_42')
// (14, 3, 'sp4_v_b_43')
// (14, 4, 'neigh_op_bnl_5')
// (14, 4, 'sp4_v_b_30')
// (14, 5, 'sp4_v_b_19')
// (14, 6, 'sp4_v_b_6')

wire n841;
// (6, 2, 'sp4_h_r_5')
// (6, 3, 'sp4_h_r_8')
// (7, 2, 'sp4_h_r_16')
// (7, 2, 'sp4_r_v_b_45')
// (7, 3, 'local_g0_5')
// (7, 3, 'lutff_1/in_2')
// (7, 3, 'sp4_h_r_21')
// (7, 3, 'sp4_r_v_b_32')
// (7, 4, 'sp4_r_v_b_21')
// (7, 5, 'sp4_r_v_b_8')
// (7, 6, 'sp4_h_r_4')
// (8, 1, 'sp4_v_t_45')
// (8, 2, 'local_g2_5')
// (8, 2, 'lutff_7/in_0')
// (8, 2, 'sp4_h_r_29')
// (8, 2, 'sp4_v_b_45')
// (8, 3, 'local_g3_0')
// (8, 3, 'lutff_7/in_0')
// (8, 3, 'sp4_h_r_32')
// (8, 3, 'sp4_v_b_32')
// (8, 4, 'local_g1_5')
// (8, 4, 'lutff_1/in_1')
// (8, 4, 'sp4_v_b_21')
// (8, 5, 'sp4_h_r_8')
// (8, 5, 'sp4_v_b_8')
// (8, 6, 'local_g0_1')
// (8, 6, 'lutff_7/in_2')
// (8, 6, 'sp4_h_r_17')
// (9, 2, 'sp4_h_r_40')
// (9, 2, 'sp4_r_v_b_37')
// (9, 3, 'local_g1_0')
// (9, 3, 'lutff_7/in_0')
// (9, 3, 'sp4_h_r_45')
// (9, 3, 'sp4_r_v_b_24')
// (9, 3, 'sp4_r_v_b_40')
// (9, 4, 'local_g3_0')
// (9, 4, 'lutff_3/in_2')
// (9, 4, 'neigh_op_tnr_0')
// (9, 4, 'sp4_r_v_b_13')
// (9, 4, 'sp4_r_v_b_29')
// (9, 4, 'sp4_r_v_b_45')
// (9, 5, 'local_g2_0')
// (9, 5, 'local_g3_0')
// (9, 5, 'lutff_0/in_0')
// (9, 5, 'lutff_5/in_2')
// (9, 5, 'lutff_7/in_2')
// (9, 5, 'neigh_op_rgt_0')
// (9, 5, 'sp4_h_r_21')
// (9, 5, 'sp4_r_v_b_0')
// (9, 5, 'sp4_r_v_b_16')
// (9, 5, 'sp4_r_v_b_32')
// (9, 6, 'neigh_op_bnr_0')
// (9, 6, 'sp4_h_r_28')
// (9, 6, 'sp4_r_v_b_21')
// (9, 6, 'sp4_r_v_b_5')
// (9, 7, 'sp4_r_v_b_8')
// (10, 1, 'sp4_v_t_37')
// (10, 2, 'sp4_h_l_40')
// (10, 2, 'sp4_v_b_37')
// (10, 2, 'sp4_v_t_40')
// (10, 3, 'sp4_h_l_45')
// (10, 3, 'sp4_r_v_b_41')
// (10, 3, 'sp4_v_b_24')
// (10, 3, 'sp4_v_b_40')
// (10, 3, 'sp4_v_t_45')
// (10, 4, 'local_g2_5')
// (10, 4, 'lutff_6/in_1')
// (10, 4, 'neigh_op_top_0')
// (10, 4, 'sp4_r_v_b_28')
// (10, 4, 'sp4_r_v_b_44')
// (10, 4, 'sp4_v_b_13')
// (10, 4, 'sp4_v_b_29')
// (10, 4, 'sp4_v_b_45')
// (10, 5, 'lutff_0/out')
// (10, 5, 'sp4_h_r_0')
// (10, 5, 'sp4_h_r_32')
// (10, 5, 'sp4_r_v_b_17')
// (10, 5, 'sp4_r_v_b_33')
// (10, 5, 'sp4_v_b_0')
// (10, 5, 'sp4_v_b_16')
// (10, 5, 'sp4_v_b_32')
// (10, 6, 'neigh_op_bot_0')
// (10, 6, 'sp4_h_r_41')
// (10, 6, 'sp4_r_v_b_20')
// (10, 6, 'sp4_r_v_b_4')
// (10, 6, 'sp4_v_b_21')
// (10, 6, 'sp4_v_b_5')
// (10, 7, 'local_g1_0')
// (10, 7, 'lutff_2/in_3')
// (10, 7, 'sp4_r_v_b_9')
// (10, 7, 'sp4_v_b_8')
// (11, 2, 'sp4_v_t_41')
// (11, 3, 'sp4_v_b_41')
// (11, 3, 'sp4_v_t_44')
// (11, 4, 'neigh_op_tnl_0')
// (11, 4, 'sp4_v_b_28')
// (11, 4, 'sp4_v_b_44')
// (11, 5, 'neigh_op_lft_0')
// (11, 5, 'sp4_h_r_13')
// (11, 5, 'sp4_h_r_45')
// (11, 5, 'sp4_v_b_17')
// (11, 5, 'sp4_v_b_33')
// (11, 6, 'neigh_op_bnl_0')
// (11, 6, 'sp4_h_l_41')
// (11, 6, 'sp4_h_r_4')
// (11, 6, 'sp4_v_b_20')
// (11, 6, 'sp4_v_b_4')
// (11, 7, 'local_g1_1')
// (11, 7, 'lutff_0/in_2')
// (11, 7, 'lutff_1/in_1')
// (11, 7, 'lutff_2/in_0')
// (11, 7, 'lutff_3/in_1')
// (11, 7, 'lutff_7/in_1')
// (11, 7, 'sp4_h_r_3')
// (11, 7, 'sp4_v_b_9')
// (12, 5, 'local_g3_0')
// (12, 5, 'lutff_2/in_1')
// (12, 5, 'sp4_h_l_45')
// (12, 5, 'sp4_h_r_24')
// (12, 6, 'local_g0_1')
// (12, 6, 'lutff_0/in_1')
// (12, 6, 'sp4_h_r_17')
// (12, 7, 'sp4_h_r_14')
// (13, 5, 'local_g2_5')
// (13, 5, 'lutff_0/in_1')
// (13, 5, 'sp4_h_r_37')
// (13, 6, 'sp4_h_r_28')
// (13, 7, 'local_g2_3')
// (13, 7, 'lutff_1/in_0')
// (13, 7, 'sp4_h_r_27')
// (14, 5, 'sp4_h_l_37')
// (14, 6, 'sp4_h_r_41')
// (14, 7, 'sp4_h_r_38')
// (15, 6, 'sp4_h_l_41')
// (15, 7, 'sp4_h_l_38')

wire n842;
// (6, 2, 'sp4_r_v_b_44')
// (6, 3, 'neigh_op_tnr_2')
// (6, 3, 'sp4_r_v_b_33')
// (6, 4, 'neigh_op_rgt_2')
// (6, 4, 'sp4_r_v_b_20')
// (6, 5, 'neigh_op_bnr_2')
// (6, 5, 'sp4_r_v_b_9')
// (7, 1, 'sp4_v_t_44')
// (7, 2, 'sp4_v_b_44')
// (7, 3, 'neigh_op_top_2')
// (7, 3, 'sp4_v_b_33')
// (7, 4, 'lutff_2/out')
// (7, 4, 'sp4_v_b_20')
// (7, 5, 'local_g0_1')
// (7, 5, 'lutff_2/in_1')
// (7, 5, 'neigh_op_bot_2')
// (7, 5, 'sp4_v_b_9')
// (8, 3, 'neigh_op_tnl_2')
// (8, 4, 'neigh_op_lft_2')
// (8, 5, 'neigh_op_bnl_2')

wire n843;
// (6, 3, 'neigh_op_tnr_1')
// (6, 4, 'neigh_op_rgt_1')
// (6, 5, 'neigh_op_bnr_1')
// (7, 3, 'neigh_op_top_1')
// (7, 4, 'lutff_1/out')
// (7, 5, 'local_g1_1')
// (7, 5, 'lutff_3/in_3')
// (7, 5, 'neigh_op_bot_1')
// (8, 3, 'neigh_op_tnl_1')
// (8, 4, 'neigh_op_lft_1')
// (8, 5, 'neigh_op_bnl_1')

wire n844;
// (6, 3, 'neigh_op_tnr_3')
// (6, 4, 'neigh_op_rgt_3')
// (6, 5, 'neigh_op_bnr_3')
// (7, 3, 'neigh_op_top_3')
// (7, 4, 'lutff_3/out')
// (7, 5, 'local_g1_3')
// (7, 5, 'lutff_4/in_0')
// (7, 5, 'neigh_op_bot_3')
// (8, 3, 'neigh_op_tnl_3')
// (8, 4, 'neigh_op_lft_3')
// (8, 5, 'neigh_op_bnl_3')

wire n845;
// (6, 3, 'neigh_op_tnr_5')
// (6, 4, 'neigh_op_rgt_5')
// (6, 5, 'neigh_op_bnr_5')
// (7, 3, 'neigh_op_top_5')
// (7, 4, 'lutff_5/out')
// (7, 5, 'local_g1_5')
// (7, 5, 'lutff_0/in_0')
// (7, 5, 'neigh_op_bot_5')
// (8, 3, 'neigh_op_tnl_5')
// (8, 4, 'neigh_op_lft_5')
// (8, 5, 'neigh_op_bnl_5')

wire n846;
// (6, 3, 'neigh_op_tnr_6')
// (6, 4, 'neigh_op_rgt_6')
// (6, 5, 'neigh_op_bnr_6')
// (7, 3, 'neigh_op_top_6')
// (7, 4, 'lutff_6/out')
// (7, 5, 'local_g0_6')
// (7, 5, 'lutff_6/in_2')
// (7, 5, 'neigh_op_bot_6')
// (8, 3, 'neigh_op_tnl_6')
// (8, 4, 'neigh_op_lft_6')
// (8, 5, 'neigh_op_bnl_6')

wire n847;
// (6, 3, 'neigh_op_tnr_7')
// (6, 4, 'neigh_op_rgt_7')
// (6, 5, 'neigh_op_bnr_7')
// (7, 3, 'neigh_op_top_7')
// (7, 4, 'local_g1_7')
// (7, 4, 'lutff_1/in_3')
// (7, 4, 'lutff_7/out')
// (7, 5, 'neigh_op_bot_7')
// (8, 3, 'neigh_op_tnl_7')
// (8, 4, 'neigh_op_lft_7')
// (8, 5, 'neigh_op_bnl_7')

wire n848;
// (6, 4, 'neigh_op_tnr_1')
// (6, 5, 'neigh_op_rgt_1')
// (6, 6, 'neigh_op_bnr_1')
// (7, 4, 'neigh_op_top_1')
// (7, 5, 'lutff_1/out')
// (7, 6, 'local_g0_1')
// (7, 6, 'lutff_7/in_0')
// (7, 6, 'neigh_op_bot_1')
// (8, 4, 'neigh_op_tnl_1')
// (8, 5, 'neigh_op_lft_1')
// (8, 6, 'neigh_op_bnl_1')

reg n849 = 0;
// (6, 4, 'neigh_op_tnr_3')
// (6, 5, 'neigh_op_rgt_3')
// (6, 5, 'sp4_r_v_b_38')
// (6, 6, 'neigh_op_bnr_3')
// (6, 6, 'sp4_r_v_b_27')
// (6, 7, 'sp4_r_v_b_14')
// (6, 8, 'sp4_r_v_b_3')
// (7, 4, 'neigh_op_top_3')
// (7, 4, 'sp4_v_t_38')
// (7, 5, 'lutff_3/out')
// (7, 5, 'sp4_v_b_38')
// (7, 6, 'neigh_op_bot_3')
// (7, 6, 'sp4_v_b_27')
// (7, 7, 'local_g1_6')
// (7, 7, 'lutff_5/in_2')
// (7, 7, 'sp4_v_b_14')
// (7, 8, 'sp4_v_b_3')
// (8, 4, 'neigh_op_tnl_3')
// (8, 5, 'neigh_op_lft_3')
// (8, 6, 'neigh_op_bnl_3')

wire n850;
// (6, 4, 'neigh_op_tnr_5')
// (6, 5, 'neigh_op_rgt_5')
// (6, 6, 'neigh_op_bnr_5')
// (7, 4, 'neigh_op_top_5')
// (7, 5, 'lutff_5/out')
// (7, 6, 'local_g0_5')
// (7, 6, 'lutff_4/in_1')
// (7, 6, 'neigh_op_bot_5')
// (8, 4, 'neigh_op_tnl_5')
// (8, 5, 'neigh_op_lft_5')
// (8, 6, 'neigh_op_bnl_5')

wire n851;
// (6, 4, 'sp4_h_r_1')
// (6, 4, 'sp4_h_r_5')
// (7, 1, 'sp4_h_r_11')
// (7, 4, 'sp4_h_r_12')
// (7, 4, 'sp4_h_r_16')
// (8, 1, 'sp4_h_r_22')
// (8, 4, 'sp4_h_r_25')
// (8, 4, 'sp4_h_r_29')
// (9, 1, 'local_g3_3')
// (9, 1, 'lutff_global/cen')
// (9, 1, 'sp4_h_r_35')
// (9, 1, 'sp4_r_v_b_42')
// (9, 1, 'sp4_r_v_b_43')
// (9, 2, 'sp4_r_v_b_30')
// (9, 2, 'sp4_r_v_b_31')
// (9, 3, 'local_g3_3')
// (9, 3, 'lutff_global/cen')
// (9, 3, 'sp4_r_v_b_18')
// (9, 3, 'sp4_r_v_b_19')
// (9, 4, 'sp4_h_r_36')
// (9, 4, 'sp4_h_r_40')
// (9, 4, 'sp4_r_v_b_6')
// (9, 4, 'sp4_r_v_b_7')
// (10, 0, 'span4_vert_42')
// (10, 0, 'span4_vert_43')
// (10, 1, 'sp4_h_r_46')
// (10, 1, 'sp4_v_b_42')
// (10, 1, 'sp4_v_b_43')
// (10, 2, 'sp4_r_v_b_40')
// (10, 2, 'sp4_v_b_30')
// (10, 2, 'sp4_v_b_31')
// (10, 3, 'local_g0_2')
// (10, 3, 'lutff_global/cen')
// (10, 3, 'neigh_op_tnr_0')
// (10, 3, 'sp4_r_v_b_29')
// (10, 3, 'sp4_v_b_18')
// (10, 3, 'sp4_v_b_19')
// (10, 4, 'neigh_op_rgt_0')
// (10, 4, 'sp4_h_l_36')
// (10, 4, 'sp4_h_l_40')
// (10, 4, 'sp4_h_r_1')
// (10, 4, 'sp4_h_r_5')
// (10, 4, 'sp4_r_v_b_16')
// (10, 4, 'sp4_v_b_6')
// (10, 4, 'sp4_v_b_7')
// (10, 5, 'neigh_op_bnr_0')
// (10, 5, 'sp4_r_v_b_5')
// (11, 1, 'sp4_h_l_46')
// (11, 1, 'sp4_v_t_40')
// (11, 2, 'sp4_v_b_40')
// (11, 3, 'neigh_op_top_0')
// (11, 3, 'sp4_v_b_29')
// (11, 4, 'lutff_0/out')
// (11, 4, 'sp4_h_r_12')
// (11, 4, 'sp4_h_r_16')
// (11, 4, 'sp4_v_b_16')
// (11, 5, 'neigh_op_bot_0')
// (11, 5, 'sp4_v_b_5')
// (12, 3, 'neigh_op_tnl_0')
// (12, 4, 'neigh_op_lft_0')
// (12, 4, 'sp4_h_r_25')
// (12, 4, 'sp4_h_r_29')
// (12, 5, 'neigh_op_bnl_0')
// (13, 4, 'sp4_h_r_36')
// (13, 4, 'sp4_h_r_40')
// (14, 4, 'sp4_h_l_36')
// (14, 4, 'sp4_h_l_40')

reg n852 = 0;
// (6, 4, 'sp4_r_v_b_42')
// (6, 5, 'sp4_r_v_b_31')
// (6, 6, 'sp4_r_v_b_18')
// (6, 7, 'sp4_r_v_b_7')
// (7, 3, 'sp4_h_r_7')
// (7, 3, 'sp4_v_t_42')
// (7, 4, 'sp4_v_b_42')
// (7, 5, 'sp4_v_b_31')
// (7, 6, 'local_g1_2')
// (7, 6, 'lutff_5/in_0')
// (7, 6, 'sp4_v_b_18')
// (7, 7, 'sp4_v_b_7')
// (8, 3, 'sp4_h_r_18')
// (8, 4, 'sp4_r_v_b_40')
// (8, 4, 'sp4_r_v_b_46')
// (8, 5, 'local_g2_3')
// (8, 5, 'lutff_2/in_1')
// (8, 5, 'sp4_r_v_b_29')
// (8, 5, 'sp4_r_v_b_35')
// (8, 6, 'local_g3_6')
// (8, 6, 'lutff_0/in_1')
// (8, 6, 'lutff_4/in_1')
// (8, 6, 'lutff_6/in_1')
// (8, 6, 'sp4_r_v_b_16')
// (8, 6, 'sp4_r_v_b_22')
// (8, 7, 'sp4_r_v_b_11')
// (8, 7, 'sp4_r_v_b_5')
// (8, 8, 'sp4_r_v_b_39')
// (8, 9, 'sp4_r_v_b_26')
// (8, 10, 'local_g2_7')
// (8, 10, 'lutff_2/in_3')
// (8, 10, 'sp4_r_v_b_15')
// (8, 11, 'sp4_r_v_b_2')
// (9, 3, 'sp4_h_r_31')
// (9, 3, 'sp4_h_r_5')
// (9, 3, 'sp4_v_t_40')
// (9, 3, 'sp4_v_t_46')
// (9, 4, 'sp4_v_b_40')
// (9, 4, 'sp4_v_b_46')
// (9, 5, 'local_g2_3')
// (9, 5, 'lutff_1/in_0')
// (9, 5, 'sp4_v_b_29')
// (9, 5, 'sp4_v_b_35')
// (9, 6, 'local_g1_6')
// (9, 6, 'lutff_4/in_1')
// (9, 6, 'sp4_v_b_16')
// (9, 6, 'sp4_v_b_22')
// (9, 7, 'local_g0_5')
// (9, 7, 'local_g1_3')
// (9, 7, 'lutff_2/in_2')
// (9, 7, 'lutff_7/in_2')
// (9, 7, 'sp4_v_b_11')
// (9, 7, 'sp4_v_b_5')
// (9, 7, 'sp4_v_t_39')
// (9, 8, 'sp4_v_b_39')
// (9, 9, 'sp4_v_b_26')
// (9, 10, 'sp4_v_b_15')
// (9, 11, 'sp4_v_b_2')
// (10, 3, 'sp4_h_r_16')
// (10, 3, 'sp4_h_r_42')
// (10, 4, 'sp4_h_r_2')
// (10, 4, 'sp4_r_v_b_41')
// (10, 4, 'sp4_r_v_b_47')
// (10, 5, 'local_g1_4')
// (10, 5, 'lutff_0/in_3')
// (10, 5, 'sp4_r_v_b_28')
// (10, 5, 'sp4_r_v_b_34')
// (10, 6, 'local_g3_1')
// (10, 6, 'lutff_2/in_0')
// (10, 6, 'lutff_3/in_3')
// (10, 6, 'lutff_5/in_3')
// (10, 6, 'sp4_r_v_b_17')
// (10, 6, 'sp4_r_v_b_23')
// (10, 7, 'sp4_r_v_b_10')
// (10, 7, 'sp4_r_v_b_4')
// (10, 8, 'sp4_r_v_b_42')
// (10, 8, 'sp4_r_v_b_47')
// (10, 9, 'sp4_r_v_b_31')
// (10, 9, 'sp4_r_v_b_34')
// (10, 10, 'sp4_r_v_b_18')
// (10, 10, 'sp4_r_v_b_23')
// (10, 11, 'sp4_r_v_b_10')
// (10, 11, 'sp4_r_v_b_7')
// (11, 3, 'local_g1_4')
// (11, 3, 'lutff_0/in_1')
// (11, 3, 'lutff_3/in_2')
// (11, 3, 'sp4_h_l_42')
// (11, 3, 'sp4_h_r_29')
// (11, 3, 'sp4_h_r_4')
// (11, 3, 'sp4_v_t_41')
// (11, 3, 'sp4_v_t_47')
// (11, 4, 'local_g0_7')
// (11, 4, 'lutff_2/in_3')
// (11, 4, 'sp4_h_r_1')
// (11, 4, 'sp4_h_r_15')
// (11, 4, 'sp4_v_b_41')
// (11, 4, 'sp4_v_b_47')
// (11, 5, 'sp4_v_b_28')
// (11, 5, 'sp4_v_b_34')
// (11, 6, 'local_g1_7')
// (11, 6, 'lutff_4/in_0')
// (11, 6, 'sp4_v_b_17')
// (11, 6, 'sp4_v_b_23')
// (11, 7, 'local_g0_2')
// (11, 7, 'lutff_6/in_0')
// (11, 7, 'sp4_v_b_10')
// (11, 7, 'sp4_v_b_4')
// (11, 7, 'sp4_v_t_42')
// (11, 7, 'sp4_v_t_47')
// (11, 8, 'sp4_v_b_42')
// (11, 8, 'sp4_v_b_47')
// (11, 9, 'sp4_v_b_31')
// (11, 9, 'sp4_v_b_34')
// (11, 10, 'local_g0_2')
// (11, 10, 'lutff_2/in_2')
// (11, 10, 'lutff_4/in_0')
// (11, 10, 'sp4_v_b_18')
// (11, 10, 'sp4_v_b_23')
// (11, 11, 'local_g1_2')
// (11, 11, 'lutff_7/in_2')
// (11, 11, 'sp4_v_b_10')
// (11, 11, 'sp4_v_b_7')
// (12, 1, 'sp4_r_v_b_33')
// (12, 2, 'local_g3_4')
// (12, 2, 'lutff_2/in_3')
// (12, 2, 'sp4_r_v_b_20')
// (12, 3, 'sp4_h_r_17')
// (12, 3, 'sp4_h_r_40')
// (12, 3, 'sp4_r_v_b_9')
// (12, 4, 'local_g0_4')
// (12, 4, 'lutff_0/in_2')
// (12, 4, 'lutff_1/in_1')
// (12, 4, 'lutff_2/in_2')
// (12, 4, 'sp4_h_r_12')
// (12, 4, 'sp4_h_r_26')
// (12, 4, 'sp4_r_v_b_44')
// (12, 5, 'local_g0_2')
// (12, 5, 'lutff_7/in_3')
// (12, 5, 'sp4_r_v_b_33')
// (12, 6, 'sp4_r_v_b_20')
// (12, 7, 'sp4_r_v_b_9')
// (13, 0, 'span4_vert_33')
// (13, 1, 'sp4_r_v_b_39')
// (13, 1, 'sp4_v_b_33')
// (13, 2, 'sp4_r_v_b_26')
// (13, 2, 'sp4_v_b_20')
// (13, 3, 'sp4_h_l_40')
// (13, 3, 'sp4_h_r_28')
// (13, 3, 'sp4_h_r_9')
// (13, 3, 'sp4_r_v_b_15')
// (13, 3, 'sp4_v_b_9')
// (13, 3, 'sp4_v_t_44')
// (13, 4, 'local_g1_2')
// (13, 4, 'lutff_2/in_3')
// (13, 4, 'sp4_h_r_25')
// (13, 4, 'sp4_h_r_39')
// (13, 4, 'sp4_r_v_b_2')
// (13, 4, 'sp4_v_b_44')
// (13, 5, 'sp4_v_b_33')
// (13, 6, 'sp4_v_b_20')
// (13, 7, 'sp4_v_b_9')
// (13, 13, 'sp4_r_v_b_39')
// (13, 14, 'sp4_r_v_b_26')
// (13, 15, 'sp4_r_v_b_15')
// (13, 16, 'local_g1_2')
// (13, 16, 'lutff_3/in_0')
// (13, 16, 'lutff_5/in_0')
// (13, 16, 'sp4_r_v_b_2')
// (14, 0, 'span4_vert_39')
// (14, 1, 'sp4_r_v_b_25')
// (14, 1, 'sp4_r_v_b_30')
// (14, 1, 'sp4_v_b_39')
// (14, 2, 'local_g2_4')
// (14, 2, 'lutff_0/in_0')
// (14, 2, 'lutff_2/in_2')
// (14, 2, 'sp4_r_v_b_12')
// (14, 2, 'sp4_r_v_b_19')
// (14, 2, 'sp4_v_b_26')
// (14, 3, 'local_g1_6')
// (14, 3, 'lutff_7/in_0')
// (14, 3, 'sp4_h_r_20')
// (14, 3, 'sp4_h_r_41')
// (14, 3, 'sp4_r_v_b_1')
// (14, 3, 'sp4_r_v_b_6')
// (14, 3, 'sp4_v_b_15')
// (14, 4, 'local_g2_4')
// (14, 4, 'lutff_0/in_2')
// (14, 4, 'sp4_h_l_39')
// (14, 4, 'sp4_h_r_2')
// (14, 4, 'sp4_h_r_36')
// (14, 4, 'sp4_r_v_b_36')
// (14, 4, 'sp4_v_b_2')
// (14, 5, 'sp4_r_v_b_25')
// (14, 6, 'sp4_r_v_b_12')
// (14, 7, 'sp4_r_v_b_1')
// (14, 12, 'sp4_h_r_8')
// (14, 12, 'sp4_v_t_39')
// (14, 13, 'sp4_v_b_39')
// (14, 14, 'sp4_v_b_26')
// (14, 15, 'sp4_v_b_15')
// (14, 16, 'sp4_v_b_2')
// (15, 0, 'span4_vert_25')
// (15, 0, 'span4_vert_30')
// (15, 1, 'sp4_v_b_25')
// (15, 1, 'sp4_v_b_30')
// (15, 2, 'sp4_v_b_12')
// (15, 2, 'sp4_v_b_19')
// (15, 3, 'sp4_h_l_41')
// (15, 3, 'sp4_h_r_1')
// (15, 3, 'sp4_h_r_33')
// (15, 3, 'sp4_v_b_1')
// (15, 3, 'sp4_v_b_6')
// (15, 3, 'sp4_v_t_36')
// (15, 4, 'sp4_h_l_36')
// (15, 4, 'sp4_h_r_1')
// (15, 4, 'sp4_h_r_15')
// (15, 4, 'sp4_v_b_36')
// (15, 5, 'sp4_v_b_25')
// (15, 6, 'sp4_v_b_12')
// (15, 7, 'sp4_v_b_1')
// (15, 12, 'sp4_h_r_21')
// (16, 3, 'sp4_h_r_12')
// (16, 3, 'sp4_h_r_44')
// (16, 4, 'sp4_h_r_12')
// (16, 4, 'sp4_h_r_26')
// (16, 4, 'sp4_r_v_b_38')
// (16, 5, 'sp4_r_v_b_27')
// (16, 6, 'sp4_r_v_b_14')
// (16, 7, 'sp4_r_v_b_3')
// (16, 12, 'sp4_h_r_32')
// (17, 1, 'sp4_r_v_b_44')
// (17, 2, 'neigh_op_tnr_2')
// (17, 2, 'sp4_r_v_b_33')
// (17, 3, 'neigh_op_rgt_2')
// (17, 3, 'sp4_h_l_44')
// (17, 3, 'sp4_h_r_25')
// (17, 3, 'sp4_h_r_9')
// (17, 3, 'sp4_r_v_b_20')
// (17, 3, 'sp4_v_t_38')
// (17, 4, 'neigh_op_bnr_2')
// (17, 4, 'sp4_h_r_25')
// (17, 4, 'sp4_h_r_39')
// (17, 4, 'sp4_r_v_b_9')
// (17, 4, 'sp4_v_b_38')
// (17, 5, 'sp4_r_v_b_37')
// (17, 5, 'sp4_v_b_27')
// (17, 6, 'sp4_r_v_b_24')
// (17, 6, 'sp4_v_b_14')
// (17, 7, 'local_g1_3')
// (17, 7, 'lutff_0/in_2')
// (17, 7, 'sp4_r_v_b_13')
// (17, 7, 'sp4_v_b_3')
// (17, 8, 'sp4_r_v_b_0')
// (17, 9, 'sp4_r_v_b_38')
// (17, 10, 'sp4_r_v_b_27')
// (17, 11, 'sp4_r_v_b_14')
// (17, 12, 'sp4_h_r_45')
// (17, 12, 'sp4_r_v_b_3')
// (18, 0, 'span4_vert_44')
// (18, 1, 'sp4_r_v_b_45')
// (18, 1, 'sp4_v_b_44')
// (18, 2, 'neigh_op_top_2')
// (18, 2, 'sp4_r_v_b_32')
// (18, 2, 'sp4_v_b_33')
// (18, 3, 'local_g3_2')
// (18, 3, 'lutff_2/in_3')
// (18, 3, 'lutff_2/out')
// (18, 3, 'sp4_h_r_20')
// (18, 3, 'sp4_h_r_36')
// (18, 3, 'sp4_r_v_b_21')
// (18, 3, 'sp4_v_b_20')
// (18, 4, 'neigh_op_bot_2')
// (18, 4, 'sp4_h_l_39')
// (18, 4, 'sp4_h_r_36')
// (18, 4, 'sp4_r_v_b_8')
// (18, 4, 'sp4_v_b_9')
// (18, 4, 'sp4_v_t_37')
// (18, 5, 'sp4_v_b_37')
// (18, 6, 'sp4_v_b_24')
// (18, 7, 'sp4_v_b_13')
// (18, 8, 'sp4_v_b_0')
// (18, 8, 'sp4_v_t_38')
// (18, 9, 'sp4_v_b_38')
// (18, 10, 'sp4_v_b_27')
// (18, 11, 'sp4_v_b_14')
// (18, 12, 'sp4_h_l_45')
// (18, 12, 'sp4_v_b_3')
// (19, 0, 'span4_vert_45')
// (19, 1, 'sp4_v_b_45')
// (19, 2, 'neigh_op_tnl_2')
// (19, 2, 'sp4_v_b_32')
// (19, 3, 'neigh_op_lft_2')
// (19, 3, 'sp4_h_l_36')
// (19, 3, 'sp4_h_r_33')
// (19, 3, 'sp4_v_b_21')
// (19, 4, 'neigh_op_bnl_2')
// (19, 4, 'sp4_h_l_36')
// (19, 4, 'sp4_v_b_8')
// (20, 3, 'sp4_h_r_44')
// (21, 3, 'sp4_h_l_44')

wire n853;
// (6, 6, 'neigh_op_tnr_0')
// (6, 7, 'neigh_op_rgt_0')
// (6, 8, 'neigh_op_bnr_0')
// (7, 6, 'neigh_op_top_0')
// (7, 7, 'local_g0_0')
// (7, 7, 'lutff_0/out')
// (7, 7, 'lutff_6/in_2')
// (7, 8, 'neigh_op_bot_0')
// (8, 6, 'neigh_op_tnl_0')
// (8, 7, 'neigh_op_lft_0')
// (8, 8, 'neigh_op_bnl_0')

wire n854;
// (6, 6, 'neigh_op_tnr_1')
// (6, 7, 'neigh_op_rgt_1')
// (6, 8, 'neigh_op_bnr_1')
// (7, 6, 'neigh_op_top_1')
// (7, 6, 'sp4_r_v_b_46')
// (7, 7, 'lutff_1/out')
// (7, 7, 'sp4_r_v_b_35')
// (7, 8, 'neigh_op_bot_1')
// (7, 8, 'sp4_r_v_b_22')
// (7, 9, 'local_g2_3')
// (7, 9, 'lutff_7/in_2')
// (7, 9, 'sp4_r_v_b_11')
// (8, 5, 'sp4_v_t_46')
// (8, 6, 'neigh_op_tnl_1')
// (8, 6, 'sp4_v_b_46')
// (8, 7, 'local_g0_1')
// (8, 7, 'lutff_6/in_1')
// (8, 7, 'neigh_op_lft_1')
// (8, 7, 'sp4_v_b_35')
// (8, 8, 'neigh_op_bnl_1')
// (8, 8, 'sp4_v_b_22')
// (8, 9, 'sp4_v_b_11')

wire n855;
// (6, 6, 'neigh_op_tnr_2')
// (6, 7, 'neigh_op_rgt_2')
// (6, 8, 'neigh_op_bnr_2')
// (7, 6, 'neigh_op_top_2')
// (7, 7, 'lutff_2/out')
// (7, 8, 'neigh_op_bot_2')
// (8, 6, 'neigh_op_tnl_2')
// (8, 7, 'local_g1_2')
// (8, 7, 'lutff_3/in_2')
// (8, 7, 'neigh_op_lft_2')
// (8, 8, 'neigh_op_bnl_2')

reg n856 = 0;
// (6, 6, 'neigh_op_tnr_3')
// (6, 7, 'neigh_op_rgt_3')
// (6, 8, 'neigh_op_bnr_3')
// (7, 6, 'neigh_op_top_3')
// (7, 7, 'local_g0_3')
// (7, 7, 'lutff_3/out')
// (7, 7, 'lutff_5/in_0')
// (7, 8, 'neigh_op_bot_3')
// (8, 6, 'neigh_op_tnl_3')
// (8, 7, 'neigh_op_lft_3')
// (8, 8, 'neigh_op_bnl_3')

wire n857;
// (6, 6, 'neigh_op_tnr_4')
// (6, 7, 'neigh_op_rgt_4')
// (6, 8, 'neigh_op_bnr_4')
// (7, 6, 'neigh_op_top_4')
// (7, 7, 'local_g2_4')
// (7, 7, 'lutff_4/out')
// (7, 7, 'lutff_6/in_0')
// (7, 8, 'neigh_op_bot_4')
// (8, 6, 'neigh_op_tnl_4')
// (8, 7, 'neigh_op_lft_4')
// (8, 8, 'neigh_op_bnl_4')

wire n858;
// (6, 6, 'neigh_op_tnr_5')
// (6, 7, 'neigh_op_rgt_5')
// (6, 8, 'neigh_op_bnr_5')
// (7, 6, 'neigh_op_top_5')
// (7, 7, 'lutff_5/out')
// (7, 7, 'sp4_h_r_10')
// (7, 8, 'neigh_op_bot_5')
// (8, 6, 'neigh_op_tnl_5')
// (8, 7, 'neigh_op_lft_5')
// (8, 7, 'sp4_h_r_23')
// (8, 8, 'neigh_op_bnl_5')
// (9, 7, 'sp4_h_r_34')
// (10, 7, 'local_g2_7')
// (10, 7, 'lutff_3/in_2')
// (10, 7, 'sp4_h_r_47')
// (11, 7, 'sp4_h_l_47')

wire n859;
// (6, 6, 'neigh_op_tnr_6')
// (6, 7, 'neigh_op_rgt_6')
// (6, 8, 'neigh_op_bnr_6')
// (7, 6, 'neigh_op_top_6')
// (7, 7, 'local_g3_6')
// (7, 7, 'lutff_1/in_2')
// (7, 7, 'lutff_6/out')
// (7, 8, 'neigh_op_bot_6')
// (8, 6, 'neigh_op_tnl_6')
// (8, 7, 'neigh_op_lft_6')
// (8, 8, 'neigh_op_bnl_6')

wire n860;
// (6, 6, 'neigh_op_tnr_7')
// (6, 7, 'neigh_op_rgt_7')
// (6, 8, 'neigh_op_bnr_7')
// (7, 6, 'neigh_op_top_7')
// (7, 7, 'lutff_7/out')
// (7, 8, 'neigh_op_bot_7')
// (8, 6, 'neigh_op_tnl_7')
// (8, 7, 'local_g0_7')
// (8, 7, 'lutff_4/in_1')
// (8, 7, 'neigh_op_lft_7')
// (8, 8, 'neigh_op_bnl_7')

wire n861;
// (6, 6, 'sp4_h_r_1')
// (7, 3, 'sp4_r_v_b_44')
// (7, 4, 'local_g2_1')
// (7, 4, 'lutff_0/in_1')
// (7, 4, 'sp4_r_v_b_33')
// (7, 5, 'sp4_r_v_b_20')
// (7, 6, 'local_g1_4')
// (7, 6, 'lutff_0/in_3')
// (7, 6, 'lutff_5/in_2')
// (7, 6, 'sp4_h_r_12')
// (7, 6, 'sp4_r_v_b_9')
// (8, 2, 'sp4_v_t_44')
// (8, 3, 'sp4_r_v_b_41')
// (8, 3, 'sp4_v_b_44')
// (8, 4, 'local_g1_4')
// (8, 4, 'lutff_3/in_0')
// (8, 4, 'sp4_r_v_b_28')
// (8, 4, 'sp4_v_b_33')
// (8, 5, 'neigh_op_tnr_2')
// (8, 5, 'sp4_r_v_b_17')
// (8, 5, 'sp4_v_b_20')
// (8, 6, 'local_g3_2')
// (8, 6, 'lutff_3/in_0')
// (8, 6, 'lutff_4/in_3')
// (8, 6, 'neigh_op_rgt_2')
// (8, 6, 'sp4_h_r_25')
// (8, 6, 'sp4_h_r_9')
// (8, 6, 'sp4_r_v_b_4')
// (8, 6, 'sp4_v_b_9')
// (8, 7, 'neigh_op_bnr_2')
// (9, 2, 'sp4_v_t_41')
// (9, 3, 'sp4_v_b_41')
// (9, 4, 'sp4_v_b_28')
// (9, 5, 'neigh_op_top_2')
// (9, 5, 'sp4_v_b_17')
// (9, 6, 'lutff_2/out')
// (9, 6, 'sp4_h_r_20')
// (9, 6, 'sp4_h_r_36')
// (9, 6, 'sp4_v_b_4')
// (9, 7, 'neigh_op_bot_2')
// (10, 5, 'local_g2_2')
// (10, 5, 'lutff_1/in_1')
// (10, 5, 'neigh_op_tnl_2')
// (10, 6, 'neigh_op_lft_2')
// (10, 6, 'sp4_h_l_36')
// (10, 6, 'sp4_h_r_33')
// (10, 7, 'neigh_op_bnl_2')
// (11, 6, 'sp4_h_r_44')
// (12, 6, 'sp4_h_l_44')

wire n862;
// (6, 6, 'sp4_r_v_b_41')
// (6, 7, 'sp4_r_v_b_28')
// (6, 8, 'neigh_op_tnr_2')
// (6, 8, 'sp4_r_v_b_17')
// (6, 9, 'neigh_op_rgt_2')
// (6, 9, 'sp4_r_v_b_4')
// (6, 10, 'neigh_op_bnr_2')
// (7, 5, 'sp4_v_t_41')
// (7, 6, 'sp4_r_v_b_40')
// (7, 6, 'sp4_v_b_41')
// (7, 7, 'local_g3_4')
// (7, 7, 'lutff_4/in_1')
// (7, 7, 'sp4_r_v_b_29')
// (7, 7, 'sp4_v_b_28')
// (7, 8, 'neigh_op_top_2')
// (7, 8, 'sp4_r_v_b_16')
// (7, 8, 'sp4_v_b_17')
// (7, 9, 'lutff_2/out')
// (7, 9, 'sp4_r_v_b_5')
// (7, 9, 'sp4_v_b_4')
// (7, 10, 'neigh_op_bot_2')
// (8, 5, 'sp4_v_t_40')
// (8, 6, 'sp4_v_b_40')
// (8, 7, 'local_g3_5')
// (8, 7, 'lutff_2/in_2')
// (8, 7, 'sp4_v_b_29')
// (8, 8, 'neigh_op_tnl_2')
// (8, 8, 'sp4_v_b_16')
// (8, 9, 'neigh_op_lft_2')
// (8, 9, 'sp4_v_b_5')
// (8, 10, 'neigh_op_bnl_2')

wire n863;
// (6, 6, 'sp4_r_v_b_43')
// (6, 7, 'sp4_r_v_b_30')
// (6, 8, 'neigh_op_tnr_3')
// (6, 8, 'sp4_r_v_b_19')
// (6, 9, 'neigh_op_rgt_3')
// (6, 9, 'sp4_r_v_b_6')
// (6, 10, 'neigh_op_bnr_3')
// (7, 5, 'sp4_v_t_43')
// (7, 6, 'sp4_r_v_b_42')
// (7, 6, 'sp4_v_b_43')
// (7, 7, 'local_g2_6')
// (7, 7, 'lutff_1/in_3')
// (7, 7, 'sp4_r_v_b_31')
// (7, 7, 'sp4_v_b_30')
// (7, 8, 'neigh_op_top_3')
// (7, 8, 'sp4_r_v_b_18')
// (7, 8, 'sp4_v_b_19')
// (7, 9, 'lutff_3/out')
// (7, 9, 'sp4_r_v_b_7')
// (7, 9, 'sp4_v_b_6')
// (7, 10, 'neigh_op_bot_3')
// (8, 5, 'sp4_v_t_42')
// (8, 6, 'sp4_v_b_42')
// (8, 7, 'local_g3_7')
// (8, 7, 'lutff_3/in_1')
// (8, 7, 'sp4_v_b_31')
// (8, 8, 'neigh_op_tnl_3')
// (8, 8, 'sp4_v_b_18')
// (8, 9, 'neigh_op_lft_3')
// (8, 9, 'sp4_v_b_7')
// (8, 10, 'neigh_op_bnl_3')

wire n864;
// (6, 6, 'sp4_r_v_b_45')
// (6, 7, 'sp4_r_v_b_32')
// (6, 8, 'neigh_op_tnr_4')
// (6, 8, 'sp4_r_v_b_21')
// (6, 9, 'neigh_op_rgt_4')
// (6, 9, 'sp4_r_v_b_8')
// (6, 10, 'neigh_op_bnr_4')
// (7, 5, 'sp4_v_t_45')
// (7, 6, 'sp4_v_b_45')
// (7, 7, 'local_g2_0')
// (7, 7, 'lutff_0/in_2')
// (7, 7, 'sp4_v_b_32')
// (7, 8, 'neigh_op_top_4')
// (7, 8, 'sp4_r_v_b_36')
// (7, 8, 'sp4_v_b_21')
// (7, 9, 'lutff_4/out')
// (7, 9, 'sp4_r_v_b_25')
// (7, 9, 'sp4_v_b_8')
// (7, 10, 'neigh_op_bot_4')
// (7, 10, 'sp4_r_v_b_12')
// (7, 11, 'sp4_r_v_b_1')
// (8, 7, 'local_g0_6')
// (8, 7, 'lutff_4/in_2')
// (8, 7, 'sp4_h_r_6')
// (8, 7, 'sp4_v_t_36')
// (8, 8, 'neigh_op_tnl_4')
// (8, 8, 'sp4_v_b_36')
// (8, 9, 'neigh_op_lft_4')
// (8, 9, 'sp4_v_b_25')
// (8, 10, 'neigh_op_bnl_4')
// (8, 10, 'sp4_v_b_12')
// (8, 11, 'sp4_v_b_1')
// (9, 7, 'sp4_h_r_19')
// (10, 7, 'sp4_h_r_30')
// (11, 7, 'sp4_h_r_43')
// (12, 7, 'sp4_h_l_43')

reg n865 = 0;
// (6, 7, 'neigh_op_tnr_1')
// (6, 8, 'neigh_op_rgt_1')
// (6, 9, 'neigh_op_bnr_1')
// (7, 7, 'local_g1_1')
// (7, 7, 'lutff_4/in_0')
// (7, 7, 'neigh_op_top_1')
// (7, 8, 'local_g3_1')
// (7, 8, 'lutff_1/in_1')
// (7, 8, 'lutff_1/out')
// (7, 9, 'neigh_op_bot_1')
// (8, 7, 'local_g2_1')
// (8, 7, 'lutff_7/in_2')
// (8, 7, 'neigh_op_tnl_1')
// (8, 8, 'neigh_op_lft_1')
// (8, 9, 'neigh_op_bnl_1')

reg n866 = 0;
// (6, 7, 'neigh_op_tnr_2')
// (6, 8, 'neigh_op_rgt_2')
// (6, 9, 'neigh_op_bnr_2')
// (7, 7, 'neigh_op_top_2')
// (7, 8, 'local_g1_2')
// (7, 8, 'lutff_2/in_1')
// (7, 8, 'lutff_2/out')
// (7, 9, 'neigh_op_bot_2')
// (8, 7, 'neigh_op_tnl_2')
// (8, 8, 'local_g1_2')
// (8, 8, 'lutff_6/in_3')
// (8, 8, 'lutff_7/in_2')
// (8, 8, 'neigh_op_lft_2')
// (8, 9, 'neigh_op_bnl_2')

reg n867 = 0;
// (6, 7, 'neigh_op_tnr_3')
// (6, 8, 'neigh_op_rgt_3')
// (6, 9, 'neigh_op_bnr_3')
// (7, 7, 'local_g1_3')
// (7, 7, 'lutff_4/in_2')
// (7, 7, 'neigh_op_top_3')
// (7, 8, 'local_g3_3')
// (7, 8, 'lutff_3/in_1')
// (7, 8, 'lutff_3/out')
// (7, 9, 'neigh_op_bot_3')
// (8, 7, 'neigh_op_tnl_3')
// (8, 8, 'local_g1_3')
// (8, 8, 'lutff_0/in_0')
// (8, 8, 'neigh_op_lft_3')
// (8, 9, 'neigh_op_bnl_3')

reg n868 = 0;
// (6, 7, 'neigh_op_tnr_4')
// (6, 8, 'neigh_op_rgt_4')
// (6, 9, 'neigh_op_bnr_4')
// (7, 7, 'local_g0_4')
// (7, 7, 'lutff_1/in_1')
// (7, 7, 'lutff_2/in_2')
// (7, 7, 'neigh_op_top_4')
// (7, 8, 'local_g3_4')
// (7, 8, 'lutff_4/in_1')
// (7, 8, 'lutff_4/out')
// (7, 9, 'neigh_op_bot_4')
// (8, 7, 'neigh_op_tnl_4')
// (8, 8, 'neigh_op_lft_4')
// (8, 9, 'neigh_op_bnl_4')

reg n869 = 0;
// (6, 7, 'neigh_op_tnr_5')
// (6, 8, 'neigh_op_rgt_5')
// (6, 9, 'neigh_op_bnr_5')
// (7, 7, 'local_g0_5')
// (7, 7, 'lutff_0/in_3')
// (7, 7, 'lutff_7/in_2')
// (7, 7, 'neigh_op_top_5')
// (7, 8, 'local_g2_5')
// (7, 8, 'lutff_5/in_2')
// (7, 8, 'lutff_5/out')
// (7, 9, 'neigh_op_bot_5')
// (8, 7, 'neigh_op_tnl_5')
// (8, 8, 'neigh_op_lft_5')
// (8, 9, 'neigh_op_bnl_5')

reg n870 = 0;
// (6, 7, 'neigh_op_tnr_6')
// (6, 8, 'neigh_op_rgt_6')
// (6, 9, 'neigh_op_bnr_6')
// (7, 7, 'neigh_op_top_6')
// (7, 8, 'local_g2_6')
// (7, 8, 'lutff_6/in_0')
// (7, 8, 'lutff_6/out')
// (7, 9, 'neigh_op_bot_6')
// (8, 7, 'neigh_op_tnl_6')
// (8, 8, 'local_g0_6')
// (8, 8, 'local_g1_6')
// (8, 8, 'lutff_3/in_1')
// (8, 8, 'lutff_7/in_0')
// (8, 8, 'neigh_op_lft_6')
// (8, 9, 'neigh_op_bnl_6')

reg n871 = 0;
// (6, 7, 'neigh_op_tnr_7')
// (6, 8, 'neigh_op_rgt_7')
// (6, 9, 'neigh_op_bnr_7')
// (7, 7, 'local_g0_7')
// (7, 7, 'lutff_6/in_1')
// (7, 7, 'neigh_op_top_7')
// (7, 8, 'local_g1_7')
// (7, 8, 'local_g2_7')
// (7, 8, 'lutff_0/in_1')
// (7, 8, 'lutff_1/in_3')
// (7, 8, 'lutff_7/in_0')
// (7, 8, 'lutff_7/out')
// (7, 9, 'neigh_op_bot_7')
// (8, 7, 'neigh_op_tnl_7')
// (8, 8, 'neigh_op_lft_7')
// (8, 9, 'neigh_op_bnl_7')

reg n872 = 0;
// (6, 7, 'sp4_r_v_b_39')
// (6, 8, 'sp4_r_v_b_26')
// (6, 9, 'neigh_op_tnr_1')
// (6, 9, 'sp4_r_v_b_15')
// (6, 10, 'neigh_op_rgt_1')
// (6, 10, 'sp4_r_v_b_2')
// (6, 11, 'neigh_op_bnr_1')
// (7, 6, 'sp4_v_t_39')
// (7, 7, 'local_g3_7')
// (7, 7, 'lutff_5/in_1')
// (7, 7, 'sp4_v_b_39')
// (7, 8, 'sp4_v_b_26')
// (7, 9, 'neigh_op_top_1')
// (7, 9, 'sp4_v_b_15')
// (7, 10, 'lutff_1/out')
// (7, 10, 'sp4_v_b_2')
// (7, 11, 'neigh_op_bot_1')
// (8, 9, 'neigh_op_tnl_1')
// (8, 10, 'neigh_op_lft_1')
// (8, 11, 'neigh_op_bnl_1')

wire n873;
// (6, 8, 'neigh_op_tnr_1')
// (6, 9, 'neigh_op_rgt_1')
// (6, 10, 'neigh_op_bnr_1')
// (7, 6, 'sp4_r_v_b_38')
// (7, 7, 'sp4_r_v_b_27')
// (7, 8, 'neigh_op_top_1')
// (7, 8, 'sp4_r_v_b_14')
// (7, 9, 'lutff_1/out')
// (7, 9, 'sp4_r_v_b_3')
// (7, 10, 'neigh_op_bot_1')
// (8, 5, 'sp4_v_t_38')
// (8, 6, 'sp4_v_b_38')
// (8, 7, 'local_g3_3')
// (8, 7, 'lutff_1/in_1')
// (8, 7, 'sp4_v_b_27')
// (8, 8, 'local_g3_1')
// (8, 8, 'lutff_7/in_1')
// (8, 8, 'neigh_op_tnl_1')
// (8, 8, 'sp4_v_b_14')
// (8, 9, 'neigh_op_lft_1')
// (8, 9, 'sp4_v_b_3')
// (8, 10, 'neigh_op_bnl_1')

wire n874;
// (6, 8, 'neigh_op_tnr_5')
// (6, 9, 'neigh_op_rgt_5')
// (6, 10, 'neigh_op_bnr_5')
// (7, 8, 'neigh_op_top_5')
// (7, 9, 'lutff_5/out')
// (7, 10, 'neigh_op_bot_5')
// (8, 8, 'neigh_op_tnl_5')
// (8, 9, 'local_g0_5')
// (8, 9, 'lutff_5/in_0')
// (8, 9, 'neigh_op_lft_5')
// (8, 10, 'neigh_op_bnl_5')

wire n875;
// (6, 8, 'neigh_op_tnr_6')
// (6, 9, 'neigh_op_rgt_6')
// (6, 10, 'neigh_op_bnr_6')
// (7, 8, 'neigh_op_top_6')
// (7, 9, 'local_g2_6')
// (7, 9, 'local_g3_6')
// (7, 9, 'lutff_0/in_1')
// (7, 9, 'lutff_1/in_3')
// (7, 9, 'lutff_6/out')
// (7, 10, 'neigh_op_bot_6')
// (8, 8, 'neigh_op_tnl_6')
// (8, 9, 'neigh_op_lft_6')
// (8, 10, 'neigh_op_bnl_6')

reg n876 = 0;
// (6, 8, 'sp4_h_r_10')
// (7, 7, 'neigh_op_tnr_1')
// (7, 8, 'neigh_op_rgt_1')
// (7, 8, 'sp4_h_r_23')
// (7, 9, 'neigh_op_bnr_1')
// (8, 7, 'neigh_op_top_1')
// (8, 8, 'lutff_1/out')
// (8, 8, 'sp4_h_r_34')
// (8, 9, 'local_g0_1')
// (8, 9, 'lutff_3/in_2')
// (8, 9, 'neigh_op_bot_1')
// (9, 5, 'sp4_r_v_b_47')
// (9, 6, 'sp4_r_v_b_34')
// (9, 7, 'neigh_op_tnl_1')
// (9, 7, 'sp4_r_v_b_23')
// (9, 8, 'neigh_op_lft_1')
// (9, 8, 'sp4_h_r_47')
// (9, 8, 'sp4_r_v_b_10')
// (9, 9, 'local_g3_1')
// (9, 9, 'lutff_1/in_1')
// (9, 9, 'neigh_op_bnl_1')
// (10, 4, 'sp4_v_t_47')
// (10, 5, 'sp4_v_b_47')
// (10, 6, 'sp4_v_b_34')
// (10, 7, 'local_g0_7')
// (10, 7, 'lutff_0/in_3')
// (10, 7, 'sp4_v_b_23')
// (10, 8, 'sp4_h_l_47')
// (10, 8, 'sp4_v_b_10')

wire n877;
// (6, 8, 'sp4_h_r_11')
// (7, 8, 'sp4_h_r_22')
// (8, 6, 'neigh_op_tnr_1')
// (8, 6, 'sp4_r_v_b_47')
// (8, 7, 'neigh_op_rgt_1')
// (8, 7, 'sp4_h_r_7')
// (8, 7, 'sp4_r_v_b_34')
// (8, 8, 'local_g3_3')
// (8, 8, 'lutff_global/cen')
// (8, 8, 'neigh_op_bnr_1')
// (8, 8, 'sp4_h_r_35')
// (8, 8, 'sp4_r_v_b_23')
// (8, 9, 'local_g2_2')
// (8, 9, 'lutff_global/cen')
// (8, 9, 'sp4_r_v_b_10')
// (9, 5, 'sp4_r_v_b_43')
// (9, 5, 'sp4_v_t_47')
// (9, 6, 'neigh_op_top_1')
// (9, 6, 'sp4_r_v_b_30')
// (9, 6, 'sp4_v_b_47')
// (9, 7, 'local_g0_2')
// (9, 7, 'lutff_1/out')
// (9, 7, 'lutff_global/cen')
// (9, 7, 'sp4_h_r_18')
// (9, 7, 'sp4_r_v_b_19')
// (9, 7, 'sp4_v_b_34')
// (9, 8, 'neigh_op_bot_1')
// (9, 8, 'sp4_h_r_46')
// (9, 8, 'sp4_r_v_b_6')
// (9, 8, 'sp4_v_b_23')
// (9, 9, 'sp4_v_b_10')
// (10, 4, 'sp4_v_t_43')
// (10, 5, 'sp4_v_b_43')
// (10, 6, 'neigh_op_tnl_1')
// (10, 6, 'sp4_v_b_30')
// (10, 7, 'neigh_op_lft_1')
// (10, 7, 'sp4_h_r_31')
// (10, 7, 'sp4_v_b_19')
// (10, 8, 'neigh_op_bnl_1')
// (10, 8, 'sp4_h_l_46')
// (10, 8, 'sp4_v_b_6')
// (11, 7, 'sp4_h_r_42')
// (12, 7, 'sp4_h_l_42')

reg n878 = 0;
// (6, 8, 'sp4_h_r_2')
// (7, 7, 'neigh_op_tnr_5')
// (7, 8, 'neigh_op_rgt_5')
// (7, 8, 'sp4_h_r_15')
// (7, 9, 'neigh_op_bnr_5')
// (8, 7, 'neigh_op_top_5')
// (8, 8, 'lutff_5/out')
// (8, 8, 'sp4_h_r_26')
// (8, 9, 'local_g1_5')
// (8, 9, 'lutff_2/in_2')
// (8, 9, 'neigh_op_bot_5')
// (9, 7, 'neigh_op_tnl_5')
// (9, 8, 'local_g3_7')
// (9, 8, 'lutff_3/in_3')
// (9, 8, 'neigh_op_lft_5')
// (9, 8, 'sp4_h_r_39')
// (9, 9, 'local_g2_5')
// (9, 9, 'lutff_6/in_1')
// (9, 9, 'neigh_op_bnl_5')
// (10, 8, 'sp4_h_l_39')

reg n879 = 0;
// (6, 9, 'neigh_op_tnr_3')
// (6, 10, 'neigh_op_rgt_3')
// (6, 11, 'neigh_op_bnr_3')
// (7, 9, 'neigh_op_top_3')
// (7, 10, 'lutff_3/out')
// (7, 11, 'neigh_op_bot_3')
// (8, 9, 'neigh_op_tnl_3')
// (8, 10, 'local_g1_3')
// (8, 10, 'lutff_6/in_2')
// (8, 10, 'neigh_op_lft_3')
// (8, 11, 'neigh_op_bnl_3')

reg n880 = 0;
// (6, 9, 'sp4_h_r_6')
// (7, 8, 'neigh_op_tnr_7')
// (7, 9, 'neigh_op_rgt_7')
// (7, 9, 'sp4_h_r_19')
// (7, 9, 'sp4_h_r_3')
// (7, 10, 'neigh_op_bnr_7')
// (8, 8, 'neigh_op_top_7')
// (8, 9, 'local_g3_7')
// (8, 9, 'lutff_1/in_1')
// (8, 9, 'lutff_7/out')
// (8, 9, 'sp4_h_r_14')
// (8, 9, 'sp4_h_r_30')
// (8, 10, 'neigh_op_bot_7')
// (9, 8, 'neigh_op_tnl_7')
// (9, 9, 'neigh_op_lft_7')
// (9, 9, 'sp4_h_r_27')
// (9, 9, 'sp4_h_r_43')
// (9, 10, 'neigh_op_bnl_7')
// (9, 10, 'sp4_r_v_b_43')
// (9, 11, 'sp4_r_v_b_30')
// (9, 12, 'sp4_r_v_b_19')
// (9, 13, 'sp4_r_v_b_6')
// (10, 9, 'local_g2_6')
// (10, 9, 'lutff_4/in_0')
// (10, 9, 'sp4_h_l_43')
// (10, 9, 'sp4_h_r_38')
// (10, 9, 'sp4_v_t_43')
// (10, 10, 'local_g3_3')
// (10, 10, 'lutff_2/in_0')
// (10, 10, 'sp4_v_b_43')
// (10, 11, 'sp4_v_b_30')
// (10, 12, 'sp4_v_b_19')
// (10, 13, 'sp4_v_b_6')
// (11, 9, 'sp4_h_l_38')

reg n881 = 0;
// (6, 10, 'neigh_op_tnr_0')
// (6, 11, 'neigh_op_rgt_0')
// (6, 12, 'neigh_op_bnr_0')
// (7, 10, 'neigh_op_top_0')
// (7, 11, 'lutff_0/out')
// (7, 12, 'local_g1_0')
// (7, 12, 'lutff_7/in_2')
// (7, 12, 'neigh_op_bot_0')
// (8, 10, 'neigh_op_tnl_0')
// (8, 11, 'neigh_op_lft_0')
// (8, 12, 'neigh_op_bnl_0')

reg n882 = 0;
// (6, 10, 'neigh_op_tnr_1')
// (6, 11, 'neigh_op_rgt_1')
// (6, 12, 'neigh_op_bnr_1')
// (7, 10, 'neigh_op_top_1')
// (7, 11, 'lutff_1/out')
// (7, 12, 'neigh_op_bot_1')
// (8, 10, 'neigh_op_tnl_1')
// (8, 11, 'local_g0_1')
// (8, 11, 'lutff_5/in_2')
// (8, 11, 'neigh_op_lft_1')
// (8, 12, 'neigh_op_bnl_1')

reg n883 = 0;
// (6, 10, 'neigh_op_tnr_2')
// (6, 11, 'neigh_op_rgt_2')
// (6, 12, 'neigh_op_bnr_2')
// (7, 10, 'neigh_op_top_2')
// (7, 11, 'lutff_2/out')
// (7, 12, 'local_g1_2')
// (7, 12, 'lutff_2/in_3')
// (7, 12, 'neigh_op_bot_2')
// (8, 10, 'neigh_op_tnl_2')
// (8, 11, 'neigh_op_lft_2')
// (8, 12, 'neigh_op_bnl_2')

reg n884 = 0;
// (6, 10, 'neigh_op_tnr_5')
// (6, 11, 'neigh_op_rgt_5')
// (6, 12, 'neigh_op_bnr_5')
// (7, 10, 'neigh_op_top_5')
// (7, 11, 'lutff_5/out')
// (7, 12, 'local_g1_5')
// (7, 12, 'lutff_2/in_2')
// (7, 12, 'neigh_op_bot_5')
// (8, 10, 'neigh_op_tnl_5')
// (8, 11, 'neigh_op_lft_5')
// (8, 12, 'neigh_op_bnl_5')

reg n885 = 0;
// (6, 11, 'neigh_op_tnr_1')
// (6, 12, 'neigh_op_rgt_1')
// (6, 13, 'neigh_op_bnr_1')
// (7, 11, 'local_g0_1')
// (7, 11, 'lutff_1/in_0')
// (7, 11, 'neigh_op_top_1')
// (7, 12, 'lutff_1/out')
// (7, 13, 'neigh_op_bot_1')
// (8, 11, 'neigh_op_tnl_1')
// (8, 12, 'neigh_op_lft_1')
// (8, 13, 'neigh_op_bnl_1')

wire n886;
// (6, 11, 'neigh_op_tnr_2')
// (6, 12, 'neigh_op_rgt_2')
// (6, 13, 'neigh_op_bnr_2')
// (7, 11, 'neigh_op_top_2')
// (7, 12, 'lutff_2/out')
// (7, 12, 'sp4_r_v_b_37')
// (7, 13, 'neigh_op_bot_2')
// (7, 13, 'sp4_r_v_b_24')
// (7, 14, 'sp4_r_v_b_13')
// (7, 15, 'sp4_r_v_b_0')
// (8, 11, 'neigh_op_tnl_2')
// (8, 11, 'sp4_v_t_37')
// (8, 12, 'neigh_op_lft_2')
// (8, 12, 'sp4_v_b_37')
// (8, 13, 'neigh_op_bnl_2')
// (8, 13, 'sp4_v_b_24')
// (8, 14, 'sp4_v_b_13')
// (8, 15, 'sp4_h_r_0')
// (8, 15, 'sp4_v_b_0')
// (9, 15, 'local_g0_5')
// (9, 15, 'lutff_2/in_3')
// (9, 15, 'sp4_h_r_13')
// (10, 15, 'sp4_h_r_24')
// (11, 15, 'sp4_h_r_37')
// (12, 15, 'sp4_h_l_37')

reg n887 = 0;
// (6, 11, 'neigh_op_tnr_3')
// (6, 12, 'neigh_op_rgt_3')
// (6, 13, 'neigh_op_bnr_3')
// (7, 11, 'neigh_op_top_3')
// (7, 12, 'lutff_3/out')
// (7, 13, 'local_g0_3')
// (7, 13, 'lutff_2/in_3')
// (7, 13, 'neigh_op_bot_3')
// (8, 11, 'neigh_op_tnl_3')
// (8, 12, 'neigh_op_lft_3')
// (8, 13, 'neigh_op_bnl_3')

reg n888 = 0;
// (6, 11, 'neigh_op_tnr_4')
// (6, 12, 'neigh_op_rgt_4')
// (6, 13, 'neigh_op_bnr_4')
// (7, 11, 'neigh_op_top_4')
// (7, 12, 'lutff_4/out')
// (7, 13, 'local_g1_4')
// (7, 13, 'lutff_5/in_2')
// (7, 13, 'neigh_op_bot_4')
// (8, 11, 'neigh_op_tnl_4')
// (8, 12, 'neigh_op_lft_4')
// (8, 13, 'neigh_op_bnl_4')

reg n889 = 0;
// (6, 11, 'neigh_op_tnr_5')
// (6, 12, 'neigh_op_rgt_5')
// (6, 13, 'neigh_op_bnr_5')
// (7, 11, 'local_g0_5')
// (7, 11, 'lutff_5/in_0')
// (7, 11, 'neigh_op_top_5')
// (7, 12, 'lutff_5/out')
// (7, 13, 'neigh_op_bot_5')
// (8, 11, 'neigh_op_tnl_5')
// (8, 12, 'neigh_op_lft_5')
// (8, 13, 'neigh_op_bnl_5')

wire n890;
// (6, 11, 'neigh_op_tnr_7')
// (6, 12, 'neigh_op_rgt_7')
// (6, 13, 'neigh_op_bnr_7')
// (7, 11, 'neigh_op_top_7')
// (7, 12, 'local_g3_7')
// (7, 12, 'lutff_2/in_0')
// (7, 12, 'lutff_7/out')
// (7, 13, 'neigh_op_bot_7')
// (8, 11, 'neigh_op_tnl_7')
// (8, 12, 'neigh_op_lft_7')
// (8, 13, 'neigh_op_bnl_7')

wire n891;
// (6, 11, 'sp4_h_r_5')
// (7, 11, 'local_g0_0')
// (7, 11, 'lutff_6/in_2')
// (7, 11, 'sp4_h_r_16')
// (8, 5, 'neigh_op_tnr_7')
// (8, 6, 'local_g2_7')
// (8, 6, 'local_g3_7')
// (8, 6, 'lutff_5/in_3')
// (8, 6, 'lutff_6/in_3')
// (8, 6, 'neigh_op_rgt_7')
// (8, 7, 'neigh_op_bnr_7')
// (8, 11, 'sp4_h_r_29')
// (9, 4, 'sp4_r_v_b_39')
// (9, 5, 'neigh_op_top_7')
// (9, 5, 'sp4_r_v_b_26')
// (9, 6, 'lutff_7/out')
// (9, 6, 'sp4_r_v_b_15')
// (9, 7, 'neigh_op_bot_7')
// (9, 7, 'sp4_r_v_b_2')
// (9, 8, 'sp4_r_v_b_40')
// (9, 9, 'sp4_r_v_b_29')
// (9, 10, 'sp4_r_v_b_16')
// (9, 11, 'sp4_h_r_40')
// (9, 11, 'sp4_r_v_b_5')
// (10, 3, 'sp4_v_t_39')
// (10, 4, 'sp4_v_b_39')
// (10, 5, 'neigh_op_tnl_7')
// (10, 5, 'sp4_v_b_26')
// (10, 6, 'neigh_op_lft_7')
// (10, 6, 'sp4_v_b_15')
// (10, 7, 'neigh_op_bnl_7')
// (10, 7, 'sp4_v_b_2')
// (10, 7, 'sp4_v_t_40')
// (10, 8, 'sp4_v_b_40')
// (10, 9, 'sp4_v_b_29')
// (10, 10, 'sp4_v_b_16')
// (10, 11, 'sp4_h_l_40')
// (10, 11, 'sp4_v_b_5')

wire n892;
// (6, 11, 'sp4_h_r_6')
// (7, 8, 'sp4_r_v_b_46')
// (7, 9, 'sp4_r_v_b_35')
// (7, 10, 'local_g3_6')
// (7, 10, 'lutff_5/in_0')
// (7, 10, 'sp4_r_v_b_22')
// (7, 11, 'local_g0_3')
// (7, 11, 'lutff_6/in_3')
// (7, 11, 'sp4_h_r_19')
// (7, 11, 'sp4_r_v_b_11')
// (8, 7, 'sp4_v_t_46')
// (8, 8, 'sp4_r_v_b_46')
// (8, 8, 'sp4_v_b_46')
// (8, 9, 'sp4_r_v_b_35')
// (8, 9, 'sp4_v_b_35')
// (8, 10, 'sp4_r_v_b_22')
// (8, 10, 'sp4_v_b_22')
// (8, 11, 'sp4_h_r_11')
// (8, 11, 'sp4_h_r_30')
// (8, 11, 'sp4_r_v_b_11')
// (8, 11, 'sp4_v_b_11')
// (9, 7, 'local_g0_3')
// (9, 7, 'lutff_1/in_2')
// (9, 7, 'sp4_h_r_11')
// (9, 7, 'sp4_v_t_46')
// (9, 8, 'sp4_v_b_46')
// (9, 9, 'sp4_v_b_35')
// (9, 10, 'sp4_v_b_22')
// (9, 11, 'sp4_h_r_22')
// (9, 11, 'sp4_h_r_43')
// (9, 11, 'sp4_h_r_6')
// (9, 11, 'sp4_v_b_11')
// (10, 7, 'sp4_h_r_22')
// (10, 10, 'neigh_op_tnr_7')
// (10, 11, 'neigh_op_rgt_7')
// (10, 11, 'sp4_h_l_43')
// (10, 11, 'sp4_h_r_19')
// (10, 11, 'sp4_h_r_3')
// (10, 11, 'sp4_h_r_35')
// (10, 12, 'neigh_op_bnr_7')
// (11, 7, 'sp4_h_r_35')
// (11, 10, 'local_g1_7')
// (11, 10, 'lutff_6/in_2')
// (11, 10, 'neigh_op_top_7')
// (11, 11, 'lutff_7/out')
// (11, 11, 'sp4_h_r_14')
// (11, 11, 'sp4_h_r_30')
// (11, 11, 'sp4_h_r_46')
// (11, 12, 'neigh_op_bot_7')
// (12, 7, 'sp4_h_r_46')
// (12, 10, 'neigh_op_tnl_7')
// (12, 11, 'neigh_op_lft_7')
// (12, 11, 'sp4_h_l_46')
// (12, 11, 'sp4_h_r_27')
// (12, 11, 'sp4_h_r_43')
// (12, 12, 'neigh_op_bnl_7')
// (13, 7, 'sp4_h_l_46')
// (13, 11, 'sp4_h_l_43')
// (13, 11, 'sp4_h_r_38')
// (14, 11, 'sp4_h_l_38')

reg n893 = 0;
// (6, 11, 'sp4_r_v_b_43')
// (6, 12, 'sp4_r_v_b_30')
// (6, 13, 'sp4_r_v_b_19')
// (6, 14, 'sp4_r_v_b_6')
// (7, 10, 'sp4_h_r_6')
// (7, 10, 'sp4_v_t_43')
// (7, 11, 'sp4_v_b_43')
// (7, 12, 'local_g2_6')
// (7, 12, 'lutff_7/in_3')
// (7, 12, 'sp4_v_b_30')
// (7, 13, 'sp4_v_b_19')
// (7, 14, 'sp4_v_b_6')
// (8, 10, 'sp4_h_r_19')
// (9, 10, 'sp4_h_r_30')
// (10, 6, 'neigh_op_tnr_2')
// (10, 7, 'neigh_op_rgt_2')
// (10, 7, 'sp4_r_v_b_36')
// (10, 8, 'neigh_op_bnr_2')
// (10, 8, 'sp4_r_v_b_25')
// (10, 9, 'sp4_r_v_b_12')
// (10, 10, 'sp4_h_r_43')
// (10, 10, 'sp4_r_v_b_1')
// (11, 6, 'neigh_op_top_2')
// (11, 6, 'sp4_v_t_36')
// (11, 7, 'lutff_2/out')
// (11, 7, 'sp4_v_b_36')
// (11, 8, 'neigh_op_bot_2')
// (11, 8, 'sp4_v_b_25')
// (11, 9, 'sp4_v_b_12')
// (11, 10, 'sp4_h_l_43')
// (11, 10, 'sp4_v_b_1')
// (12, 6, 'neigh_op_tnl_2')
// (12, 7, 'neigh_op_lft_2')
// (12, 8, 'neigh_op_bnl_2')

reg n894 = 0;
// (6, 12, 'neigh_op_tnr_0')
// (6, 13, 'neigh_op_rgt_0')
// (6, 14, 'neigh_op_bnr_0')
// (7, 12, 'local_g0_0')
// (7, 12, 'lutff_7/in_1')
// (7, 12, 'neigh_op_top_0')
// (7, 13, 'lutff_0/out')
// (7, 14, 'neigh_op_bot_0')
// (8, 12, 'neigh_op_tnl_0')
// (8, 13, 'neigh_op_lft_0')
// (8, 14, 'neigh_op_bnl_0')

reg n895 = 0;
// (6, 12, 'neigh_op_tnr_1')
// (6, 13, 'neigh_op_rgt_1')
// (6, 14, 'neigh_op_bnr_1')
// (7, 12, 'neigh_op_top_1')
// (7, 13, 'local_g2_1')
// (7, 13, 'lutff_1/out')
// (7, 13, 'lutff_4/in_3')
// (7, 14, 'neigh_op_bot_1')
// (8, 12, 'neigh_op_tnl_1')
// (8, 13, 'neigh_op_lft_1')
// (8, 14, 'neigh_op_bnl_1')

reg n896 = 0;
// (6, 12, 'neigh_op_tnr_2')
// (6, 13, 'neigh_op_rgt_2')
// (6, 14, 'neigh_op_bnr_2')
// (7, 12, 'neigh_op_top_2')
// (7, 13, 'lutff_2/out')
// (7, 14, 'neigh_op_bot_2')
// (8, 12, 'neigh_op_tnl_2')
// (8, 13, 'local_g0_2')
// (8, 13, 'lutff_4/in_2')
// (8, 13, 'neigh_op_lft_2')
// (8, 14, 'neigh_op_bnl_2')

reg n897 = 0;
// (6, 12, 'neigh_op_tnr_3')
// (6, 13, 'neigh_op_rgt_3')
// (6, 14, 'neigh_op_bnr_3')
// (7, 12, 'neigh_op_top_3')
// (7, 13, 'lutff_3/out')
// (7, 14, 'neigh_op_bot_3')
// (8, 12, 'neigh_op_tnl_3')
// (8, 13, 'local_g0_3')
// (8, 13, 'lutff_4/in_3')
// (8, 13, 'neigh_op_lft_3')
// (8, 14, 'neigh_op_bnl_3')

wire n898;
// (6, 12, 'neigh_op_tnr_4')
// (6, 12, 'sp4_r_v_b_37')
// (6, 13, 'neigh_op_rgt_4')
// (6, 13, 'sp4_r_v_b_24')
// (6, 14, 'neigh_op_bnr_4')
// (6, 14, 'sp4_r_v_b_13')
// (6, 15, 'sp4_r_v_b_0')
// (7, 11, 'sp4_h_r_5')
// (7, 11, 'sp4_v_t_37')
// (7, 12, 'neigh_op_top_4')
// (7, 12, 'sp4_v_b_37')
// (7, 13, 'lutff_4/out')
// (7, 13, 'sp4_v_b_24')
// (7, 14, 'neigh_op_bot_4')
// (7, 14, 'sp4_v_b_13')
// (7, 15, 'sp4_v_b_0')
// (8, 11, 'sp4_h_r_16')
// (8, 12, 'neigh_op_tnl_4')
// (8, 13, 'neigh_op_lft_4')
// (8, 14, 'neigh_op_bnl_4')
// (9, 11, 'local_g3_5')
// (9, 11, 'lutff_5/in_3')
// (9, 11, 'sp4_h_r_29')
// (10, 11, 'sp4_h_r_40')
// (11, 11, 'sp4_h_l_40')

reg n899 = 0;
// (6, 12, 'neigh_op_tnr_5')
// (6, 13, 'neigh_op_rgt_5')
// (6, 14, 'neigh_op_bnr_5')
// (7, 12, 'neigh_op_top_5')
// (7, 13, 'local_g3_5')
// (7, 13, 'lutff_4/in_2')
// (7, 13, 'lutff_5/out')
// (7, 14, 'neigh_op_bot_5')
// (8, 12, 'neigh_op_tnl_5')
// (8, 13, 'neigh_op_lft_5')
// (8, 14, 'neigh_op_bnl_5')

reg n900 = 0;
// (6, 12, 'neigh_op_tnr_6')
// (6, 13, 'neigh_op_rgt_6')
// (6, 14, 'neigh_op_bnr_6')
// (7, 12, 'neigh_op_top_6')
// (7, 13, 'local_g0_6')
// (7, 13, 'lutff_4/in_0')
// (7, 13, 'lutff_6/out')
// (7, 14, 'neigh_op_bot_6')
// (8, 12, 'neigh_op_tnl_6')
// (8, 13, 'neigh_op_lft_6')
// (8, 14, 'neigh_op_bnl_6')

reg n901 = 0;
// (6, 12, 'neigh_op_tnr_7')
// (6, 13, 'neigh_op_rgt_7')
// (6, 14, 'neigh_op_bnr_7')
// (7, 12, 'local_g0_7')
// (7, 12, 'lutff_7/in_0')
// (7, 12, 'neigh_op_top_7')
// (7, 13, 'lutff_7/out')
// (7, 14, 'neigh_op_bot_7')
// (8, 12, 'neigh_op_tnl_7')
// (8, 13, 'neigh_op_lft_7')
// (8, 14, 'neigh_op_bnl_7')

wire n902;
// (6, 12, 'sp4_h_r_1')
// (7, 12, 'local_g1_4')
// (7, 12, 'lutff_6/in_1')
// (7, 12, 'sp4_h_r_12')
// (8, 11, 'neigh_op_tnr_2')
// (8, 12, 'neigh_op_rgt_2')
// (8, 12, 'sp4_h_r_25')
// (8, 13, 'neigh_op_bnr_2')
// (9, 11, 'neigh_op_top_2')
// (9, 12, 'lutff_2/out')
// (9, 12, 'sp4_h_r_36')
// (9, 13, 'neigh_op_bot_2')
// (10, 11, 'neigh_op_tnl_2')
// (10, 12, 'neigh_op_lft_2')
// (10, 12, 'sp4_h_l_36')
// (10, 13, 'neigh_op_bnl_2')

reg n903 = 0;
// (6, 13, 'neigh_op_tnr_1')
// (6, 14, 'neigh_op_rgt_1')
// (6, 15, 'neigh_op_bnr_1')
// (7, 13, 'neigh_op_top_1')
// (7, 14, 'local_g2_1')
// (7, 14, 'lutff_0/in_1')
// (7, 14, 'lutff_1/out')
// (7, 14, 'lutff_6/in_1')
// (7, 15, 'neigh_op_bot_1')
// (8, 13, 'neigh_op_tnl_1')
// (8, 14, 'neigh_op_lft_1')
// (8, 15, 'neigh_op_bnl_1')

reg n904 = 0;
// (6, 13, 'neigh_op_tnr_2')
// (6, 14, 'neigh_op_rgt_2')
// (6, 14, 'sp4_h_r_9')
// (6, 15, 'neigh_op_bnr_2')
// (7, 13, 'neigh_op_top_2')
// (7, 14, 'local_g2_2')
// (7, 14, 'lutff_2/in_2')
// (7, 14, 'lutff_2/out')
// (7, 14, 'sp4_h_r_20')
// (7, 14, 'sp4_r_v_b_37')
// (7, 15, 'neigh_op_bot_2')
// (7, 15, 'sp4_r_v_b_24')
// (7, 16, 'sp4_r_v_b_13')
// (7, 17, 'sp4_r_v_b_0')
// (8, 13, 'neigh_op_tnl_2')
// (8, 13, 'sp4_h_r_0')
// (8, 13, 'sp4_v_t_37')
// (8, 14, 'neigh_op_lft_2')
// (8, 14, 'sp4_h_r_33')
// (8, 14, 'sp4_v_b_37')
// (8, 15, 'neigh_op_bnl_2')
// (8, 15, 'sp4_v_b_24')
// (8, 16, 'sp4_v_b_13')
// (8, 17, 'sp4_v_b_0')
// (9, 13, 'sp4_h_r_13')
// (9, 14, 'sp4_h_r_44')
// (10, 13, 'local_g2_0')
// (10, 13, 'lutff_5/in_3')
// (10, 13, 'sp4_h_r_24')
// (10, 14, 'sp4_h_l_44')
// (10, 14, 'sp4_h_r_9')
// (11, 13, 'sp4_h_r_37')
// (11, 14, 'local_g1_4')
// (11, 14, 'lutff_7/in_0')
// (11, 14, 'sp4_h_r_20')
// (12, 13, 'sp4_h_l_37')
// (12, 14, 'sp4_h_r_33')
// (13, 14, 'sp4_h_r_44')
// (14, 14, 'sp4_h_l_44')

reg n905 = 0;
// (6, 13, 'neigh_op_tnr_4')
// (6, 14, 'neigh_op_rgt_4')
// (6, 15, 'neigh_op_bnr_4')
// (7, 13, 'neigh_op_top_4')
// (7, 14, 'local_g0_4')
// (7, 14, 'lutff_0/in_2')
// (7, 14, 'lutff_4/out')
// (7, 14, 'lutff_6/in_2')
// (7, 15, 'neigh_op_bot_4')
// (8, 13, 'neigh_op_tnl_4')
// (8, 14, 'neigh_op_lft_4')
// (8, 15, 'neigh_op_bnl_4')

wire n906;
// (6, 13, 'neigh_op_tnr_6')
// (6, 14, 'neigh_op_rgt_6')
// (6, 15, 'neigh_op_bnr_6')
// (7, 13, 'neigh_op_top_6')
// (7, 14, 'local_g1_6')
// (7, 14, 'lutff_1/in_0')
// (7, 14, 'lutff_6/out')
// (7, 15, 'neigh_op_bot_6')
// (8, 13, 'neigh_op_tnl_6')
// (8, 14, 'neigh_op_lft_6')
// (8, 15, 'neigh_op_bnl_6')

reg n907 = 0;
// (6, 13, 'sp4_h_r_5')
// (7, 13, 'sp4_h_r_16')
// (8, 13, 'local_g3_5')
// (8, 13, 'lutff_6/in_0')
// (8, 13, 'sp4_h_r_29')
// (8, 20, 'neigh_op_tnr_4')
// (8, 21, 'neigh_op_rgt_4')
// (8, 22, 'neigh_op_bnr_4')
// (9, 6, 'sp4_r_v_b_45')
// (9, 7, 'sp4_r_v_b_32')
// (9, 8, 'sp4_r_v_b_21')
// (9, 9, 'local_g2_0')
// (9, 9, 'lutff_0/in_2')
// (9, 9, 'sp4_r_v_b_8')
// (9, 10, 'sp4_r_v_b_45')
// (9, 11, 'sp4_r_v_b_32')
// (9, 12, 'sp4_r_v_b_21')
// (9, 13, 'sp4_h_r_40')
// (9, 13, 'sp4_r_v_b_8')
// (9, 14, 'sp4_r_v_b_40')
// (9, 15, 'sp4_r_v_b_29')
// (9, 16, 'sp4_r_v_b_16')
// (9, 17, 'local_g1_5')
// (9, 17, 'lutff_7/in_3')
// (9, 17, 'sp4_r_v_b_5')
// (9, 18, 'sp4_r_v_b_44')
// (9, 19, 'local_g2_1')
// (9, 19, 'lutff_2/in_3')
// (9, 19, 'lutff_4/in_3')
// (9, 19, 'sp4_r_v_b_33')
// (9, 20, 'local_g0_4')
// (9, 20, 'lutff_7/in_1')
// (9, 20, 'neigh_op_top_4')
// (9, 20, 'sp4_r_v_b_20')
// (9, 21, 'lutff_4/out')
// (9, 21, 'sp4_r_v_b_9')
// (9, 22, 'local_g1_4')
// (9, 22, 'lutff_4/in_1')
// (9, 22, 'neigh_op_bot_4')
// (10, 5, 'sp4_v_t_45')
// (10, 6, 'sp4_v_b_45')
// (10, 7, 'sp4_v_b_32')
// (10, 8, 'sp4_v_b_21')
// (10, 9, 'sp4_v_b_8')
// (10, 9, 'sp4_v_t_45')
// (10, 10, 'sp4_v_b_45')
// (10, 11, 'sp4_v_b_32')
// (10, 12, 'sp4_v_b_21')
// (10, 13, 'sp4_h_l_40')
// (10, 13, 'sp4_v_b_8')
// (10, 13, 'sp4_v_t_40')
// (10, 14, 'sp4_v_b_40')
// (10, 15, 'sp4_v_b_29')
// (10, 16, 'sp4_v_b_16')
// (10, 17, 'sp4_v_b_5')
// (10, 17, 'sp4_v_t_44')
// (10, 18, 'sp4_v_b_44')
// (10, 19, 'local_g2_1')
// (10, 19, 'lutff_5/in_0')
// (10, 19, 'sp4_v_b_33')
// (10, 20, 'neigh_op_tnl_4')
// (10, 20, 'sp4_v_b_20')
// (10, 21, 'neigh_op_lft_4')
// (10, 21, 'sp4_v_b_9')
// (10, 22, 'neigh_op_bnl_4')

reg n908 = 0;
// (6, 13, 'sp4_h_r_7')
// (7, 13, 'local_g1_2')
// (7, 13, 'lutff_4/in_1')
// (7, 13, 'sp4_h_r_18')
// (8, 12, 'neigh_op_tnr_5')
// (8, 13, 'neigh_op_rgt_5')
// (8, 13, 'sp4_h_r_31')
// (8, 14, 'neigh_op_bnr_5')
// (9, 12, 'neigh_op_top_5')
// (9, 13, 'lutff_5/out')
// (9, 13, 'sp4_h_r_42')
// (9, 14, 'neigh_op_bot_5')
// (10, 12, 'neigh_op_tnl_5')
// (10, 13, 'neigh_op_lft_5')
// (10, 13, 'sp4_h_l_42')
// (10, 14, 'neigh_op_bnl_5')

wire n909;
// (6, 13, 'sp4_r_v_b_46')
// (6, 14, 'sp4_r_v_b_35')
// (6, 15, 'sp4_r_v_b_22')
// (6, 16, 'sp4_r_v_b_11')
// (6, 17, 'sp4_r_v_b_46')
// (6, 18, 'sp4_r_v_b_35')
// (6, 19, 'sp4_r_v_b_22')
// (6, 20, 'sp4_r_v_b_11')
// (7, 12, 'sp4_v_t_46')
// (7, 13, 'sp4_v_b_46')
// (7, 14, 'sp4_v_b_35')
// (7, 15, 'local_g1_6')
// (7, 15, 'lutff_5/in_2')
// (7, 15, 'sp4_v_b_22')
// (7, 16, 'sp4_v_b_11')
// (7, 16, 'sp4_v_t_46')
// (7, 17, 'sp4_v_b_46')
// (7, 18, 'sp4_v_b_35')
// (7, 19, 'sp4_v_b_22')
// (7, 20, 'local_g0_3')
// (7, 20, 'lutff_5/in_2')
// (7, 20, 'sp4_h_r_11')
// (7, 20, 'sp4_v_b_11')
// (8, 17, 'sp4_r_v_b_38')
// (8, 18, 'sp4_r_v_b_27')
// (8, 19, 'local_g2_6')
// (8, 19, 'lutff_5/in_1')
// (8, 19, 'sp4_r_v_b_14')
// (8, 20, 'sp4_h_r_22')
// (8, 20, 'sp4_r_v_b_3')
// (9, 14, 'sp4_r_v_b_43')
// (9, 15, 'sp4_r_v_b_30')
// (9, 16, 'local_g3_3')
// (9, 16, 'lutff_5/in_1')
// (9, 16, 'sp4_r_v_b_19')
// (9, 16, 'sp4_v_t_38')
// (9, 17, 'sp4_r_v_b_6')
// (9, 17, 'sp4_v_b_38')
// (9, 18, 'sp4_r_v_b_38')
// (9, 18, 'sp4_v_b_27')
// (9, 19, 'neigh_op_tnr_7')
// (9, 19, 'sp4_r_v_b_27')
// (9, 19, 'sp4_v_b_14')
// (9, 20, 'neigh_op_rgt_7')
// (9, 20, 'sp4_h_r_3')
// (9, 20, 'sp4_h_r_35')
// (9, 20, 'sp4_r_v_b_14')
// (9, 20, 'sp4_v_b_3')
// (9, 21, 'neigh_op_bnr_7')
// (9, 21, 'sp4_r_v_b_3')
// (10, 13, 'sp4_v_t_43')
// (10, 14, 'sp4_v_b_43')
// (10, 15, 'sp4_v_b_30')
// (10, 16, 'sp4_v_b_19')
// (10, 17, 'sp4_v_b_6')
// (10, 17, 'sp4_v_t_38')
// (10, 18, 'sp4_v_b_38')
// (10, 19, 'neigh_op_top_7')
// (10, 19, 'sp4_v_b_27')
// (10, 20, 'lutff_7/out')
// (10, 20, 'sp4_h_r_14')
// (10, 20, 'sp4_h_r_46')
// (10, 20, 'sp4_v_b_14')
// (10, 21, 'neigh_op_bot_7')
// (10, 21, 'sp4_v_b_3')
// (11, 19, 'neigh_op_tnl_7')
// (11, 20, 'neigh_op_lft_7')
// (11, 20, 'sp4_h_l_46')
// (11, 20, 'sp4_h_r_27')
// (11, 21, 'neigh_op_bnl_7')
// (12, 20, 'sp4_h_r_38')
// (13, 20, 'sp4_h_l_38')

reg n910 = 0;
// (6, 14, 'sp4_r_v_b_36')
// (6, 15, 'sp4_r_v_b_25')
// (6, 16, 'sp4_r_v_b_12')
// (6, 17, 'sp4_r_v_b_1')
// (7, 12, 'neigh_op_tnr_1')
// (7, 12, 'sp4_r_v_b_47')
// (7, 13, 'neigh_op_rgt_1')
// (7, 13, 'sp4_h_r_7')
// (7, 13, 'sp4_r_v_b_34')
// (7, 13, 'sp4_v_t_36')
// (7, 14, 'neigh_op_bnr_1')
// (7, 14, 'sp4_r_v_b_23')
// (7, 14, 'sp4_v_b_36')
// (7, 15, 'local_g3_1')
// (7, 15, 'lutff_1/in_1')
// (7, 15, 'sp4_r_v_b_10')
// (7, 15, 'sp4_v_b_25')
// (7, 16, 'sp4_v_b_12')
// (7, 17, 'sp4_v_b_1')
// (8, 11, 'sp4_v_t_47')
// (8, 12, 'neigh_op_top_1')
// (8, 12, 'sp4_v_b_47')
// (8, 13, 'lutff_1/out')
// (8, 13, 'sp4_h_r_18')
// (8, 13, 'sp4_v_b_34')
// (8, 14, 'local_g1_1')
// (8, 14, 'lutff_1/in_1')
// (8, 14, 'lutff_4/in_2')
// (8, 14, 'neigh_op_bot_1')
// (8, 14, 'sp4_v_b_23')
// (8, 15, 'local_g0_2')
// (8, 15, 'lutff_1/in_1')
// (8, 15, 'sp4_v_b_10')
// (9, 12, 'neigh_op_tnl_1')
// (9, 13, 'local_g0_1')
// (9, 13, 'lutff_0/in_1')
// (9, 13, 'neigh_op_lft_1')
// (9, 13, 'sp4_h_r_31')
// (9, 14, 'neigh_op_bnl_1')
// (10, 13, 'sp4_h_r_42')
// (11, 13, 'sp4_h_l_42')

wire n911;
// (6, 14, 'sp4_r_v_b_44')
// (6, 15, 'sp4_r_v_b_33')
// (6, 16, 'sp4_r_v_b_20')
// (6, 17, 'sp4_r_v_b_9')
// (6, 18, 'sp4_r_v_b_47')
// (6, 19, 'sp4_r_v_b_34')
// (6, 20, 'sp4_r_v_b_23')
// (6, 21, 'sp4_r_v_b_10')
// (7, 13, 'sp4_v_t_44')
// (7, 14, 'sp4_v_b_44')
// (7, 15, 'sp4_v_b_33')
// (7, 16, 'local_g0_4')
// (7, 16, 'lutff_0/in_2')
// (7, 16, 'sp4_v_b_20')
// (7, 17, 'sp4_h_r_4')
// (7, 17, 'sp4_v_b_9')
// (7, 17, 'sp4_v_t_47')
// (7, 18, 'sp4_v_b_47')
// (7, 19, 'sp4_v_b_34')
// (7, 20, 'sp4_v_b_23')
// (7, 21, 'local_g0_2')
// (7, 21, 'lutff_0/in_2')
// (7, 21, 'sp4_v_b_10')
// (8, 16, 'neigh_op_tnr_6')
// (8, 17, 'neigh_op_rgt_6')
// (8, 17, 'sp4_h_r_17')
// (8, 17, 'sp4_r_v_b_44')
// (8, 18, 'neigh_op_bnr_6')
// (8, 18, 'sp4_r_v_b_33')
// (8, 19, 'sp4_r_v_b_20')
// (8, 20, 'local_g2_1')
// (8, 20, 'lutff_0/in_1')
// (8, 20, 'sp4_r_v_b_9')
// (9, 16, 'neigh_op_top_6')
// (9, 16, 'sp4_v_t_44')
// (9, 17, 'local_g0_6')
// (9, 17, 'lutff_0/in_2')
// (9, 17, 'lutff_6/out')
// (9, 17, 'sp4_h_r_28')
// (9, 17, 'sp4_v_b_44')
// (9, 18, 'neigh_op_bot_6')
// (9, 18, 'sp4_v_b_33')
// (9, 19, 'sp4_v_b_20')
// (9, 20, 'sp4_v_b_9')
// (10, 16, 'neigh_op_tnl_6')
// (10, 17, 'neigh_op_lft_6')
// (10, 17, 'sp4_h_r_41')
// (10, 18, 'neigh_op_bnl_6')
// (11, 17, 'sp4_h_l_41')

wire n912;
// (6, 15, 'neigh_op_tnr_1')
// (6, 16, 'neigh_op_rgt_1')
// (6, 17, 'neigh_op_bnr_1')
// (7, 15, 'neigh_op_top_1')
// (7, 16, 'lutff_1/out')
// (7, 17, 'neigh_op_bot_1')
// (8, 15, 'neigh_op_tnl_1')
// (8, 16, 'local_g0_1')
// (8, 16, 'lutff_1/in_2')
// (8, 16, 'neigh_op_lft_1')
// (8, 17, 'neigh_op_bnl_1')

wire n913;
// (6, 15, 'neigh_op_tnr_2')
// (6, 16, 'neigh_op_rgt_2')
// (6, 16, 'sp4_h_r_9')
// (6, 16, 'sp4_r_v_b_36')
// (6, 17, 'neigh_op_bnr_2')
// (6, 17, 'sp4_r_v_b_25')
// (6, 18, 'sp4_r_v_b_12')
// (6, 19, 'sp4_r_v_b_1')
// (7, 15, 'neigh_op_top_2')
// (7, 15, 'sp4_v_t_36')
// (7, 16, 'lutff_2/out')
// (7, 16, 'sp4_h_r_20')
// (7, 16, 'sp4_v_b_36')
// (7, 17, 'neigh_op_bot_2')
// (7, 17, 'sp4_v_b_25')
// (7, 18, 'local_g1_4')
// (7, 18, 'lutff_6/in_1')
// (7, 18, 'sp4_v_b_12')
// (7, 19, 'sp4_v_b_1')
// (8, 15, 'local_g2_2')
// (8, 15, 'lutff_6/in_2')
// (8, 15, 'neigh_op_tnl_2')
// (8, 16, 'neigh_op_lft_2')
// (8, 16, 'sp4_h_r_33')
// (8, 17, 'local_g2_2')
// (8, 17, 'lutff_6/in_2')
// (8, 17, 'neigh_op_bnl_2')
// (9, 16, 'sp4_h_r_44')
// (9, 17, 'sp4_r_v_b_39')
// (9, 18, 'local_g0_2')
// (9, 18, 'lutff_6/in_2')
// (9, 18, 'sp4_r_v_b_26')
// (9, 19, 'sp4_r_v_b_15')
// (9, 20, 'sp4_r_v_b_2')
// (10, 16, 'sp4_h_l_44')
// (10, 16, 'sp4_v_t_39')
// (10, 17, 'sp4_v_b_39')
// (10, 18, 'sp4_v_b_26')
// (10, 19, 'sp4_v_b_15')
// (10, 20, 'sp4_v_b_2')

wire n914;
// (6, 16, 'neigh_op_tnr_0')
// (6, 17, 'neigh_op_rgt_0')
// (6, 18, 'neigh_op_bnr_0')
// (7, 15, 'sp4_r_v_b_41')
// (7, 16, 'neigh_op_top_0')
// (7, 16, 'sp4_r_v_b_28')
// (7, 17, 'lutff_0/out')
// (7, 17, 'sp4_r_v_b_17')
// (7, 18, 'local_g0_0')
// (7, 18, 'lutff_2/in_2')
// (7, 18, 'neigh_op_bot_0')
// (7, 18, 'sp4_r_v_b_4')
// (8, 14, 'sp4_v_t_41')
// (8, 15, 'local_g3_1')
// (8, 15, 'lutff_2/in_2')
// (8, 15, 'sp4_v_b_41')
// (8, 16, 'neigh_op_tnl_0')
// (8, 16, 'sp4_v_b_28')
// (8, 17, 'local_g1_0')
// (8, 17, 'lutff_2/in_1')
// (8, 17, 'neigh_op_lft_0')
// (8, 17, 'sp4_v_b_17')
// (8, 18, 'neigh_op_bnl_0')
// (8, 18, 'sp4_h_r_10')
// (8, 18, 'sp4_v_b_4')
// (9, 18, 'local_g0_7')
// (9, 18, 'lutff_2/in_1')
// (9, 18, 'sp4_h_r_23')
// (10, 18, 'sp4_h_r_34')
// (11, 18, 'sp4_h_r_47')
// (12, 18, 'sp4_h_l_47')

wire n915;
// (6, 16, 'neigh_op_tnr_3')
// (6, 17, 'neigh_op_rgt_3')
// (6, 18, 'neigh_op_bnr_3')
// (7, 14, 'sp4_r_v_b_42')
// (7, 15, 'sp4_r_v_b_31')
// (7, 15, 'sp4_r_v_b_47')
// (7, 16, 'neigh_op_top_3')
// (7, 16, 'sp4_r_v_b_18')
// (7, 16, 'sp4_r_v_b_34')
// (7, 17, 'lutff_3/out')
// (7, 17, 'sp4_r_v_b_23')
// (7, 17, 'sp4_r_v_b_7')
// (7, 18, 'local_g0_3')
// (7, 18, 'lutff_4/in_1')
// (7, 18, 'neigh_op_bot_3')
// (7, 18, 'sp4_r_v_b_10')
// (8, 13, 'sp4_v_t_42')
// (8, 14, 'sp4_v_b_42')
// (8, 14, 'sp4_v_t_47')
// (8, 15, 'local_g3_7')
// (8, 15, 'lutff_4/in_2')
// (8, 15, 'sp4_v_b_31')
// (8, 15, 'sp4_v_b_47')
// (8, 16, 'neigh_op_tnl_3')
// (8, 16, 'sp4_v_b_18')
// (8, 16, 'sp4_v_b_34')
// (8, 17, 'local_g1_3')
// (8, 17, 'lutff_4/in_2')
// (8, 17, 'neigh_op_lft_3')
// (8, 17, 'sp4_v_b_23')
// (8, 17, 'sp4_v_b_7')
// (8, 18, 'neigh_op_bnl_3')
// (8, 18, 'sp4_h_r_4')
// (8, 18, 'sp4_v_b_10')
// (9, 18, 'local_g1_1')
// (9, 18, 'lutff_4/in_2')
// (9, 18, 'sp4_h_r_17')
// (10, 18, 'sp4_h_r_28')
// (11, 18, 'sp4_h_r_41')
// (12, 18, 'sp4_h_l_41')

wire n916;
// (6, 16, 'neigh_op_tnr_5')
// (6, 17, 'neigh_op_rgt_5')
// (6, 18, 'neigh_op_bnr_5')
// (7, 16, 'neigh_op_top_5')
// (7, 17, 'local_g0_2')
// (7, 17, 'lutff_5/out')
// (7, 17, 'lutff_global/cen')
// (7, 17, 'sp4_h_r_10')
// (7, 18, 'neigh_op_bot_5')
// (8, 16, 'neigh_op_tnl_5')
// (8, 17, 'neigh_op_lft_5')
// (8, 17, 'sp4_h_r_23')
// (8, 18, 'neigh_op_bnl_5')
// (9, 17, 'sp4_h_r_34')
// (10, 17, 'sp4_h_r_47')
// (11, 17, 'sp4_h_l_47')

wire n917;
// (6, 16, 'neigh_op_tnr_6')
// (6, 17, 'neigh_op_rgt_6')
// (6, 18, 'neigh_op_bnr_6')
// (7, 15, 'sp4_r_v_b_37')
// (7, 16, 'neigh_op_top_6')
// (7, 16, 'sp4_r_v_b_24')
// (7, 17, 'lutff_6/out')
// (7, 17, 'sp4_r_v_b_13')
// (7, 18, 'local_g1_6')
// (7, 18, 'lutff_5/in_2')
// (7, 18, 'neigh_op_bot_6')
// (7, 18, 'sp4_r_v_b_0')
// (8, 14, 'sp4_v_t_37')
// (8, 15, 'local_g2_5')
// (8, 15, 'lutff_5/in_2')
// (8, 15, 'sp4_v_b_37')
// (8, 16, 'neigh_op_tnl_6')
// (8, 16, 'sp4_v_b_24')
// (8, 17, 'local_g1_6')
// (8, 17, 'lutff_5/in_2')
// (8, 17, 'neigh_op_lft_6')
// (8, 17, 'sp4_v_b_13')
// (8, 18, 'neigh_op_bnl_6')
// (8, 18, 'sp4_h_r_0')
// (8, 18, 'sp4_v_b_0')
// (9, 18, 'local_g0_5')
// (9, 18, 'lutff_5/in_2')
// (9, 18, 'sp4_h_r_13')
// (10, 18, 'sp4_h_r_24')
// (11, 18, 'sp4_h_r_37')
// (12, 18, 'sp4_h_l_37')

wire n918;
// (6, 16, 'neigh_op_tnr_7')
// (6, 17, 'neigh_op_rgt_7')
// (6, 18, 'neigh_op_bnr_7')
// (7, 15, 'sp4_r_v_b_39')
// (7, 16, 'neigh_op_top_7')
// (7, 16, 'sp4_r_v_b_26')
// (7, 17, 'lutff_7/out')
// (7, 17, 'sp4_r_v_b_15')
// (7, 18, 'local_g0_7')
// (7, 18, 'lutff_3/in_2')
// (7, 18, 'neigh_op_bot_7')
// (7, 18, 'sp4_r_v_b_2')
// (8, 14, 'sp4_v_t_39')
// (8, 15, 'local_g2_7')
// (8, 15, 'lutff_3/in_2')
// (8, 15, 'sp4_v_b_39')
// (8, 16, 'neigh_op_tnl_7')
// (8, 16, 'sp4_v_b_26')
// (8, 17, 'local_g0_7')
// (8, 17, 'lutff_3/in_2')
// (8, 17, 'neigh_op_lft_7')
// (8, 17, 'sp4_v_b_15')
// (8, 18, 'neigh_op_bnl_7')
// (8, 18, 'sp4_h_r_2')
// (8, 18, 'sp4_v_b_2')
// (9, 18, 'local_g1_7')
// (9, 18, 'lutff_3/in_1')
// (9, 18, 'sp4_h_r_15')
// (10, 18, 'sp4_h_r_26')
// (11, 18, 'sp4_h_r_39')
// (12, 18, 'sp4_h_l_39')

wire n919;
// (6, 17, 'sp4_r_v_b_38')
// (6, 18, 'sp4_r_v_b_27')
// (6, 19, 'sp4_r_v_b_14')
// (6, 20, 'sp4_r_v_b_3')
// (7, 15, 'local_g2_7')
// (7, 15, 'lutff_4/in_1')
// (7, 15, 'neigh_op_tnr_7')
// (7, 16, 'neigh_op_rgt_7')
// (7, 16, 'sp4_h_r_3')
// (7, 16, 'sp4_r_v_b_46')
// (7, 16, 'sp4_v_t_38')
// (7, 17, 'neigh_op_bnr_7')
// (7, 17, 'sp4_r_v_b_35')
// (7, 17, 'sp4_v_b_38')
// (7, 18, 'sp4_r_v_b_22')
// (7, 18, 'sp4_v_b_27')
// (7, 19, 'sp4_r_v_b_11')
// (7, 19, 'sp4_v_b_14')
// (7, 20, 'local_g1_3')
// (7, 20, 'lutff_4/in_2')
// (7, 20, 'sp4_v_b_3')
// (8, 15, 'neigh_op_top_7')
// (8, 15, 'sp4_v_t_46')
// (8, 16, 'lutff_7/out')
// (8, 16, 'sp4_h_r_14')
// (8, 16, 'sp4_v_b_46')
// (8, 17, 'neigh_op_bot_7')
// (8, 17, 'sp4_v_b_35')
// (8, 18, 'sp4_v_b_22')
// (8, 19, 'local_g0_3')
// (8, 19, 'lutff_4/in_1')
// (8, 19, 'sp4_v_b_11')
// (9, 15, 'neigh_op_tnl_7')
// (9, 16, 'local_g0_7')
// (9, 16, 'lutff_4/in_1')
// (9, 16, 'neigh_op_lft_7')
// (9, 16, 'sp4_h_r_27')
// (9, 17, 'neigh_op_bnl_7')
// (10, 16, 'sp4_h_r_38')
// (11, 16, 'sp4_h_l_38')

wire n920;
// (6, 17, 'sp4_r_v_b_40')
// (6, 18, 'sp4_r_v_b_29')
// (6, 19, 'sp4_r_v_b_16')
// (6, 20, 'sp4_r_v_b_5')
// (7, 15, 'local_g3_3')
// (7, 15, 'lutff_6/in_2')
// (7, 15, 'neigh_op_tnr_3')
// (7, 16, 'neigh_op_rgt_3')
// (7, 16, 'sp4_h_r_11')
// (7, 16, 'sp4_v_t_40')
// (7, 17, 'neigh_op_bnr_3')
// (7, 17, 'sp4_v_b_40')
// (7, 18, 'sp4_v_b_29')
// (7, 19, 'sp4_v_b_16')
// (7, 20, 'local_g0_5')
// (7, 20, 'lutff_6/in_1')
// (7, 20, 'sp4_v_b_5')
// (8, 15, 'neigh_op_top_3')
// (8, 16, 'lutff_3/out')
// (8, 16, 'sp4_h_r_22')
// (8, 16, 'sp4_r_v_b_39')
// (8, 17, 'neigh_op_bot_3')
// (8, 17, 'sp4_r_v_b_26')
// (8, 18, 'sp4_r_v_b_15')
// (8, 19, 'local_g1_2')
// (8, 19, 'lutff_6/in_1')
// (8, 19, 'sp4_r_v_b_2')
// (9, 15, 'neigh_op_tnl_3')
// (9, 15, 'sp4_v_t_39')
// (9, 16, 'local_g0_3')
// (9, 16, 'lutff_6/in_1')
// (9, 16, 'neigh_op_lft_3')
// (9, 16, 'sp4_h_r_35')
// (9, 16, 'sp4_v_b_39')
// (9, 17, 'neigh_op_bnl_3')
// (9, 17, 'sp4_v_b_26')
// (9, 18, 'sp4_v_b_15')
// (9, 19, 'sp4_v_b_2')
// (10, 16, 'sp4_h_r_46')
// (11, 16, 'sp4_h_l_46')

wire n921;
// (6, 17, 'sp4_r_v_b_42')
// (6, 18, 'sp4_r_v_b_31')
// (6, 19, 'sp4_r_v_b_18')
// (6, 20, 'sp4_r_v_b_7')
// (7, 15, 'local_g3_6')
// (7, 15, 'lutff_2/in_1')
// (7, 15, 'neigh_op_tnr_6')
// (7, 16, 'neigh_op_rgt_6')
// (7, 16, 'sp4_h_r_1')
// (7, 16, 'sp4_v_t_42')
// (7, 17, 'neigh_op_bnr_6')
// (7, 17, 'sp4_v_b_42')
// (7, 18, 'sp4_v_b_31')
// (7, 19, 'sp4_v_b_18')
// (7, 20, 'local_g1_7')
// (7, 20, 'lutff_2/in_2')
// (7, 20, 'sp4_v_b_7')
// (8, 15, 'neigh_op_top_6')
// (8, 16, 'lutff_6/out')
// (8, 16, 'sp4_h_r_12')
// (8, 16, 'sp4_r_v_b_45')
// (8, 17, 'neigh_op_bot_6')
// (8, 17, 'sp4_r_v_b_32')
// (8, 18, 'sp4_r_v_b_21')
// (8, 19, 'local_g2_0')
// (8, 19, 'lutff_2/in_2')
// (8, 19, 'sp4_r_v_b_8')
// (9, 15, 'neigh_op_tnl_6')
// (9, 15, 'sp4_v_t_45')
// (9, 16, 'local_g1_6')
// (9, 16, 'lutff_2/in_1')
// (9, 16, 'neigh_op_lft_6')
// (9, 16, 'sp4_h_r_25')
// (9, 16, 'sp4_v_b_45')
// (9, 17, 'neigh_op_bnl_6')
// (9, 17, 'sp4_v_b_32')
// (9, 18, 'sp4_v_b_21')
// (9, 19, 'sp4_v_b_8')
// (10, 16, 'sp4_h_r_36')
// (11, 16, 'sp4_h_l_36')

wire n922;
// (6, 17, 'sp4_r_v_b_44')
// (6, 18, 'sp4_r_v_b_33')
// (6, 19, 'sp4_r_v_b_20')
// (6, 20, 'sp4_r_v_b_9')
// (7, 15, 'local_g2_2')
// (7, 15, 'lutff_0/in_2')
// (7, 15, 'neigh_op_tnr_2')
// (7, 16, 'neigh_op_rgt_2')
// (7, 16, 'sp4_h_r_9')
// (7, 16, 'sp4_v_t_44')
// (7, 17, 'neigh_op_bnr_2')
// (7, 17, 'sp4_v_b_44')
// (7, 18, 'sp4_v_b_33')
// (7, 19, 'sp4_v_b_20')
// (7, 20, 'local_g0_1')
// (7, 20, 'lutff_0/in_1')
// (7, 20, 'sp4_v_b_9')
// (8, 15, 'neigh_op_top_2')
// (8, 16, 'lutff_2/out')
// (8, 16, 'sp4_h_r_20')
// (8, 16, 'sp4_r_v_b_37')
// (8, 17, 'neigh_op_bot_2')
// (8, 17, 'sp4_r_v_b_24')
// (8, 18, 'sp4_r_v_b_13')
// (8, 19, 'local_g1_0')
// (8, 19, 'lutff_0/in_1')
// (8, 19, 'sp4_r_v_b_0')
// (9, 15, 'neigh_op_tnl_2')
// (9, 15, 'sp4_v_t_37')
// (9, 16, 'local_g1_2')
// (9, 16, 'lutff_0/in_1')
// (9, 16, 'neigh_op_lft_2')
// (9, 16, 'sp4_h_r_33')
// (9, 16, 'sp4_v_b_37')
// (9, 17, 'neigh_op_bnl_2')
// (9, 17, 'sp4_v_b_24')
// (9, 18, 'sp4_v_b_13')
// (9, 19, 'sp4_v_b_0')
// (10, 16, 'sp4_h_r_44')
// (11, 16, 'sp4_h_l_44')

wire n923;
// (6, 18, 'neigh_op_tnr_4')
// (6, 19, 'neigh_op_rgt_4')
// (6, 20, 'neigh_op_bnr_4')
// (7, 16, 'sp4_r_v_b_44')
// (7, 17, 'sp4_r_v_b_33')
// (7, 18, 'neigh_op_top_4')
// (7, 18, 'sp4_r_v_b_20')
// (7, 19, 'local_g1_4')
// (7, 19, 'lutff_0/in_1')
// (7, 19, 'lutff_4/out')
// (7, 19, 'sp4_h_r_8')
// (7, 19, 'sp4_r_v_b_9')
// (7, 20, 'neigh_op_bot_4')
// (8, 15, 'sp4_v_t_44')
// (8, 16, 'local_g3_4')
// (8, 16, 'lutff_0/in_1')
// (8, 16, 'sp4_v_b_44')
// (8, 17, 'sp4_v_b_33')
// (8, 18, 'local_g2_4')
// (8, 18, 'lutff_0/in_2')
// (8, 18, 'neigh_op_tnl_4')
// (8, 18, 'sp4_v_b_20')
// (8, 19, 'neigh_op_lft_4')
// (8, 19, 'sp4_h_r_21')
// (8, 19, 'sp4_v_b_9')
// (8, 20, 'neigh_op_bnl_4')
// (9, 19, 'local_g2_0')
// (9, 19, 'lutff_0/in_2')
// (9, 19, 'sp4_h_r_32')
// (10, 19, 'sp4_h_r_45')
// (11, 19, 'sp4_h_l_45')

wire n924;
// (6, 20, 'neigh_op_tnr_1')
// (6, 21, 'neigh_op_rgt_1')
// (6, 22, 'neigh_op_bnr_1')
// (7, 19, 'sp4_r_v_b_43')
// (7, 20, 'neigh_op_top_1')
// (7, 20, 'sp4_r_v_b_30')
// (7, 21, 'lutff_1/out')
// (7, 21, 'sp4_h_r_2')
// (7, 21, 'sp4_r_v_b_19')
// (7, 22, 'neigh_op_bot_1')
// (7, 22, 'sp4_r_v_b_6')
// (8, 18, 'sp4_v_t_43')
// (8, 19, 'sp4_v_b_43')
// (8, 20, 'neigh_op_tnl_1')
// (8, 20, 'sp4_v_b_30')
// (8, 21, 'local_g1_1')
// (8, 21, 'lutff_0/in_0')
// (8, 21, 'lutff_2/in_0')
// (8, 21, 'neigh_op_lft_1')
// (8, 21, 'sp4_h_r_15')
// (8, 21, 'sp4_v_b_19')
// (8, 22, 'local_g2_1')
// (8, 22, 'lutff_0/in_3')
// (8, 22, 'lutff_3/in_0')
// (8, 22, 'lutff_7/in_2')
// (8, 22, 'neigh_op_bnl_1')
// (8, 22, 'sp4_h_r_0')
// (8, 22, 'sp4_v_b_6')
// (9, 21, 'local_g2_2')
// (9, 21, 'lutff_2/in_2')
// (9, 21, 'lutff_3/in_3')
// (9, 21, 'lutff_6/in_0')
// (9, 21, 'sp4_h_r_26')
// (9, 22, 'local_g0_5')
// (9, 22, 'local_g1_5')
// (9, 22, 'lutff_6/in_1')
// (9, 22, 'lutff_7/in_1')
// (9, 22, 'sp4_h_r_13')
// (10, 21, 'sp4_h_r_39')
// (10, 22, 'sp4_h_r_24')
// (11, 21, 'sp4_h_l_39')
// (11, 22, 'sp4_h_r_37')
// (12, 22, 'sp4_h_l_37')

wire n925;
// (6, 20, 'neigh_op_tnr_2')
// (6, 21, 'neigh_op_rgt_2')
// (6, 22, 'neigh_op_bnr_2')
// (7, 20, 'neigh_op_top_2')
// (7, 21, 'lutff_2/out')
// (7, 22, 'neigh_op_bot_2')
// (8, 20, 'local_g3_2')
// (8, 20, 'lutff_2/in_3')
// (8, 20, 'lutff_3/in_2')
// (8, 20, 'lutff_4/in_3')
// (8, 20, 'lutff_5/in_0')
// (8, 20, 'neigh_op_tnl_2')
// (8, 21, 'local_g0_2')
// (8, 21, 'local_g1_2')
// (8, 21, 'lutff_3/in_0')
// (8, 21, 'lutff_6/in_0')
// (8, 21, 'neigh_op_lft_2')
// (8, 22, 'neigh_op_bnl_2')

wire n926;
// (6, 20, 'neigh_op_tnr_3')
// (6, 21, 'neigh_op_rgt_3')
// (6, 22, 'neigh_op_bnr_3')
// (7, 20, 'neigh_op_top_3')
// (7, 21, 'lutff_3/out')
// (7, 21, 'sp4_r_v_b_39')
// (7, 22, 'neigh_op_bot_3')
// (7, 22, 'sp4_r_v_b_26')
// (7, 23, 'sp4_r_v_b_15')
// (7, 24, 'sp4_r_v_b_2')
// (8, 20, 'neigh_op_tnl_3')
// (8, 20, 'sp4_v_t_39')
// (8, 21, 'local_g3_7')
// (8, 21, 'lutff_1/in_1')
// (8, 21, 'neigh_op_lft_3')
// (8, 21, 'sp4_v_b_39')
// (8, 22, 'neigh_op_bnl_3')
// (8, 22, 'sp4_v_b_26')
// (8, 23, 'sp4_v_b_15')
// (8, 24, 'sp4_v_b_2')

wire n927;
// (6, 20, 'neigh_op_tnr_5')
// (6, 21, 'neigh_op_rgt_5')
// (6, 22, 'neigh_op_bnr_5')
// (7, 20, 'neigh_op_top_5')
// (7, 21, 'local_g0_5')
// (7, 21, 'lutff_4/in_3')
// (7, 21, 'lutff_5/out')
// (7, 22, 'neigh_op_bot_5')
// (8, 20, 'neigh_op_tnl_5')
// (8, 21, 'neigh_op_lft_5')
// (8, 22, 'neigh_op_bnl_5')

wire n928;
// (6, 20, 'neigh_op_tnr_6')
// (6, 21, 'neigh_op_rgt_6')
// (6, 22, 'neigh_op_bnr_6')
// (7, 20, 'neigh_op_top_6')
// (7, 21, 'lutff_6/out')
// (7, 22, 'neigh_op_bot_6')
// (8, 20, 'neigh_op_tnl_6')
// (8, 21, 'local_g0_6')
// (8, 21, 'lutff_7/in_3')
// (8, 21, 'neigh_op_lft_6')
// (8, 22, 'neigh_op_bnl_6')

wire n929;
// (6, 20, 'neigh_op_tnr_7')
// (6, 21, 'neigh_op_rgt_7')
// (6, 21, 'sp4_h_r_3')
// (6, 22, 'neigh_op_bnr_7')
// (7, 20, 'neigh_op_top_7')
// (7, 21, 'lutff_7/out')
// (7, 21, 'sp4_h_r_14')
// (7, 22, 'neigh_op_bot_7')
// (8, 20, 'neigh_op_tnl_7')
// (8, 21, 'local_g2_3')
// (8, 21, 'lutff_5/in_2')
// (8, 21, 'neigh_op_lft_7')
// (8, 21, 'sp4_h_r_27')
// (8, 22, 'neigh_op_bnl_7')
// (9, 21, 'sp4_h_r_38')
// (10, 21, 'sp4_h_l_38')

wire n930;
// (6, 20, 'sp4_h_r_9')
// (7, 20, 'sp4_h_r_20')
// (8, 20, 'local_g3_1')
// (8, 20, 'lutff_4/in_0')
// (8, 20, 'sp4_h_r_33')
// (9, 17, 'sp4_r_v_b_44')
// (9, 18, 'neigh_op_tnr_2')
// (9, 18, 'sp4_r_v_b_33')
// (9, 19, 'neigh_op_rgt_2')
// (9, 19, 'sp4_r_v_b_20')
// (9, 20, 'neigh_op_bnr_2')
// (9, 20, 'sp4_h_r_44')
// (9, 20, 'sp4_r_v_b_9')
// (10, 16, 'sp4_v_t_44')
// (10, 17, 'sp4_v_b_44')
// (10, 18, 'neigh_op_top_2')
// (10, 18, 'sp4_v_b_33')
// (10, 19, 'local_g3_2')
// (10, 19, 'lutff_2/out')
// (10, 19, 'lutff_3/in_0')
// (10, 19, 'sp4_v_b_20')
// (10, 20, 'neigh_op_bot_2')
// (10, 20, 'sp4_h_l_44')
// (10, 20, 'sp4_v_b_9')
// (11, 18, 'neigh_op_tnl_2')
// (11, 19, 'neigh_op_lft_2')
// (11, 20, 'neigh_op_bnl_2')

reg n931 = 0;
// (6, 21, 'sp4_h_r_10')
// (7, 14, 'sp4_r_v_b_39')
// (7, 15, 'sp4_r_v_b_26')
// (7, 16, 'sp4_r_v_b_15')
// (7, 17, 'sp4_r_v_b_2')
// (7, 18, 'sp4_r_v_b_39')
// (7, 19, 'sp4_r_v_b_26')
// (7, 20, 'neigh_op_tnr_1')
// (7, 20, 'sp4_r_v_b_15')
// (7, 21, 'neigh_op_rgt_1')
// (7, 21, 'sp4_h_r_23')
// (7, 21, 'sp4_r_v_b_2')
// (7, 22, 'neigh_op_bnr_1')
// (8, 10, 'sp12_h_r_1')
// (8, 10, 'sp12_v_t_22')
// (8, 11, 'sp12_v_b_22')
// (8, 12, 'sp12_v_b_21')
// (8, 13, 'sp12_v_b_18')
// (8, 13, 'sp4_v_t_39')
// (8, 14, 'local_g3_7')
// (8, 14, 'lutff_6/in_0')
// (8, 14, 'sp12_v_b_17')
// (8, 14, 'sp4_v_b_39')
// (8, 15, 'sp12_v_b_14')
// (8, 15, 'sp4_v_b_26')
// (8, 16, 'local_g0_7')
// (8, 16, 'lutff_3/in_2')
// (8, 16, 'sp12_v_b_13')
// (8, 16, 'sp4_v_b_15')
// (8, 17, 'sp12_v_b_10')
// (8, 17, 'sp4_v_b_2')
// (8, 17, 'sp4_v_t_39')
// (8, 18, 'sp12_v_b_9')
// (8, 18, 'sp4_r_v_b_38')
// (8, 18, 'sp4_v_b_39')
// (8, 19, 'sp12_v_b_6')
// (8, 19, 'sp4_r_v_b_27')
// (8, 19, 'sp4_v_b_26')
// (8, 20, 'neigh_op_top_1')
// (8, 20, 'sp12_v_b_5')
// (8, 20, 'sp4_r_v_b_14')
// (8, 20, 'sp4_v_b_15')
// (8, 21, 'lutff_1/out')
// (8, 21, 'sp12_v_b_2')
// (8, 21, 'sp4_h_r_34')
// (8, 21, 'sp4_r_v_b_3')
// (8, 21, 'sp4_v_b_2')
// (8, 22, 'neigh_op_bot_1')
// (8, 22, 'sp12_v_b_1')
// (9, 10, 'sp12_h_r_2')
// (9, 17, 'sp4_v_t_38')
// (9, 18, 'sp4_r_v_b_47')
// (9, 18, 'sp4_v_b_38')
// (9, 19, 'local_g3_3')
// (9, 19, 'lutff_2/in_2')
// (9, 19, 'lutff_7/in_1')
// (9, 19, 'sp4_r_v_b_34')
// (9, 19, 'sp4_v_b_27')
// (9, 20, 'local_g3_1')
// (9, 20, 'lutff_6/in_2')
// (9, 20, 'neigh_op_tnl_1')
// (9, 20, 'sp4_r_v_b_23')
// (9, 20, 'sp4_v_b_14')
// (9, 21, 'neigh_op_lft_1')
// (9, 21, 'sp4_h_r_47')
// (9, 21, 'sp4_r_v_b_10')
// (9, 21, 'sp4_v_b_3')
// (9, 22, 'local_g2_1')
// (9, 22, 'lutff_3/in_2')
// (9, 22, 'neigh_op_bnl_1')
// (10, 10, 'local_g0_5')
// (10, 10, 'lutff_6/in_1')
// (10, 10, 'sp12_h_r_5')
// (10, 17, 'sp4_v_t_47')
// (10, 18, 'sp4_v_b_47')
// (10, 19, 'local_g2_2')
// (10, 19, 'lutff_4/in_0')
// (10, 19, 'sp4_v_b_34')
// (10, 20, 'sp4_v_b_23')
// (10, 21, 'sp4_h_l_47')
// (10, 21, 'sp4_v_b_10')
// (11, 10, 'sp12_h_r_6')
// (12, 10, 'sp12_h_r_9')
// (13, 10, 'sp12_h_r_10')
// (14, 10, 'sp12_h_r_13')
// (15, 10, 'sp12_h_r_14')
// (16, 10, 'sp12_h_r_17')
// (17, 10, 'sp12_h_r_18')
// (18, 10, 'sp12_h_r_21')
// (19, 10, 'sp12_h_r_22')
// (20, 10, 'sp12_h_l_22')

reg n932 = 0;
// (6, 21, 'sp4_h_r_4')
// (7, 20, 'neigh_op_tnr_6')
// (7, 20, 'sp4_r_v_b_41')
// (7, 21, 'neigh_op_rgt_6')
// (7, 21, 'sp4_h_r_17')
// (7, 21, 'sp4_r_v_b_28')
// (7, 22, 'neigh_op_bnr_6')
// (7, 22, 'sp4_r_v_b_17')
// (7, 23, 'sp4_r_v_b_4')
// (8, 11, 'sp4_r_v_b_46')
// (8, 12, 'sp4_r_v_b_35')
// (8, 13, 'sp4_r_v_b_22')
// (8, 14, 'local_g2_3')
// (8, 14, 'lutff_7/in_0')
// (8, 14, 'sp4_r_v_b_11')
// (8, 15, 'sp4_r_v_b_45')
// (8, 16, 'sp4_r_v_b_32')
// (8, 17, 'sp4_r_v_b_21')
// (8, 18, 'sp4_r_v_b_8')
// (8, 19, 'sp4_h_r_4')
// (8, 19, 'sp4_r_v_b_37')
// (8, 19, 'sp4_v_t_41')
// (8, 20, 'neigh_op_top_6')
// (8, 20, 'sp4_r_v_b_24')
// (8, 20, 'sp4_v_b_41')
// (8, 21, 'lutff_6/out')
// (8, 21, 'sp4_h_r_28')
// (8, 21, 'sp4_r_v_b_13')
// (8, 21, 'sp4_v_b_28')
// (8, 22, 'neigh_op_bot_6')
// (8, 22, 'sp4_r_v_b_0')
// (8, 22, 'sp4_v_b_17')
// (8, 23, 'sp4_v_b_4')
// (9, 10, 'sp4_v_t_46')
// (9, 11, 'sp4_v_b_46')
// (9, 12, 'sp4_v_b_35')
// (9, 13, 'sp4_v_b_22')
// (9, 14, 'sp4_v_b_11')
// (9, 14, 'sp4_v_t_45')
// (9, 15, 'sp4_v_b_45')
// (9, 16, 'sp4_v_b_32')
// (9, 17, 'local_g0_5')
// (9, 17, 'lutff_6/in_1')
// (9, 17, 'sp4_v_b_21')
// (9, 18, 'sp4_v_b_8')
// (9, 18, 'sp4_v_t_37')
// (9, 19, 'local_g2_5')
// (9, 19, 'lutff_2/in_1')
// (9, 19, 'lutff_7/in_0')
// (9, 19, 'sp4_h_r_17')
// (9, 19, 'sp4_v_b_37')
// (9, 20, 'neigh_op_tnl_6')
// (9, 20, 'sp4_v_b_24')
// (9, 21, 'local_g3_1')
// (9, 21, 'lutff_0/in_2')
// (9, 21, 'neigh_op_lft_6')
// (9, 21, 'sp4_h_r_41')
// (9, 21, 'sp4_v_b_13')
// (9, 22, 'local_g2_6')
// (9, 22, 'lutff_5/in_1')
// (9, 22, 'neigh_op_bnl_6')
// (9, 22, 'sp4_v_b_0')
// (10, 19, 'local_g2_4')
// (10, 19, 'lutff_1/in_3')
// (10, 19, 'sp4_h_r_28')
// (10, 21, 'sp4_h_l_41')
// (11, 19, 'sp4_h_r_41')
// (12, 19, 'sp4_h_l_41')

reg n933 = 0;
// (7, 0, 'logic_op_tnr_0')
// (7, 1, 'neigh_op_rgt_0')
// (7, 2, 'neigh_op_bnr_0')
// (8, 0, 'logic_op_top_0')
// (8, 1, 'local_g3_0')
// (8, 1, 'lutff_0/out')
// (8, 1, 'lutff_6/in_1')
// (8, 2, 'neigh_op_bot_0')
// (9, 0, 'logic_op_tnl_0')
// (9, 1, 'neigh_op_lft_0')
// (9, 2, 'neigh_op_bnl_0')

wire n934;
// (7, 0, 'logic_op_tnr_1')
// (7, 1, 'neigh_op_rgt_1')
// (7, 2, 'neigh_op_bnr_1')
// (8, 0, 'logic_op_top_1')
// (8, 1, 'lutff_1/out')
// (8, 2, 'local_g1_1')
// (8, 2, 'lutff_2/in_0')
// (8, 2, 'neigh_op_bot_1')
// (9, 0, 'logic_op_tnl_1')
// (9, 1, 'neigh_op_lft_1')
// (9, 2, 'neigh_op_bnl_1')

reg n935 = 0;
// (7, 0, 'logic_op_tnr_2')
// (7, 1, 'local_g2_2')
// (7, 1, 'lutff_2/in_0')
// (7, 1, 'neigh_op_rgt_2')
// (7, 2, 'neigh_op_bnr_2')
// (8, 0, 'logic_op_top_2')
// (8, 1, 'lutff_2/out')
// (8, 2, 'neigh_op_bot_2')
// (9, 0, 'logic_op_tnl_2')
// (9, 1, 'neigh_op_lft_2')
// (9, 2, 'neigh_op_bnl_2')

wire n936;
// (7, 0, 'logic_op_tnr_3')
// (7, 1, 'neigh_op_rgt_3')
// (7, 2, 'neigh_op_bnr_3')
// (8, 0, 'logic_op_top_3')
// (8, 1, 'lutff_3/out')
// (8, 2, 'local_g0_3')
// (8, 2, 'lutff_6/in_3')
// (8, 2, 'neigh_op_bot_3')
// (9, 0, 'logic_op_tnl_3')
// (9, 1, 'neigh_op_lft_3')
// (9, 2, 'neigh_op_bnl_3')

reg n937 = 0;
// (7, 0, 'logic_op_tnr_4')
// (7, 1, 'local_g2_4')
// (7, 1, 'lutff_2/in_2')
// (7, 1, 'neigh_op_rgt_4')
// (7, 2, 'neigh_op_bnr_4')
// (8, 0, 'logic_op_top_4')
// (8, 1, 'lutff_4/out')
// (8, 2, 'neigh_op_bot_4')
// (9, 0, 'logic_op_tnl_4')
// (9, 1, 'neigh_op_lft_4')
// (9, 2, 'neigh_op_bnl_4')

reg n938 = 0;
// (7, 0, 'logic_op_tnr_5')
// (7, 1, 'neigh_op_rgt_5')
// (7, 2, 'neigh_op_bnr_5')
// (8, 0, 'logic_op_top_5')
// (8, 1, 'local_g1_5')
// (8, 1, 'lutff_5/out')
// (8, 1, 'lutff_6/in_2')
// (8, 2, 'neigh_op_bot_5')
// (9, 0, 'logic_op_tnl_5')
// (9, 1, 'neigh_op_lft_5')
// (9, 2, 'neigh_op_bnl_5')

wire n939;
// (7, 0, 'logic_op_tnr_6')
// (7, 1, 'neigh_op_rgt_6')
// (7, 2, 'local_g0_6')
// (7, 2, 'lutff_0/in_2')
// (7, 2, 'neigh_op_bnr_6')
// (8, 0, 'logic_op_top_6')
// (8, 1, 'lutff_6/out')
// (8, 2, 'neigh_op_bot_6')
// (9, 0, 'logic_op_tnl_6')
// (9, 1, 'neigh_op_lft_6')
// (9, 2, 'neigh_op_bnl_6')

wire n940;
// (7, 0, 'logic_op_tnr_7')
// (7, 1, 'neigh_op_rgt_7')
// (7, 2, 'local_g0_7')
// (7, 2, 'lutff_1/in_2')
// (7, 2, 'neigh_op_bnr_7')
// (8, 0, 'logic_op_top_7')
// (8, 1, 'lutff_7/out')
// (8, 2, 'neigh_op_bot_7')
// (9, 0, 'logic_op_tnl_7')
// (9, 1, 'neigh_op_lft_7')
// (9, 2, 'neigh_op_bnl_7')

wire n941;
// (7, 1, 'neigh_op_tnr_1')
// (7, 2, 'neigh_op_rgt_1')
// (7, 3, 'neigh_op_bnr_1')
// (8, 1, 'neigh_op_top_1')
// (8, 2, 'local_g0_2')
// (8, 2, 'lutff_1/out')
// (8, 2, 'lutff_6/in_0')
// (8, 2, 'sp4_h_r_2')
// (8, 3, 'neigh_op_bot_1')
// (9, 1, 'neigh_op_tnl_1')
// (9, 2, 'neigh_op_lft_1')
// (9, 2, 'sp4_h_r_15')
// (9, 3, 'neigh_op_bnl_1')
// (10, 2, 'sp4_h_r_26')
// (11, 2, 'sp4_h_r_39')
// (12, 2, 'sp4_h_l_39')

wire n942;
// (7, 1, 'neigh_op_tnr_2')
// (7, 2, 'local_g2_2')
// (7, 2, 'lutff_4/in_0')
// (7, 2, 'neigh_op_rgt_2')
// (7, 3, 'local_g0_2')
// (7, 3, 'lutff_6/in_2')
// (7, 3, 'neigh_op_bnr_2')
// (8, 1, 'neigh_op_top_2')
// (8, 2, 'lutff_2/out')
// (8, 3, 'neigh_op_bot_2')
// (9, 1, 'neigh_op_tnl_2')
// (9, 2, 'neigh_op_lft_2')
// (9, 3, 'neigh_op_bnl_2')

wire n943;
// (7, 1, 'neigh_op_tnr_3')
// (7, 2, 'local_g2_3')
// (7, 2, 'lutff_5/in_0')
// (7, 2, 'neigh_op_rgt_3')
// (7, 3, 'neigh_op_bnr_3')
// (8, 1, 'neigh_op_top_3')
// (8, 1, 'sp4_r_v_b_18')
// (8, 2, 'local_g1_7')
// (8, 2, 'lutff_1/in_3')
// (8, 2, 'lutff_3/out')
// (8, 2, 'sp4_r_v_b_7')
// (8, 3, 'neigh_op_bot_3')
// (9, 0, 'span4_vert_18')
// (9, 1, 'neigh_op_tnl_3')
// (9, 1, 'sp4_v_b_18')
// (9, 2, 'neigh_op_lft_3')
// (9, 2, 'sp4_v_b_7')
// (9, 3, 'neigh_op_bnl_3')

reg n944 = 0;
// (7, 1, 'neigh_op_tnr_4')
// (7, 2, 'neigh_op_rgt_4')
// (7, 2, 'sp4_r_v_b_40')
// (7, 3, 'neigh_op_bnr_4')
// (7, 3, 'sp4_r_v_b_29')
// (7, 4, 'sp4_r_v_b_16')
// (7, 5, 'sp4_r_v_b_5')
// (8, 1, 'neigh_op_top_4')
// (8, 1, 'sp4_v_t_40')
// (8, 2, 'local_g3_4')
// (8, 2, 'lutff_4/out')
// (8, 2, 'lutff_5/in_0')
// (8, 2, 'sp4_v_b_40')
// (8, 3, 'neigh_op_bot_4')
// (8, 3, 'sp4_v_b_29')
// (8, 4, 'local_g1_0')
// (8, 4, 'lutff_1/in_2')
// (8, 4, 'sp4_v_b_16')
// (8, 5, 'sp4_v_b_5')
// (9, 1, 'neigh_op_tnl_4')
// (9, 2, 'neigh_op_lft_4')
// (9, 3, 'neigh_op_bnl_4')

wire n945;
// (7, 1, 'neigh_op_tnr_5')
// (7, 2, 'neigh_op_rgt_5')
// (7, 3, 'neigh_op_bnr_5')
// (8, 1, 'neigh_op_top_5')
// (8, 2, 'local_g1_5')
// (8, 2, 'lutff_3/in_1')
// (8, 2, 'lutff_5/out')
// (8, 3, 'neigh_op_bot_5')
// (9, 1, 'neigh_op_tnl_5')
// (9, 2, 'neigh_op_lft_5')
// (9, 3, 'neigh_op_bnl_5')

wire n946;
// (7, 1, 'neigh_op_tnr_7')
// (7, 2, 'neigh_op_rgt_7')
// (7, 3, 'neigh_op_bnr_7')
// (8, 1, 'neigh_op_top_7')
// (8, 2, 'lutff_7/out')
// (8, 3, 'local_g0_7')
// (8, 3, 'lutff_4/in_3')
// (8, 3, 'neigh_op_bot_7')
// (9, 1, 'neigh_op_tnl_7')
// (9, 2, 'neigh_op_lft_7')
// (9, 3, 'neigh_op_bnl_7')

wire n947;
// (7, 1, 'sp4_r_v_b_47')
// (7, 2, 'sp4_r_v_b_34')
// (7, 3, 'neigh_op_tnr_5')
// (7, 3, 'sp4_r_v_b_23')
// (7, 4, 'neigh_op_rgt_5')
// (7, 4, 'sp4_r_v_b_10')
// (7, 5, 'neigh_op_bnr_5')
// (8, 0, 'span4_vert_47')
// (8, 1, 'sp4_v_b_47')
// (8, 2, 'local_g3_2')
// (8, 2, 'lutff_7/in_2')
// (8, 2, 'sp4_v_b_34')
// (8, 3, 'neigh_op_top_5')
// (8, 3, 'sp4_v_b_23')
// (8, 4, 'lutff_5/out')
// (8, 4, 'sp4_v_b_10')
// (8, 5, 'neigh_op_bot_5')
// (9, 3, 'neigh_op_tnl_5')
// (9, 4, 'neigh_op_lft_5')
// (9, 5, 'neigh_op_bnl_5')

wire n948;
// (7, 2, 'local_g3_0')
// (7, 2, 'lutff_4/in_1')
// (7, 2, 'neigh_op_tnr_0')
// (7, 3, 'local_g2_0')
// (7, 3, 'lutff_6/in_0')
// (7, 3, 'neigh_op_rgt_0')
// (7, 4, 'neigh_op_bnr_0')
// (8, 2, 'neigh_op_top_0')
// (8, 3, 'lutff_0/out')
// (8, 4, 'neigh_op_bot_0')
// (9, 2, 'neigh_op_tnl_0')
// (9, 3, 'neigh_op_lft_0')
// (9, 4, 'neigh_op_bnl_0')

wire n949;
// (7, 2, 'local_g3_1')
// (7, 2, 'lutff_5/in_3')
// (7, 2, 'neigh_op_tnr_1')
// (7, 3, 'neigh_op_rgt_1')
// (7, 4, 'neigh_op_bnr_1')
// (8, 2, 'local_g0_1')
// (8, 2, 'lutff_1/in_0')
// (8, 2, 'neigh_op_top_1')
// (8, 3, 'lutff_1/out')
// (8, 4, 'neigh_op_bot_1')
// (9, 2, 'neigh_op_tnl_1')
// (9, 3, 'neigh_op_lft_1')
// (9, 4, 'neigh_op_bnl_1')

wire n950;
// (7, 2, 'neigh_op_tnr_2')
// (7, 3, 'neigh_op_rgt_2')
// (7, 4, 'local_g0_2')
// (7, 4, 'lutff_5/in_3')
// (7, 4, 'neigh_op_bnr_2')
// (8, 2, 'neigh_op_top_2')
// (8, 3, 'lutff_2/out')
// (8, 4, 'neigh_op_bot_2')
// (9, 2, 'neigh_op_tnl_2')
// (9, 3, 'neigh_op_lft_2')
// (9, 4, 'neigh_op_bnl_2')

reg n951 = 0;
// (7, 2, 'neigh_op_tnr_3')
// (7, 3, 'neigh_op_rgt_3')
// (7, 4, 'neigh_op_bnr_3')
// (8, 1, 'sp4_r_v_b_31')
// (8, 2, 'local_g1_3')
// (8, 2, 'lutff_7/in_3')
// (8, 2, 'neigh_op_top_3')
// (8, 2, 'sp4_r_v_b_18')
// (8, 3, 'lutff_3/out')
// (8, 3, 'sp4_r_v_b_7')
// (8, 4, 'neigh_op_bot_3')
// (9, 0, 'span4_vert_31')
// (9, 1, 'local_g3_7')
// (9, 1, 'lutff_4/in_0')
// (9, 1, 'sp4_v_b_31')
// (9, 2, 'neigh_op_tnl_3')
// (9, 2, 'sp4_v_b_18')
// (9, 3, 'neigh_op_lft_3')
// (9, 3, 'sp4_v_b_7')
// (9, 4, 'neigh_op_bnl_3')

wire n952;
// (7, 2, 'neigh_op_tnr_4')
// (7, 3, 'neigh_op_rgt_4')
// (7, 4, 'local_g0_4')
// (7, 4, 'lutff_2/in_2')
// (7, 4, 'neigh_op_bnr_4')
// (8, 2, 'neigh_op_top_4')
// (8, 3, 'lutff_4/out')
// (8, 4, 'neigh_op_bot_4')
// (9, 2, 'neigh_op_tnl_4')
// (9, 3, 'neigh_op_lft_4')
// (9, 4, 'neigh_op_bnl_4')

reg n953 = 0;
// (7, 2, 'neigh_op_tnr_5')
// (7, 3, 'neigh_op_rgt_5')
// (7, 4, 'neigh_op_bnr_5')
// (8, 2, 'local_g0_5')
// (8, 2, 'lutff_5/in_2')
// (8, 2, 'neigh_op_top_5')
// (8, 3, 'local_g1_5')
// (8, 3, 'lutff_5/out')
// (8, 3, 'lutff_7/in_1')
// (8, 4, 'neigh_op_bot_5')
// (9, 2, 'neigh_op_tnl_5')
// (9, 3, 'neigh_op_lft_5')
// (9, 4, 'neigh_op_bnl_5')

reg n954 = 0;
// (7, 2, 'neigh_op_tnr_6')
// (7, 3, 'local_g3_6')
// (7, 3, 'lutff_1/in_0')
// (7, 3, 'neigh_op_rgt_6')
// (7, 4, 'neigh_op_bnr_6')
// (8, 1, 'sp4_r_v_b_37')
// (8, 2, 'neigh_op_top_6')
// (8, 2, 'sp4_r_v_b_24')
// (8, 3, 'lutff_6/out')
// (8, 3, 'sp4_r_v_b_13')
// (8, 4, 'neigh_op_bot_6')
// (8, 4, 'sp4_r_v_b_0')
// (9, 0, 'span4_vert_37')
// (9, 1, 'local_g2_5')
// (9, 1, 'lutff_4/in_1')
// (9, 1, 'sp4_v_b_37')
// (9, 2, 'neigh_op_tnl_6')
// (9, 2, 'sp4_v_b_24')
// (9, 3, 'neigh_op_lft_6')
// (9, 3, 'sp4_v_b_13')
// (9, 4, 'neigh_op_bnl_6')
// (9, 4, 'sp4_v_b_0')

wire n955;
// (7, 2, 'neigh_op_tnr_7')
// (7, 3, 'neigh_op_rgt_7')
// (7, 4, 'local_g0_7')
// (7, 4, 'lutff_5/in_2')
// (7, 4, 'neigh_op_bnr_7')
// (8, 2, 'neigh_op_top_7')
// (8, 3, 'lutff_7/out')
// (8, 4, 'neigh_op_bot_7')
// (9, 2, 'neigh_op_tnl_7')
// (9, 3, 'neigh_op_lft_7')
// (9, 4, 'neigh_op_bnl_7')

wire n956;
// (7, 2, 'sp4_h_r_3')
// (7, 4, 'sp4_r_v_b_44')
// (7, 5, 'sp4_r_v_b_33')
// (7, 6, 'sp4_r_v_b_20')
// (7, 7, 'sp4_r_v_b_9')
// (8, 2, 'sp4_h_r_14')
// (8, 3, 'sp4_h_r_3')
// (8, 3, 'sp4_v_t_44')
// (8, 4, 'sp4_v_b_44')
// (8, 5, 'local_g3_1')
// (8, 5, 'lutff_4/in_0')
// (8, 5, 'sp4_v_b_33')
// (8, 6, 'local_g0_4')
// (8, 6, 'lutff_1/in_1')
// (8, 6, 'sp4_v_b_20')
// (8, 7, 'sp4_v_b_9')
// (9, 2, 'local_g2_3')
// (9, 2, 'lutff_4/in_3')
// (9, 2, 'sp4_h_r_27')
// (9, 3, 'sp4_h_r_14')
// (10, 2, 'local_g2_3')
// (10, 2, 'lutff_3/in_0')
// (10, 2, 'lutff_4/in_1')
// (10, 2, 'neigh_op_tnr_3')
// (10, 2, 'sp4_h_r_38')
// (10, 3, 'local_g3_3')
// (10, 3, 'lutff_6/in_0')
// (10, 3, 'neigh_op_rgt_3')
// (10, 3, 'sp4_h_r_11')
// (10, 3, 'sp4_h_r_27')
// (10, 3, 'sp4_r_v_b_38')
// (10, 4, 'local_g0_3')
// (10, 4, 'local_g1_3')
// (10, 4, 'lutff_1/in_1')
// (10, 4, 'lutff_2/in_1')
// (10, 4, 'lutff_3/in_3')
// (10, 4, 'neigh_op_bnr_3')
// (10, 4, 'sp4_r_v_b_27')
// (10, 5, 'local_g2_6')
// (10, 5, 'lutff_7/in_1')
// (10, 5, 'sp4_r_v_b_14')
// (10, 6, 'sp4_r_v_b_3')
// (11, 1, 'sp4_r_v_b_47')
// (11, 2, 'local_g1_3')
// (11, 2, 'lutff_2/in_0')
// (11, 2, 'neigh_op_top_3')
// (11, 2, 'sp4_h_l_38')
// (11, 2, 'sp4_r_v_b_34')
// (11, 2, 'sp4_v_t_38')
// (11, 3, 'lutff_3/out')
// (11, 3, 'sp4_h_r_22')
// (11, 3, 'sp4_h_r_38')
// (11, 3, 'sp4_r_v_b_23')
// (11, 3, 'sp4_r_v_b_39')
// (11, 3, 'sp4_v_b_38')
// (11, 4, 'neigh_op_bot_3')
// (11, 4, 'sp4_r_v_b_10')
// (11, 4, 'sp4_r_v_b_26')
// (11, 4, 'sp4_v_b_27')
// (11, 5, 'sp4_r_v_b_15')
// (11, 5, 'sp4_r_v_b_36')
// (11, 5, 'sp4_v_b_14')
// (11, 6, 'sp4_r_v_b_2')
// (11, 6, 'sp4_r_v_b_25')
// (11, 6, 'sp4_v_b_3')
// (11, 7, 'sp4_r_v_b_12')
// (11, 8, 'sp4_r_v_b_1')
// (12, 0, 'span4_vert_47')
// (12, 1, 'sp4_v_b_47')
// (12, 2, 'neigh_op_tnl_3')
// (12, 2, 'sp4_v_b_34')
// (12, 2, 'sp4_v_t_39')
// (12, 3, 'neigh_op_lft_3')
// (12, 3, 'sp4_h_l_38')
// (12, 3, 'sp4_h_r_35')
// (12, 3, 'sp4_v_b_23')
// (12, 3, 'sp4_v_b_39')
// (12, 4, 'local_g3_3')
// (12, 4, 'lutff_5/in_3')
// (12, 4, 'neigh_op_bnl_3')
// (12, 4, 'sp4_v_b_10')
// (12, 4, 'sp4_v_b_26')
// (12, 4, 'sp4_v_t_36')
// (12, 5, 'local_g1_7')
// (12, 5, 'lutff_6/in_2')
// (12, 5, 'sp4_v_b_15')
// (12, 5, 'sp4_v_b_36')
// (12, 6, 'local_g1_2')
// (12, 6, 'lutff_1/in_0')
// (12, 6, 'lutff_3/in_0')
// (12, 6, 'lutff_7/in_0')
// (12, 6, 'sp4_v_b_2')
// (12, 6, 'sp4_v_b_25')
// (12, 7, 'local_g0_4')
// (12, 7, 'lutff_7/in_1')
// (12, 7, 'sp4_v_b_12')
// (12, 8, 'sp4_v_b_1')
// (13, 3, 'sp4_h_r_46')
// (13, 4, 'sp4_r_v_b_46')
// (13, 5, 'local_g2_3')
// (13, 5, 'lutff_0/in_3')
// (13, 5, 'sp4_r_v_b_35')
// (13, 6, 'sp4_r_v_b_22')
// (13, 7, 'sp4_r_v_b_11')
// (14, 3, 'sp4_h_l_46')
// (14, 3, 'sp4_v_t_46')
// (14, 4, 'local_g2_6')
// (14, 4, 'lutff_2/in_0')
// (14, 4, 'sp4_v_b_46')
// (14, 5, 'local_g2_3')
// (14, 5, 'lutff_1/in_0')
// (14, 5, 'sp4_v_b_35')
// (14, 6, 'sp4_v_b_22')
// (14, 7, 'local_g0_3')
// (14, 7, 'lutff_5/in_0')
// (14, 7, 'sp4_v_b_11')

wire n957;
// (7, 2, 'sp4_r_v_b_38')
// (7, 3, 'neigh_op_tnr_7')
// (7, 3, 'sp4_r_v_b_27')
// (7, 4, 'neigh_op_rgt_7')
// (7, 4, 'sp4_r_v_b_14')
// (7, 5, 'neigh_op_bnr_7')
// (7, 5, 'sp4_r_v_b_3')
// (8, 1, 'sp4_v_t_38')
// (8, 2, 'local_g3_6')
// (8, 2, 'lutff_1/in_2')
// (8, 2, 'sp4_v_b_38')
// (8, 3, 'neigh_op_top_7')
// (8, 3, 'sp4_v_b_27')
// (8, 4, 'lutff_7/out')
// (8, 4, 'sp4_v_b_14')
// (8, 5, 'neigh_op_bot_7')
// (8, 5, 'sp4_v_b_3')
// (9, 3, 'neigh_op_tnl_7')
// (9, 4, 'neigh_op_lft_7')
// (9, 5, 'neigh_op_bnl_7')

wire n958;
// (7, 2, 'sp4_r_v_b_41')
// (7, 3, 'local_g0_4')
// (7, 3, 'lutff_3/in_3')
// (7, 3, 'sp4_r_v_b_28')
// (7, 4, 'local_g2_2')
// (7, 4, 'lutff_0/in_0')
// (7, 4, 'neigh_op_tnr_2')
// (7, 4, 'sp4_r_v_b_17')
// (7, 5, 'local_g2_2')
// (7, 5, 'lutff_7/in_3')
// (7, 5, 'neigh_op_rgt_2')
// (7, 5, 'sp4_r_v_b_4')
// (7, 6, 'neigh_op_bnr_2')
// (8, 1, 'sp4_v_t_41')
// (8, 2, 'sp4_v_b_41')
// (8, 3, 'sp4_v_b_28')
// (8, 4, 'local_g0_1')
// (8, 4, 'lutff_3/in_2')
// (8, 4, 'neigh_op_top_2')
// (8, 4, 'sp4_v_b_17')
// (8, 5, 'local_g1_2')
// (8, 5, 'lutff_2/out')
// (8, 5, 'lutff_3/in_2')
// (8, 5, 'lutff_5/in_2')
// (8, 5, 'sp4_v_b_4')
// (8, 6, 'neigh_op_bot_2')
// (9, 4, 'neigh_op_tnl_2')
// (9, 5, 'neigh_op_lft_2')
// (9, 6, 'neigh_op_bnl_2')

wire n959;
// (7, 3, 'local_g1_3')
// (7, 3, 'lutff_1/in_3')
// (7, 3, 'sp4_h_r_3')
// (8, 3, 'sp4_h_r_14')
// (9, 2, 'neigh_op_tnr_3')
// (9, 3, 'neigh_op_rgt_3')
// (9, 3, 'sp4_h_r_27')
// (9, 4, 'neigh_op_bnr_3')
// (10, 2, 'neigh_op_top_3')
// (10, 3, 'lutff_3/out')
// (10, 3, 'sp4_h_r_38')
// (10, 4, 'neigh_op_bot_3')
// (11, 2, 'neigh_op_tnl_3')
// (11, 3, 'neigh_op_lft_3')
// (11, 3, 'sp4_h_l_38')
// (11, 4, 'neigh_op_bnl_3')

wire n960;
// (7, 3, 'local_g3_7')
// (7, 3, 'lutff_3/in_1')
// (7, 3, 'sp4_r_v_b_47')
// (7, 4, 'sp4_r_v_b_34')
// (7, 5, 'local_g3_7')
// (7, 5, 'lutff_7/in_1')
// (7, 5, 'sp4_r_v_b_23')
// (7, 6, 'sp4_r_v_b_10')
// (8, 2, 'sp4_v_t_47')
// (8, 3, 'sp4_v_b_47')
// (8, 4, 'sp4_v_b_34')
// (8, 5, 'sp4_v_b_23')
// (8, 6, 'local_g0_2')
// (8, 6, 'lutff_0/in_0')
// (8, 6, 'sp4_h_r_10')
// (8, 6, 'sp4_v_b_10')
// (9, 3, 'sp4_r_v_b_39')
// (9, 4, 'sp4_r_v_b_26')
// (9, 5, 'neigh_op_tnr_1')
// (9, 5, 'sp4_r_v_b_15')
// (9, 6, 'neigh_op_rgt_1')
// (9, 6, 'sp4_h_r_23')
// (9, 6, 'sp4_r_v_b_2')
// (9, 7, 'neigh_op_bnr_1')
// (10, 2, 'sp4_h_r_7')
// (10, 2, 'sp4_v_t_39')
// (10, 3, 'sp4_v_b_39')
// (10, 4, 'sp4_v_b_26')
// (10, 5, 'neigh_op_top_1')
// (10, 5, 'sp4_v_b_15')
// (10, 6, 'lutff_1/out')
// (10, 6, 'sp4_h_r_34')
// (10, 6, 'sp4_v_b_2')
// (10, 7, 'neigh_op_bot_1')
// (11, 2, 'local_g0_2')
// (11, 2, 'lutff_0/in_2')
// (11, 2, 'sp4_h_r_18')
// (11, 5, 'neigh_op_tnl_1')
// (11, 6, 'neigh_op_lft_1')
// (11, 6, 'sp4_h_r_47')
// (11, 7, 'neigh_op_bnl_1')
// (12, 2, 'sp4_h_r_31')
// (12, 6, 'sp4_h_l_47')
// (13, 2, 'sp4_h_r_42')
// (14, 2, 'sp4_h_l_42')

reg n961 = 0;
// (7, 3, 'neigh_op_tnr_0')
// (7, 4, 'neigh_op_rgt_0')
// (7, 5, 'neigh_op_bnr_0')
// (8, 3, 'neigh_op_top_0')
// (8, 3, 'sp4_r_v_b_44')
// (8, 4, 'local_g2_0')
// (8, 4, 'lutff_0/out')
// (8, 4, 'lutff_6/in_2')
// (8, 4, 'sp4_r_v_b_33')
// (8, 5, 'neigh_op_bot_0')
// (8, 5, 'sp4_r_v_b_20')
// (8, 6, 'sp4_r_v_b_9')
// (9, 2, 'local_g1_1')
// (9, 2, 'lutff_3/in_3')
// (9, 2, 'sp4_h_r_9')
// (9, 2, 'sp4_v_t_44')
// (9, 3, 'neigh_op_tnl_0')
// (9, 3, 'sp4_v_b_44')
// (9, 4, 'neigh_op_lft_0')
// (9, 4, 'sp4_v_b_33')
// (9, 5, 'neigh_op_bnl_0')
// (9, 5, 'sp4_v_b_20')
// (9, 6, 'sp4_v_b_9')
// (10, 2, 'sp4_h_r_20')
// (11, 2, 'sp4_h_r_33')
// (12, 2, 'sp4_h_r_44')
// (13, 2, 'sp4_h_l_44')

wire n962;
// (7, 3, 'neigh_op_tnr_1')
// (7, 4, 'local_g3_1')
// (7, 4, 'lutff_7/in_3')
// (7, 4, 'neigh_op_rgt_1')
// (7, 5, 'neigh_op_bnr_1')
// (8, 3, 'neigh_op_top_1')
// (8, 4, 'lutff_1/out')
// (8, 5, 'neigh_op_bot_1')
// (9, 3, 'neigh_op_tnl_1')
// (9, 4, 'neigh_op_lft_1')
// (9, 5, 'neigh_op_bnl_1')

wire n963;
// (7, 3, 'neigh_op_tnr_2')
// (7, 4, 'neigh_op_rgt_2')
// (7, 5, 'local_g1_2')
// (7, 5, 'lutff_5/in_0')
// (7, 5, 'neigh_op_bnr_2')
// (8, 3, 'neigh_op_top_2')
// (8, 4, 'lutff_2/out')
// (8, 5, 'neigh_op_bot_2')
// (9, 3, 'neigh_op_tnl_2')
// (9, 4, 'neigh_op_lft_2')
// (9, 5, 'neigh_op_bnl_2')

reg n964 = 0;
// (7, 3, 'neigh_op_tnr_4')
// (7, 4, 'neigh_op_rgt_4')
// (7, 5, 'neigh_op_bnr_4')
// (8, 1, 'sp4_r_v_b_44')
// (8, 2, 'sp4_r_v_b_33')
// (8, 3, 'neigh_op_top_4')
// (8, 3, 'sp4_r_v_b_20')
// (8, 4, 'local_g2_4')
// (8, 4, 'lutff_2/in_0')
// (8, 4, 'lutff_4/out')
// (8, 4, 'sp4_r_v_b_9')
// (8, 5, 'neigh_op_bot_4')
// (9, 0, 'span4_vert_44')
// (9, 1, 'sp4_v_b_44')
// (9, 2, 'local_g2_1')
// (9, 2, 'lutff_3/in_0')
// (9, 2, 'sp4_v_b_33')
// (9, 3, 'neigh_op_tnl_4')
// (9, 3, 'sp4_v_b_20')
// (9, 4, 'neigh_op_lft_4')
// (9, 4, 'sp4_v_b_9')
// (9, 5, 'neigh_op_bnl_4')

wire n965;
// (7, 3, 'neigh_op_tnr_6')
// (7, 4, 'local_g3_6')
// (7, 4, 'lutff_3/in_0')
// (7, 4, 'neigh_op_rgt_6')
// (7, 5, 'neigh_op_bnr_6')
// (8, 3, 'neigh_op_top_6')
// (8, 4, 'lutff_6/out')
// (8, 5, 'neigh_op_bot_6')
// (9, 3, 'neigh_op_tnl_6')
// (9, 4, 'neigh_op_lft_6')
// (9, 5, 'neigh_op_bnl_6')

reg n966 = 0;
// (7, 3, 'sp4_h_r_0')
// (8, 2, 'neigh_op_tnr_4')
// (8, 3, 'neigh_op_rgt_4')
// (8, 3, 'sp4_h_r_13')
// (8, 4, 'local_g0_4')
// (8, 4, 'lutff_5/in_1')
// (8, 4, 'neigh_op_bnr_4')
// (9, 2, 'neigh_op_top_4')
// (9, 3, 'lutff_4/out')
// (9, 3, 'sp4_h_r_24')
// (9, 4, 'neigh_op_bot_4')
// (10, 1, 'sp4_r_v_b_30')
// (10, 2, 'neigh_op_tnl_4')
// (10, 2, 'sp4_r_v_b_19')
// (10, 3, 'neigh_op_lft_4')
// (10, 3, 'sp4_h_r_37')
// (10, 3, 'sp4_r_v_b_6')
// (10, 4, 'neigh_op_bnl_4')
// (11, 0, 'span4_vert_30')
// (11, 1, 'sp4_v_b_30')
// (11, 2, 'local_g0_3')
// (11, 2, 'lutff_3/in_2')
// (11, 2, 'sp4_v_b_19')
// (11, 3, 'sp4_h_l_37')
// (11, 3, 'sp4_v_b_6')

wire n967;
// (7, 3, 'sp4_r_v_b_42')
// (7, 4, 'local_g1_3')
// (7, 4, 'lutff_0/in_2')
// (7, 4, 'sp4_h_r_11')
// (7, 4, 'sp4_r_v_b_31')
// (7, 5, 'sp4_r_v_b_18')
// (7, 6, 'local_g1_7')
// (7, 6, 'lutff_0/in_2')
// (7, 6, 'lutff_5/in_1')
// (7, 6, 'sp4_r_v_b_7')
// (8, 2, 'sp4_v_t_42')
// (8, 3, 'sp4_v_b_42')
// (8, 4, 'sp4_h_r_22')
// (8, 4, 'sp4_v_b_31')
// (8, 5, 'sp4_v_b_18')
// (8, 6, 'sp4_h_r_2')
// (8, 6, 'sp4_v_b_7')
// (9, 4, 'sp4_h_r_35')
// (9, 6, 'local_g1_7')
// (9, 6, 'lutff_5/in_3')
// (9, 6, 'sp4_h_r_15')
// (10, 4, 'sp4_h_r_46')
// (10, 6, 'sp4_h_r_26')
// (11, 4, 'sp4_h_l_46')
// (11, 4, 'sp4_h_r_11')
// (11, 6, 'sp4_h_r_39')
// (12, 4, 'sp4_h_r_22')
// (12, 6, 'sp4_h_l_39')
// (12, 6, 'sp4_h_r_2')
// (13, 4, 'sp4_h_r_35')
// (13, 6, 'sp4_h_r_15')
// (14, 1, 'sp4_r_v_b_46')
// (14, 2, 'local_g3_3')
// (14, 2, 'lutff_0/in_2')
// (14, 2, 'neigh_op_tnr_3')
// (14, 2, 'sp4_r_v_b_35')
// (14, 3, 'neigh_op_rgt_3')
// (14, 3, 'sp4_r_v_b_22')
// (14, 4, 'neigh_op_bnr_3')
// (14, 4, 'sp4_h_r_46')
// (14, 4, 'sp4_r_v_b_11')
// (14, 6, 'sp4_h_r_26')
// (15, 0, 'span4_vert_46')
// (15, 1, 'sp4_v_b_46')
// (15, 2, 'neigh_op_top_3')
// (15, 2, 'sp4_v_b_35')
// (15, 3, 'lutff_3/out')
// (15, 3, 'sp4_r_v_b_39')
// (15, 3, 'sp4_v_b_22')
// (15, 4, 'neigh_op_bot_3')
// (15, 4, 'sp4_h_l_46')
// (15, 4, 'sp4_r_v_b_26')
// (15, 4, 'sp4_v_b_11')
// (15, 5, 'sp4_r_v_b_15')
// (15, 6, 'sp4_h_r_39')
// (15, 6, 'sp4_r_v_b_2')
// (16, 2, 'neigh_op_tnl_3')
// (16, 2, 'sp4_v_t_39')
// (16, 3, 'neigh_op_lft_3')
// (16, 3, 'sp4_v_b_39')
// (16, 4, 'neigh_op_bnl_3')
// (16, 4, 'sp4_v_b_26')
// (16, 5, 'sp4_v_b_15')
// (16, 6, 'sp4_h_l_39')
// (16, 6, 'sp4_v_b_2')

reg n968 = 0;
// (7, 4, 'neigh_op_tnr_0')
// (7, 5, 'neigh_op_rgt_0')
// (7, 6, 'neigh_op_bnr_0')
// (8, 2, 'sp4_r_v_b_36')
// (8, 3, 'sp4_r_v_b_25')
// (8, 4, 'neigh_op_top_0')
// (8, 4, 'sp4_r_v_b_12')
// (8, 5, 'lutff_0/out')
// (8, 5, 'sp4_r_v_b_1')
// (8, 6, 'neigh_op_bot_0')
// (9, 1, 'sp4_v_t_36')
// (9, 2, 'local_g2_4')
// (9, 2, 'lutff_6/in_2')
// (9, 2, 'sp4_v_b_36')
// (9, 3, 'sp4_v_b_25')
// (9, 4, 'neigh_op_tnl_0')
// (9, 4, 'sp4_v_b_12')
// (9, 5, 'local_g1_0')
// (9, 5, 'lutff_4/in_1')
// (9, 5, 'neigh_op_lft_0')
// (9, 5, 'sp4_v_b_1')
// (9, 6, 'neigh_op_bnl_0')

reg n969 = 0;
// (7, 4, 'neigh_op_tnr_1')
// (7, 5, 'neigh_op_rgt_1')
// (7, 6, 'neigh_op_bnr_1')
// (8, 2, 'sp4_r_v_b_38')
// (8, 3, 'sp4_r_v_b_27')
// (8, 4, 'neigh_op_top_1')
// (8, 4, 'sp4_r_v_b_14')
// (8, 5, 'local_g1_1')
// (8, 5, 'lutff_1/out')
// (8, 5, 'lutff_6/in_0')
// (8, 5, 'sp4_r_v_b_3')
// (8, 6, 'neigh_op_bot_1')
// (9, 1, 'sp4_v_t_38')
// (9, 2, 'local_g3_6')
// (9, 2, 'lutff_6/in_1')
// (9, 2, 'sp4_v_b_38')
// (9, 3, 'sp4_v_b_27')
// (9, 4, 'neigh_op_tnl_1')
// (9, 4, 'sp4_v_b_14')
// (9, 5, 'neigh_op_lft_1')
// (9, 5, 'sp4_v_b_3')
// (9, 6, 'neigh_op_bnl_1')

wire n970;
// (7, 4, 'neigh_op_tnr_4')
// (7, 5, 'neigh_op_rgt_4')
// (7, 6, 'local_g0_4')
// (7, 6, 'lutff_2/in_0')
// (7, 6, 'neigh_op_bnr_4')
// (8, 4, 'neigh_op_top_4')
// (8, 5, 'lutff_4/out')
// (8, 6, 'neigh_op_bot_4')
// (9, 4, 'neigh_op_tnl_4')
// (9, 5, 'neigh_op_lft_4')
// (9, 6, 'neigh_op_bnl_4')

wire n971;
// (7, 4, 'neigh_op_tnr_7')
// (7, 5, 'neigh_op_rgt_7')
// (7, 6, 'neigh_op_bnr_7')
// (8, 4, 'local_g0_7')
// (8, 4, 'lutff_2/in_3')
// (8, 4, 'lutff_6/in_3')
// (8, 4, 'neigh_op_top_7')
// (8, 5, 'local_g0_7')
// (8, 5, 'lutff_6/in_3')
// (8, 5, 'lutff_7/out')
// (8, 6, 'neigh_op_bot_7')
// (9, 4, 'neigh_op_tnl_7')
// (9, 5, 'neigh_op_lft_7')
// (9, 6, 'neigh_op_bnl_7')

wire n972;
// (7, 4, 'sp4_h_r_2')
// (8, 4, 'local_g1_7')
// (8, 4, 'lutff_5/in_3')
// (8, 4, 'sp4_h_r_15')
// (9, 2, 'neigh_op_tnr_7')
// (9, 3, 'neigh_op_rgt_7')
// (9, 4, 'neigh_op_bnr_7')
// (9, 4, 'sp4_h_r_26')
// (10, 1, 'sp4_r_v_b_39')
// (10, 2, 'neigh_op_top_7')
// (10, 2, 'sp4_r_v_b_26')
// (10, 3, 'lutff_7/out')
// (10, 3, 'sp4_r_v_b_15')
// (10, 4, 'neigh_op_bot_7')
// (10, 4, 'sp4_h_r_39')
// (10, 4, 'sp4_r_v_b_2')
// (11, 0, 'span4_vert_39')
// (11, 1, 'sp4_v_b_39')
// (11, 2, 'neigh_op_tnl_7')
// (11, 2, 'sp4_v_b_26')
// (11, 3, 'neigh_op_lft_7')
// (11, 3, 'sp4_v_b_15')
// (11, 4, 'neigh_op_bnl_7')
// (11, 4, 'sp4_h_l_39')
// (11, 4, 'sp4_v_b_2')

wire n973;
// (7, 4, 'sp4_h_r_3')
// (8, 4, 'local_g0_6')
// (8, 4, 'lutff_3/in_1')
// (8, 4, 'sp4_h_r_14')
// (8, 5, 'sp4_r_v_b_46')
// (8, 6, 'local_g0_0')
// (8, 6, 'lutff_3/in_1')
// (8, 6, 'lutff_4/in_0')
// (8, 6, 'sp4_r_v_b_35')
// (8, 7, 'sp4_r_v_b_22')
// (8, 8, 'sp4_r_v_b_11')
// (9, 4, 'sp4_h_r_11')
// (9, 4, 'sp4_h_r_27')
// (9, 4, 'sp4_v_t_46')
// (9, 5, 'sp4_v_b_46')
// (9, 6, 'local_g2_3')
// (9, 6, 'lutff_7/in_0')
// (9, 6, 'sp4_v_b_35')
// (9, 7, 'local_g0_6')
// (9, 7, 'local_g1_6')
// (9, 7, 'lutff_1/in_1')
// (9, 7, 'lutff_2/in_3')
// (9, 7, 'sp4_v_b_22')
// (9, 8, 'sp4_v_b_11')
// (10, 4, 'sp4_h_r_22')
// (10, 4, 'sp4_h_r_38')
// (11, 3, 'neigh_op_tnr_7')
// (11, 4, 'neigh_op_rgt_7')
// (11, 4, 'sp4_h_l_38')
// (11, 4, 'sp4_h_r_3')
// (11, 4, 'sp4_h_r_35')
// (11, 5, 'neigh_op_bnr_7')
// (12, 3, 'neigh_op_top_7')
// (12, 4, 'local_g2_7')
// (12, 4, 'lutff_1/in_2')
// (12, 4, 'lutff_7/out')
// (12, 4, 'sp4_h_r_14')
// (12, 4, 'sp4_h_r_46')
// (12, 5, 'neigh_op_bot_7')
// (13, 3, 'neigh_op_tnl_7')
// (13, 4, 'neigh_op_lft_7')
// (13, 4, 'sp4_h_l_46')
// (13, 4, 'sp4_h_r_27')
// (13, 5, 'neigh_op_bnl_7')
// (14, 4, 'sp4_h_r_38')
// (15, 4, 'sp4_h_l_38')

wire n974;
// (7, 4, 'sp4_h_r_7')
// (8, 4, 'local_g0_2')
// (8, 4, 'lutff_1/in_3')
// (8, 4, 'sp4_h_r_18')
// (9, 3, 'neigh_op_tnr_5')
// (9, 4, 'neigh_op_rgt_5')
// (9, 4, 'sp4_h_r_31')
// (9, 5, 'neigh_op_bnr_5')
// (10, 3, 'neigh_op_top_5')
// (10, 4, 'lutff_5/out')
// (10, 4, 'sp4_h_r_42')
// (10, 5, 'neigh_op_bot_5')
// (11, 3, 'neigh_op_tnl_5')
// (11, 4, 'neigh_op_lft_5')
// (11, 4, 'sp4_h_l_42')
// (11, 5, 'neigh_op_bnl_5')

wire n975;
// (7, 5, 'local_g0_5')
// (7, 5, 'lutff_7/in_0')
// (7, 5, 'sp4_h_r_5')
// (8, 5, 'sp4_h_r_16')
// (9, 5, 'sp4_h_r_29')
// (10, 4, 'neigh_op_tnr_1')
// (10, 5, 'local_g2_1')
// (10, 5, 'lutff_1/in_0')
// (10, 5, 'neigh_op_rgt_1')
// (10, 5, 'sp4_h_r_40')
// (10, 6, 'local_g1_1')
// (10, 6, 'lutff_3/in_1')
// (10, 6, 'neigh_op_bnr_1')
// (11, 4, 'local_g1_1')
// (11, 4, 'lutff_2/in_2')
// (11, 4, 'neigh_op_top_1')
// (11, 5, 'lutff_1/out')
// (11, 5, 'sp4_h_l_40')
// (11, 5, 'sp4_h_r_2')
// (11, 6, 'neigh_op_bot_1')
// (12, 4, 'neigh_op_tnl_1')
// (12, 5, 'neigh_op_lft_1')
// (12, 5, 'sp4_h_r_15')
// (12, 6, 'neigh_op_bnl_1')
// (13, 5, 'sp4_h_r_26')
// (14, 5, 'sp4_h_r_39')
// (15, 5, 'sp4_h_l_39')

wire n976;
// (7, 5, 'local_g3_2')
// (7, 5, 'lutff_7/in_2')
// (7, 5, 'neigh_op_tnr_2')
// (7, 6, 'local_g3_2')
// (7, 6, 'lutff_0/in_1')
// (7, 6, 'neigh_op_rgt_2')
// (7, 7, 'neigh_op_bnr_2')
// (8, 5, 'local_g0_2')
// (8, 5, 'lutff_3/in_3')
// (8, 5, 'lutff_5/in_3')
// (8, 5, 'neigh_op_top_2')
// (8, 6, 'lutff_2/out')
// (8, 7, 'neigh_op_bot_2')
// (9, 5, 'neigh_op_tnl_2')
// (9, 6, 'neigh_op_lft_2')
// (9, 7, 'neigh_op_bnl_2')

wire n977;
// (7, 5, 'neigh_op_tnr_1')
// (7, 6, 'local_g3_1')
// (7, 6, 'lutff_0/in_0')
// (7, 6, 'neigh_op_rgt_1')
// (7, 7, 'neigh_op_bnr_1')
// (8, 5, 'neigh_op_top_1')
// (8, 6, 'lutff_1/out')
// (8, 7, 'neigh_op_bot_1')
// (9, 5, 'neigh_op_tnl_1')
// (9, 6, 'neigh_op_lft_1')
// (9, 7, 'neigh_op_bnl_1')

wire n978;
// (7, 5, 'neigh_op_tnr_3')
// (7, 6, 'neigh_op_rgt_3')
// (7, 7, 'neigh_op_bnr_3')
// (8, 5, 'neigh_op_top_3')
// (8, 6, 'local_g1_3')
// (8, 6, 'lutff_3/out')
// (8, 6, 'lutff_7/in_3')
// (8, 7, 'neigh_op_bot_3')
// (9, 5, 'neigh_op_tnl_3')
// (9, 6, 'neigh_op_lft_3')
// (9, 7, 'neigh_op_bnl_3')

wire n979;
// (7, 5, 'sp4_h_r_0')
// (8, 2, 'sp4_h_r_10')
// (8, 5, 'sp4_h_r_13')
// (9, 2, 'sp4_h_r_23')
// (9, 2, 'sp4_r_v_b_47')
// (9, 3, 'sp4_r_v_b_34')
// (9, 4, 'sp4_r_v_b_23')
// (9, 5, 'sp4_h_r_24')
// (9, 5, 'sp4_r_v_b_10')
// (10, 1, 'sp4_r_v_b_35')
// (10, 1, 'sp4_v_t_47')
// (10, 2, 'local_g2_2')
// (10, 2, 'lutff_global/cen')
// (10, 2, 'sp4_h_r_34')
// (10, 2, 'sp4_r_v_b_22')
// (10, 2, 'sp4_r_v_b_43')
// (10, 2, 'sp4_v_b_47')
// (10, 3, 'sp4_r_v_b_11')
// (10, 3, 'sp4_r_v_b_30')
// (10, 3, 'sp4_v_b_34')
// (10, 4, 'local_g3_3')
// (10, 4, 'lutff_global/cen')
// (10, 4, 'neigh_op_tnr_0')
// (10, 4, 'sp4_r_v_b_19')
// (10, 4, 'sp4_r_v_b_45')
// (10, 4, 'sp4_v_b_23')
// (10, 5, 'local_g0_2')
// (10, 5, 'lutff_global/cen')
// (10, 5, 'neigh_op_rgt_0')
// (10, 5, 'sp4_h_r_37')
// (10, 5, 'sp4_h_r_5')
// (10, 5, 'sp4_r_v_b_32')
// (10, 5, 'sp4_r_v_b_6')
// (10, 5, 'sp4_v_b_10')
// (10, 6, 'neigh_op_bnr_0')
// (10, 6, 'sp4_r_v_b_21')
// (10, 7, 'sp4_r_v_b_8')
// (11, 0, 'span12_vert_8')
// (11, 0, 'span4_vert_35')
// (11, 1, 'sp12_v_b_8')
// (11, 1, 'sp4_v_b_35')
// (11, 1, 'sp4_v_t_43')
// (11, 2, 'sp12_v_b_7')
// (11, 2, 'sp4_h_r_47')
// (11, 2, 'sp4_v_b_22')
// (11, 2, 'sp4_v_b_43')
// (11, 3, 'local_g1_3')
// (11, 3, 'lutff_global/cen')
// (11, 3, 'sp12_v_b_4')
// (11, 3, 'sp4_r_v_b_41')
// (11, 3, 'sp4_v_b_11')
// (11, 3, 'sp4_v_b_30')
// (11, 3, 'sp4_v_t_45')
// (11, 4, 'local_g3_3')
// (11, 4, 'lutff_global/cen')
// (11, 4, 'neigh_op_top_0')
// (11, 4, 'sp12_v_b_3')
// (11, 4, 'sp4_r_v_b_28')
// (11, 4, 'sp4_v_b_19')
// (11, 4, 'sp4_v_b_45')
// (11, 5, 'lutff_0/out')
// (11, 5, 'sp12_v_b_0')
// (11, 5, 'sp4_h_l_37')
// (11, 5, 'sp4_h_r_0')
// (11, 5, 'sp4_h_r_16')
// (11, 5, 'sp4_r_v_b_17')
// (11, 5, 'sp4_v_b_32')
// (11, 5, 'sp4_v_b_6')
// (11, 6, 'neigh_op_bot_0')
// (11, 6, 'sp4_r_v_b_4')
// (11, 6, 'sp4_v_b_21')
// (11, 7, 'sp4_v_b_8')
// (12, 2, 'sp4_h_l_47')
// (12, 2, 'sp4_v_t_41')
// (12, 3, 'sp4_v_b_41')
// (12, 4, 'neigh_op_tnl_0')
// (12, 4, 'sp4_v_b_28')
// (12, 5, 'neigh_op_lft_0')
// (12, 5, 'sp4_h_r_13')
// (12, 5, 'sp4_h_r_29')
// (12, 5, 'sp4_v_b_17')
// (12, 6, 'neigh_op_bnl_0')
// (12, 6, 'sp4_v_b_4')
// (13, 5, 'sp4_h_r_24')
// (13, 5, 'sp4_h_r_40')
// (14, 5, 'sp4_h_l_40')
// (14, 5, 'sp4_h_r_37')
// (15, 5, 'sp4_h_l_37')

wire n980;
// (7, 5, 'sp4_h_r_4')
// (8, 5, 'local_g0_1')
// (8, 5, 'lutff_5/in_0')
// (8, 5, 'sp4_h_r_17')
// (9, 5, 'sp4_h_r_28')
// (10, 2, 'sp4_r_v_b_36')
// (10, 3, 'sp4_r_v_b_25')
// (10, 4, 'sp4_r_v_b_12')
// (10, 5, 'sp4_h_r_41')
// (10, 5, 'sp4_r_v_b_1')
// (10, 6, 'local_g2_4')
// (10, 6, 'lutff_5/in_1')
// (10, 6, 'sp4_r_v_b_36')
// (10, 7, 'sp4_r_v_b_25')
// (10, 8, 'sp4_r_v_b_12')
// (10, 9, 'sp4_r_v_b_1')
// (11, 1, 'sp4_v_t_36')
// (11, 2, 'sp4_v_b_36')
// (11, 3, 'local_g3_1')
// (11, 3, 'lutff_0/in_0')
// (11, 3, 'sp4_v_b_25')
// (11, 4, 'sp4_v_b_12')
// (11, 5, 'sp4_h_l_41')
// (11, 5, 'sp4_h_r_1')
// (11, 5, 'sp4_v_b_1')
// (11, 5, 'sp4_v_t_36')
// (11, 6, 'sp4_v_b_36')
// (11, 7, 'sp4_v_b_25')
// (11, 8, 'sp4_v_b_12')
// (11, 9, 'sp4_v_b_1')
// (12, 5, 'sp4_h_r_12')
// (13, 4, 'local_g2_2')
// (13, 4, 'lutff_2/in_2')
// (13, 4, 'neigh_op_tnr_2')
// (13, 5, 'neigh_op_rgt_2')
// (13, 5, 'sp4_h_r_25')
// (13, 6, 'neigh_op_bnr_2')
// (14, 4, 'neigh_op_top_2')
// (14, 5, 'lutff_2/out')
// (14, 5, 'sp4_h_r_36')
// (14, 6, 'neigh_op_bot_2')
// (15, 4, 'neigh_op_tnl_2')
// (15, 5, 'neigh_op_lft_2')
// (15, 5, 'sp4_h_l_36')
// (15, 6, 'neigh_op_bnl_2')

wire n981;
// (7, 6, 'neigh_op_tnr_6')
// (7, 7, 'neigh_op_rgt_6')
// (7, 8, 'local_g0_6')
// (7, 8, 'local_g1_6')
// (7, 8, 'lutff_1/in_0')
// (7, 8, 'lutff_2/in_0')
// (7, 8, 'lutff_3/in_0')
// (7, 8, 'lutff_4/in_0')
// (7, 8, 'lutff_5/in_0')
// (7, 8, 'lutff_6/in_2')
// (7, 8, 'lutff_7/in_2')
// (7, 8, 'neigh_op_bnr_6')
// (8, 6, 'neigh_op_top_6')
// (8, 7, 'lutff_6/out')
// (8, 8, 'neigh_op_bot_6')
// (9, 6, 'neigh_op_tnl_6')
// (9, 7, 'neigh_op_lft_6')
// (9, 8, 'neigh_op_bnl_6')

wire n982;
// (7, 6, 'neigh_op_tnr_7')
// (7, 7, 'neigh_op_rgt_7')
// (7, 8, 'neigh_op_bnr_7')
// (8, 6, 'neigh_op_top_7')
// (8, 7, 'local_g2_7')
// (8, 7, 'lutff_0/in_1')
// (8, 7, 'lutff_7/out')
// (8, 8, 'neigh_op_bot_7')
// (9, 6, 'neigh_op_tnl_7')
// (9, 7, 'neigh_op_lft_7')
// (9, 8, 'neigh_op_bnl_7')

wire n983;
// (7, 6, 'sp4_h_r_1')
// (8, 6, 'local_g1_4')
// (8, 6, 'lutff_5/in_0')
// (8, 6, 'sp4_h_r_12')
// (9, 6, 'sp4_h_r_25')
// (10, 3, 'sp4_r_v_b_36')
// (10, 4, 'neigh_op_tnr_6')
// (10, 4, 'sp4_r_v_b_25')
// (10, 5, 'neigh_op_rgt_6')
// (10, 5, 'sp4_r_v_b_12')
// (10, 6, 'neigh_op_bnr_6')
// (10, 6, 'sp4_h_r_36')
// (10, 6, 'sp4_r_v_b_1')
// (11, 2, 'sp4_v_t_36')
// (11, 3, 'sp4_v_b_36')
// (11, 4, 'neigh_op_top_6')
// (11, 4, 'sp4_v_b_25')
// (11, 5, 'lutff_6/out')
// (11, 5, 'sp4_v_b_12')
// (11, 6, 'local_g1_6')
// (11, 6, 'lutff_0/in_1')
// (11, 6, 'neigh_op_bot_6')
// (11, 6, 'sp4_h_l_36')
// (11, 6, 'sp4_v_b_1')
// (12, 4, 'neigh_op_tnl_6')
// (12, 5, 'neigh_op_lft_6')
// (12, 6, 'neigh_op_bnl_6')

wire n984;
// (7, 6, 'sp4_h_r_7')
// (8, 6, 'sp4_h_r_18')
// (9, 3, 'sp4_r_v_b_47')
// (9, 4, 'sp4_r_v_b_34')
// (9, 5, 'neigh_op_tnr_5')
// (9, 5, 'sp4_r_v_b_23')
// (9, 5, 'sp4_r_v_b_39')
// (9, 6, 'neigh_op_rgt_5')
// (9, 6, 'sp4_h_r_31')
// (9, 6, 'sp4_r_v_b_10')
// (9, 6, 'sp4_r_v_b_26')
// (9, 7, 'neigh_op_bnr_5')
// (9, 7, 'sp4_r_v_b_15')
// (9, 7, 'sp4_r_v_b_43')
// (9, 8, 'sp4_r_v_b_2')
// (9, 8, 'sp4_r_v_b_30')
// (9, 9, 'sp4_r_v_b_19')
// (9, 9, 'sp4_r_v_b_39')
// (9, 9, 'sp4_r_v_b_40')
// (9, 10, 'local_g1_6')
// (9, 10, 'lutff_6/in_1')
// (9, 10, 'sp4_r_v_b_26')
// (9, 10, 'sp4_r_v_b_29')
// (9, 10, 'sp4_r_v_b_6')
// (9, 11, 'local_g3_0')
// (9, 11, 'lutff_7/in_0')
// (9, 11, 'sp4_r_v_b_15')
// (9, 11, 'sp4_r_v_b_16')
// (9, 11, 'sp4_r_v_b_39')
// (9, 11, 'sp4_r_v_b_43')
// (9, 12, 'sp4_r_v_b_2')
// (9, 12, 'sp4_r_v_b_26')
// (9, 12, 'sp4_r_v_b_30')
// (9, 12, 'sp4_r_v_b_5')
// (9, 13, 'local_g2_7')
// (9, 13, 'lutff_2/in_1')
// (9, 13, 'sp4_r_v_b_15')
// (9, 13, 'sp4_r_v_b_19')
// (9, 13, 'sp4_r_v_b_39')
// (9, 14, 'sp4_r_v_b_2')
// (9, 14, 'sp4_r_v_b_26')
// (9, 14, 'sp4_r_v_b_6')
// (9, 15, 'local_g2_7')
// (9, 15, 'lutff_3/in_2')
// (9, 15, 'lutff_5/in_0')
// (9, 15, 'sp4_r_v_b_15')
// (9, 16, 'sp4_r_v_b_2')
// (10, 0, 'span12_vert_21')
// (10, 1, 'sp12_v_b_21')
// (10, 2, 'sp12_v_b_18')
// (10, 2, 'sp4_v_t_47')
// (10, 3, 'sp12_v_b_17')
// (10, 3, 'sp4_v_b_47')
// (10, 4, 'sp12_v_b_14')
// (10, 4, 'sp4_v_b_34')
// (10, 4, 'sp4_v_t_39')
// (10, 5, 'neigh_op_top_5')
// (10, 5, 'sp12_v_b_13')
// (10, 5, 'sp4_v_b_23')
// (10, 5, 'sp4_v_b_39')
// (10, 6, 'lutff_5/out')
// (10, 6, 'sp12_v_b_10')
// (10, 6, 'sp4_h_r_42')
// (10, 6, 'sp4_r_v_b_43')
// (10, 6, 'sp4_v_b_10')
// (10, 6, 'sp4_v_b_26')
// (10, 6, 'sp4_v_t_43')
// (10, 7, 'local_g1_5')
// (10, 7, 'lutff_6/in_0')
// (10, 7, 'neigh_op_bot_5')
// (10, 7, 'sp12_v_b_9')
// (10, 7, 'sp4_r_v_b_30')
// (10, 7, 'sp4_r_v_b_37')
// (10, 7, 'sp4_v_b_15')
// (10, 7, 'sp4_v_b_43')
// (10, 8, 'local_g0_2')
// (10, 8, 'lutff_6/in_2')
// (10, 8, 'sp12_v_b_6')
// (10, 8, 'sp4_r_v_b_19')
// (10, 8, 'sp4_r_v_b_24')
// (10, 8, 'sp4_v_b_2')
// (10, 8, 'sp4_v_b_30')
// (10, 8, 'sp4_v_t_39')
// (10, 8, 'sp4_v_t_40')
// (10, 9, 'sp12_v_b_5')
// (10, 9, 'sp4_r_v_b_13')
// (10, 9, 'sp4_r_v_b_6')
// (10, 9, 'sp4_v_b_19')
// (10, 9, 'sp4_v_b_39')
// (10, 9, 'sp4_v_b_40')
// (10, 10, 'local_g2_2')
// (10, 10, 'lutff_0/in_0')
// (10, 10, 'sp12_v_b_2')
// (10, 10, 'sp4_r_v_b_0')
// (10, 10, 'sp4_r_v_b_39')
// (10, 10, 'sp4_v_b_26')
// (10, 10, 'sp4_v_b_29')
// (10, 10, 'sp4_v_b_6')
// (10, 10, 'sp4_v_t_39')
// (10, 10, 'sp4_v_t_43')
// (10, 11, 'local_g2_1')
// (10, 11, 'lutff_7/in_2')
// (10, 11, 'sp12_v_b_1')
// (10, 11, 'sp4_r_v_b_26')
// (10, 11, 'sp4_r_v_b_38')
// (10, 11, 'sp4_v_b_15')
// (10, 11, 'sp4_v_b_16')
// (10, 11, 'sp4_v_b_39')
// (10, 11, 'sp4_v_b_43')
// (10, 12, 'sp4_r_v_b_15')
// (10, 12, 'sp4_r_v_b_27')
// (10, 12, 'sp4_v_b_2')
// (10, 12, 'sp4_v_b_26')
// (10, 12, 'sp4_v_b_30')
// (10, 12, 'sp4_v_b_5')
// (10, 12, 'sp4_v_t_39')
// (10, 13, 'local_g1_2')
// (10, 13, 'lutff_5/in_2')
// (10, 13, 'lutff_7/in_0')
// (10, 13, 'sp4_r_v_b_14')
// (10, 13, 'sp4_r_v_b_2')
// (10, 13, 'sp4_v_b_15')
// (10, 13, 'sp4_v_b_19')
// (10, 13, 'sp4_v_b_39')
// (10, 14, 'local_g0_6')
// (10, 14, 'lutff_7/in_1')
// (10, 14, 'sp4_r_v_b_3')
// (10, 14, 'sp4_v_b_2')
// (10, 14, 'sp4_v_b_26')
// (10, 14, 'sp4_v_b_6')
// (10, 15, 'local_g0_7')
// (10, 15, 'lutff_1/in_0')
// (10, 15, 'lutff_2/in_3')
// (10, 15, 'lutff_5/in_0')
// (10, 15, 'sp4_v_b_15')
// (10, 16, 'sp4_v_b_2')
// (11, 5, 'neigh_op_tnl_5')
// (11, 5, 'sp4_v_t_43')
// (11, 6, 'neigh_op_lft_5')
// (11, 6, 'sp4_h_l_42')
// (11, 6, 'sp4_v_b_43')
// (11, 6, 'sp4_v_t_37')
// (11, 7, 'local_g2_5')
// (11, 7, 'lutff_4/in_1')
// (11, 7, 'neigh_op_bnl_5')
// (11, 7, 'sp4_v_b_30')
// (11, 7, 'sp4_v_b_37')
// (11, 8, 'local_g1_3')
// (11, 8, 'lutff_2/in_0')
// (11, 8, 'lutff_7/in_3')
// (11, 8, 'sp4_v_b_19')
// (11, 8, 'sp4_v_b_24')
// (11, 9, 'local_g1_6')
// (11, 9, 'lutff_4/in_3')
// (11, 9, 'sp4_v_b_13')
// (11, 9, 'sp4_v_b_6')
// (11, 9, 'sp4_v_t_39')
// (11, 10, 'sp4_v_b_0')
// (11, 10, 'sp4_v_b_39')
// (11, 10, 'sp4_v_t_38')
// (11, 11, 'sp4_v_b_26')
// (11, 11, 'sp4_v_b_38')
// (11, 12, 'sp4_v_b_15')
// (11, 12, 'sp4_v_b_27')
// (11, 13, 'sp4_v_b_14')
// (11, 13, 'sp4_v_b_2')
// (11, 14, 'local_g1_3')
// (11, 14, 'lutff_5/in_3')
// (11, 14, 'sp4_v_b_3')

wire n985;
// (7, 6, 'sp4_r_v_b_47')
// (7, 7, 'sp4_r_v_b_34')
// (7, 8, 'neigh_op_tnr_5')
// (7, 8, 'sp4_r_v_b_23')
// (7, 9, 'neigh_op_rgt_5')
// (7, 9, 'sp4_r_v_b_10')
// (7, 10, 'neigh_op_bnr_5')
// (8, 5, 'sp4_v_t_47')
// (8, 6, 'sp4_v_b_47')
// (8, 7, 'local_g2_2')
// (8, 7, 'lutff_5/in_1')
// (8, 7, 'sp4_v_b_34')
// (8, 8, 'local_g1_5')
// (8, 8, 'lutff_7/in_3')
// (8, 8, 'neigh_op_top_5')
// (8, 8, 'sp4_v_b_23')
// (8, 9, 'lutff_5/out')
// (8, 9, 'sp4_v_b_10')
// (8, 10, 'neigh_op_bot_5')
// (9, 8, 'neigh_op_tnl_5')
// (9, 9, 'neigh_op_lft_5')
// (9, 10, 'neigh_op_bnl_5')

wire n986;
// (7, 7, 'local_g2_7')
// (7, 7, 'lutff_6/in_3')
// (7, 7, 'neigh_op_tnr_7')
// (7, 8, 'neigh_op_rgt_7')
// (7, 9, 'neigh_op_bnr_7')
// (8, 7, 'neigh_op_top_7')
// (8, 8, 'lutff_7/out')
// (8, 9, 'neigh_op_bot_7')
// (9, 7, 'neigh_op_tnl_7')
// (9, 8, 'neigh_op_lft_7')
// (9, 9, 'neigh_op_bnl_7')

wire n987;
// (7, 7, 'neigh_op_tnr_0')
// (7, 8, 'neigh_op_rgt_0')
// (7, 9, 'neigh_op_bnr_0')
// (8, 7, 'local_g1_0')
// (8, 7, 'lutff_2/in_1')
// (8, 7, 'neigh_op_top_0')
// (8, 8, 'lutff_0/out')
// (8, 9, 'neigh_op_bot_0')
// (9, 7, 'neigh_op_tnl_0')
// (9, 8, 'neigh_op_lft_0')
// (9, 9, 'neigh_op_bnl_0')

wire n988;
// (7, 7, 'neigh_op_tnr_3')
// (7, 8, 'neigh_op_rgt_3')
// (7, 9, 'neigh_op_bnr_3')
// (8, 7, 'local_g0_3')
// (8, 7, 'lutff_5/in_2')
// (8, 7, 'neigh_op_top_3')
// (8, 8, 'lutff_3/out')
// (8, 9, 'neigh_op_bot_3')
// (9, 7, 'neigh_op_tnl_3')
// (9, 8, 'neigh_op_lft_3')
// (9, 9, 'neigh_op_bnl_3')

reg n989 = 0;
// (7, 7, 'neigh_op_tnr_4')
// (7, 8, 'neigh_op_rgt_4')
// (7, 9, 'neigh_op_bnr_4')
// (8, 7, 'neigh_op_top_4')
// (8, 8, 'lutff_4/out')
// (8, 8, 'sp4_r_v_b_41')
// (8, 9, 'local_g1_4')
// (8, 9, 'lutff_4/in_1')
// (8, 9, 'neigh_op_bot_4')
// (8, 9, 'sp4_r_v_b_28')
// (8, 10, 'sp4_r_v_b_17')
// (8, 11, 'sp4_r_v_b_4')
// (9, 7, 'neigh_op_tnl_4')
// (9, 7, 'sp4_v_t_41')
// (9, 8, 'local_g0_4')
// (9, 8, 'lutff_6/in_2')
// (9, 8, 'neigh_op_lft_4')
// (9, 8, 'sp4_v_b_41')
// (9, 9, 'neigh_op_bnl_4')
// (9, 9, 'sp4_v_b_28')
// (9, 10, 'local_g1_1')
// (9, 10, 'lutff_5/in_1')
// (9, 10, 'sp4_v_b_17')
// (9, 11, 'sp4_v_b_4')

wire n990;
// (7, 7, 'neigh_op_tnr_6')
// (7, 8, 'neigh_op_rgt_6')
// (7, 9, 'neigh_op_bnr_6')
// (8, 7, 'local_g1_6')
// (8, 7, 'lutff_1/in_2')
// (8, 7, 'neigh_op_top_6')
// (8, 8, 'lutff_6/out')
// (8, 9, 'neigh_op_bot_6')
// (9, 7, 'neigh_op_tnl_6')
// (9, 8, 'neigh_op_lft_6')
// (9, 9, 'neigh_op_bnl_6')

wire n991;
// (7, 8, 'lutff_1/cout')
// (7, 8, 'lutff_2/in_3')

wire n992;
// (7, 8, 'lutff_2/cout')
// (7, 8, 'lutff_3/in_3')

wire n993;
// (7, 8, 'lutff_3/cout')
// (7, 8, 'lutff_4/in_3')

wire n994;
// (7, 8, 'lutff_4/cout')
// (7, 8, 'lutff_5/in_3')

wire n995;
// (7, 8, 'lutff_5/cout')
// (7, 8, 'lutff_6/in_3')

wire n996;
// (7, 8, 'neigh_op_tnr_1')
// (7, 9, 'local_g2_1')
// (7, 9, 'lutff_1/in_2')
// (7, 9, 'neigh_op_rgt_1')
// (7, 10, 'neigh_op_bnr_1')
// (8, 8, 'neigh_op_top_1')
// (8, 9, 'lutff_1/out')
// (8, 10, 'neigh_op_bot_1')
// (9, 8, 'neigh_op_tnl_1')
// (9, 9, 'neigh_op_lft_1')
// (9, 10, 'neigh_op_bnl_1')

wire n997;
// (7, 8, 'neigh_op_tnr_2')
// (7, 9, 'local_g2_2')
// (7, 9, 'lutff_2/in_2')
// (7, 9, 'neigh_op_rgt_2')
// (7, 10, 'neigh_op_bnr_2')
// (8, 8, 'neigh_op_top_2')
// (8, 9, 'lutff_2/out')
// (8, 10, 'neigh_op_bot_2')
// (9, 8, 'neigh_op_tnl_2')
// (9, 9, 'neigh_op_lft_2')
// (9, 10, 'neigh_op_bnl_2')

wire n998;
// (7, 8, 'neigh_op_tnr_3')
// (7, 9, 'local_g3_3')
// (7, 9, 'lutff_3/in_1')
// (7, 9, 'neigh_op_rgt_3')
// (7, 10, 'neigh_op_bnr_3')
// (8, 8, 'neigh_op_top_3')
// (8, 9, 'lutff_3/out')
// (8, 10, 'neigh_op_bot_3')
// (9, 8, 'neigh_op_tnl_3')
// (9, 9, 'neigh_op_lft_3')
// (9, 10, 'neigh_op_bnl_3')

wire n999;
// (7, 8, 'neigh_op_tnr_4')
// (7, 9, 'local_g3_4')
// (7, 9, 'lutff_4/in_1')
// (7, 9, 'neigh_op_rgt_4')
// (7, 10, 'neigh_op_bnr_4')
// (8, 8, 'neigh_op_top_4')
// (8, 9, 'lutff_4/out')
// (8, 10, 'neigh_op_bot_4')
// (9, 8, 'neigh_op_tnl_4')
// (9, 9, 'neigh_op_lft_4')
// (9, 10, 'neigh_op_bnl_4')

reg n1000 = 0;
// (7, 8, 'neigh_op_tnr_6')
// (7, 9, 'neigh_op_rgt_6')
// (7, 9, 'sp4_h_r_1')
// (7, 10, 'neigh_op_bnr_6')
// (8, 8, 'neigh_op_top_6')
// (8, 9, 'local_g0_6')
// (8, 9, 'lutff_5/in_1')
// (8, 9, 'lutff_6/out')
// (8, 9, 'sp4_h_r_12')
// (8, 10, 'neigh_op_bot_6')
// (9, 8, 'neigh_op_tnl_6')
// (9, 9, 'neigh_op_lft_6')
// (9, 9, 'sp4_h_r_25')
// (9, 10, 'neigh_op_bnl_6')
// (10, 9, 'local_g2_4')
// (10, 9, 'lutff_5/in_3')
// (10, 9, 'lutff_6/in_2')
// (10, 9, 'sp4_h_r_36')
// (11, 9, 'sp4_h_l_36')

wire n1001;
// (7, 8, 'sp4_r_v_b_47')
// (7, 9, 'sp4_r_v_b_34')
// (7, 10, 'local_g3_7')
// (7, 10, 'lutff_5/in_1')
// (7, 10, 'sp4_r_v_b_23')
// (7, 11, 'sp4_r_v_b_10')
// (8, 7, 'sp4_h_r_10')
// (8, 7, 'sp4_v_t_47')
// (8, 8, 'sp4_v_b_47')
// (8, 9, 'sp4_v_b_34')
// (8, 10, 'local_g1_7')
// (8, 10, 'lutff_2/in_2')
// (8, 10, 'sp4_v_b_23')
// (8, 11, 'sp4_v_b_10')
// (9, 7, 'sp4_h_r_23')
// (10, 5, 'sp4_h_r_11')
// (10, 7, 'sp4_h_r_34')
// (11, 4, 'local_g1_5')
// (11, 4, 'lutff_7/in_3')
// (11, 4, 'sp4_h_r_5')
// (11, 5, 'sp4_h_r_22')
// (11, 7, 'sp4_h_r_47')
// (12, 4, 'sp4_h_r_16')
// (12, 5, 'local_g2_3')
// (12, 5, 'lutff_7/in_0')
// (12, 5, 'sp4_h_r_35')
// (12, 7, 'sp4_h_l_47')
// (12, 7, 'sp4_h_r_7')
// (13, 2, 'sp4_r_v_b_45')
// (13, 3, 'sp4_r_v_b_32')
// (13, 4, 'sp4_h_r_29')
// (13, 4, 'sp4_r_v_b_21')
// (13, 5, 'sp4_h_r_46')
// (13, 5, 'sp4_r_v_b_8')
// (13, 7, 'sp4_h_r_18')
// (14, 1, 'sp4_v_t_45')
// (14, 2, 'local_g3_5')
// (14, 2, 'lutff_2/in_0')
// (14, 2, 'sp4_v_b_45')
// (14, 3, 'sp4_v_b_32')
// (14, 4, 'neigh_op_tnr_7')
// (14, 4, 'sp4_h_r_40')
// (14, 4, 'sp4_v_b_21')
// (14, 5, 'neigh_op_rgt_7')
// (14, 5, 'sp4_h_l_46')
// (14, 5, 'sp4_h_r_3')
// (14, 5, 'sp4_r_v_b_46')
// (14, 5, 'sp4_v_b_8')
// (14, 6, 'neigh_op_bnr_7')
// (14, 6, 'sp4_r_v_b_35')
// (14, 7, 'sp4_h_r_31')
// (14, 7, 'sp4_r_v_b_22')
// (14, 8, 'sp4_r_v_b_11')
// (15, 4, 'neigh_op_top_7')
// (15, 4, 'sp4_h_l_40')
// (15, 4, 'sp4_r_v_b_42')
// (15, 4, 'sp4_v_t_46')
// (15, 5, 'lutff_7/out')
// (15, 5, 'sp4_h_r_14')
// (15, 5, 'sp4_r_v_b_31')
// (15, 5, 'sp4_v_b_46')
// (15, 6, 'neigh_op_bot_7')
// (15, 6, 'sp4_r_v_b_18')
// (15, 6, 'sp4_v_b_35')
// (15, 7, 'sp4_h_r_42')
// (15, 7, 'sp4_r_v_b_7')
// (15, 7, 'sp4_v_b_22')
// (15, 8, 'sp4_v_b_11')
// (16, 3, 'sp4_v_t_42')
// (16, 4, 'neigh_op_tnl_7')
// (16, 4, 'sp4_v_b_42')
// (16, 5, 'neigh_op_lft_7')
// (16, 5, 'sp4_h_r_27')
// (16, 5, 'sp4_v_b_31')
// (16, 6, 'neigh_op_bnl_7')
// (16, 6, 'sp4_v_b_18')
// (16, 7, 'sp4_h_l_42')
// (16, 7, 'sp4_v_b_7')
// (17, 5, 'sp4_h_r_38')
// (18, 5, 'sp4_h_l_38')

wire n1002;
// (7, 9, 'lutff_1/cout')
// (7, 9, 'lutff_2/in_3')

wire n1003;
// (7, 9, 'lutff_2/cout')
// (7, 9, 'lutff_3/in_3')

wire n1004;
// (7, 9, 'lutff_3/cout')
// (7, 9, 'lutff_4/in_3')

wire n1005;
// (7, 9, 'lutff_4/cout')
// (7, 9, 'lutff_5/in_3')

reg n1006 = 0;
// (7, 9, 'neigh_op_tnr_0')
// (7, 10, 'neigh_op_rgt_0')
// (7, 11, 'neigh_op_bnr_0')
// (8, 9, 'neigh_op_top_0')
// (8, 10, 'local_g3_0')
// (8, 10, 'lutff_0/out')
// (8, 10, 'lutff_6/in_3')
// (8, 11, 'neigh_op_bot_0')
// (9, 9, 'neigh_op_tnl_0')
// (9, 10, 'neigh_op_lft_0')
// (9, 11, 'neigh_op_bnl_0')

reg n1007 = 0;
// (7, 9, 'neigh_op_tnr_1')
// (7, 10, 'neigh_op_rgt_1')
// (7, 11, 'neigh_op_bnr_1')
// (8, 9, 'neigh_op_top_1')
// (8, 10, 'lutff_1/out')
// (8, 11, 'neigh_op_bot_1')
// (9, 9, 'neigh_op_tnl_1')
// (9, 10, 'local_g0_1')
// (9, 10, 'lutff_2/in_1')
// (9, 10, 'neigh_op_lft_1')
// (9, 11, 'neigh_op_bnl_1')

reg n1008 = 0;
// (7, 9, 'neigh_op_tnr_3')
// (7, 10, 'neigh_op_rgt_3')
// (7, 11, 'neigh_op_bnr_3')
// (8, 9, 'neigh_op_top_3')
// (8, 10, 'lutff_3/out')
// (8, 11, 'neigh_op_bot_3')
// (9, 9, 'neigh_op_tnl_3')
// (9, 10, 'local_g0_3')
// (9, 10, 'lutff_4/in_3')
// (9, 10, 'neigh_op_lft_3')
// (9, 11, 'neigh_op_bnl_3')

reg n1009 = 0;
// (7, 9, 'neigh_op_tnr_4')
// (7, 10, 'neigh_op_rgt_4')
// (7, 11, 'neigh_op_bnr_4')
// (8, 9, 'neigh_op_top_4')
// (8, 10, 'local_g0_4')
// (8, 10, 'lutff_4/out')
// (8, 10, 'lutff_6/in_0')
// (8, 11, 'neigh_op_bot_4')
// (9, 9, 'neigh_op_tnl_4')
// (9, 10, 'neigh_op_lft_4')
// (9, 11, 'neigh_op_bnl_4')

wire n1010;
// (7, 9, 'neigh_op_tnr_6')
// (7, 10, 'neigh_op_rgt_6')
// (7, 10, 'sp4_h_r_1')
// (7, 11, 'neigh_op_bnr_6')
// (8, 9, 'neigh_op_top_6')
// (8, 10, 'lutff_6/out')
// (8, 10, 'sp4_h_r_12')
// (8, 11, 'neigh_op_bot_6')
// (9, 9, 'neigh_op_tnl_6')
// (9, 10, 'neigh_op_lft_6')
// (9, 10, 'sp4_h_r_25')
// (9, 11, 'neigh_op_bnl_6')
// (10, 10, 'local_g3_4')
// (10, 10, 'lutff_3/in_2')
// (10, 10, 'sp4_h_r_36')
// (11, 10, 'sp4_h_l_36')

reg n1011 = 0;
// (7, 9, 'neigh_op_tnr_7')
// (7, 10, 'neigh_op_rgt_7')
// (7, 11, 'neigh_op_bnr_7')
// (8, 9, 'neigh_op_top_7')
// (8, 10, 'lutff_7/out')
// (8, 11, 'local_g1_7')
// (8, 11, 'lutff_5/in_3')
// (8, 11, 'neigh_op_bot_7')
// (9, 9, 'neigh_op_tnl_7')
// (9, 10, 'neigh_op_lft_7')
// (9, 11, 'neigh_op_bnl_7')

reg n1012 = 0;
// (7, 10, 'neigh_op_tnr_0')
// (7, 11, 'neigh_op_rgt_0')
// (7, 12, 'neigh_op_bnr_0')
// (8, 10, 'neigh_op_top_0')
// (8, 11, 'local_g3_0')
// (8, 11, 'lutff_0/out')
// (8, 11, 'lutff_5/in_0')
// (8, 12, 'neigh_op_bot_0')
// (9, 10, 'neigh_op_tnl_0')
// (9, 11, 'neigh_op_lft_0')
// (9, 12, 'neigh_op_bnl_0')

reg n1013 = 0;
// (7, 10, 'neigh_op_tnr_1')
// (7, 11, 'neigh_op_rgt_1')
// (7, 12, 'neigh_op_bnr_1')
// (8, 10, 'neigh_op_top_1')
// (8, 10, 'sp4_r_v_b_46')
// (8, 11, 'lutff_1/out')
// (8, 11, 'sp4_r_v_b_35')
// (8, 12, 'neigh_op_bot_1')
// (8, 12, 'sp4_r_v_b_22')
// (8, 13, 'local_g2_3')
// (8, 13, 'lutff_4/in_1')
// (8, 13, 'sp4_r_v_b_11')
// (9, 9, 'sp4_v_t_46')
// (9, 10, 'neigh_op_tnl_1')
// (9, 10, 'sp4_v_b_46')
// (9, 11, 'neigh_op_lft_1')
// (9, 11, 'sp4_v_b_35')
// (9, 12, 'neigh_op_bnl_1')
// (9, 12, 'sp4_v_b_22')
// (9, 13, 'sp4_v_b_11')

reg n1014 = 0;
// (7, 10, 'neigh_op_tnr_2')
// (7, 11, 'neigh_op_rgt_2')
// (7, 12, 'neigh_op_bnr_2')
// (8, 10, 'neigh_op_top_2')
// (8, 11, 'local_g1_2')
// (8, 11, 'lutff_2/out')
// (8, 11, 'lutff_4/in_1')
// (8, 12, 'neigh_op_bot_2')
// (9, 10, 'neigh_op_tnl_2')
// (9, 11, 'neigh_op_lft_2')
// (9, 12, 'neigh_op_bnl_2')

reg n1015 = 0;
// (7, 10, 'neigh_op_tnr_3')
// (7, 11, 'neigh_op_rgt_3')
// (7, 12, 'neigh_op_bnr_3')
// (8, 10, 'neigh_op_top_3')
// (8, 11, 'local_g3_3')
// (8, 11, 'lutff_3/out')
// (8, 11, 'lutff_4/in_0')
// (8, 12, 'neigh_op_bot_3')
// (9, 10, 'neigh_op_tnl_3')
// (9, 11, 'neigh_op_lft_3')
// (9, 12, 'neigh_op_bnl_3')

wire n1016;
// (7, 10, 'neigh_op_tnr_4')
// (7, 11, 'neigh_op_rgt_4')
// (7, 12, 'neigh_op_bnr_4')
// (8, 10, 'neigh_op_top_4')
// (8, 11, 'local_g0_4')
// (8, 11, 'lutff_4/out')
// (8, 11, 'lutff_5/in_1')
// (8, 12, 'neigh_op_bot_4')
// (9, 10, 'neigh_op_tnl_4')
// (9, 11, 'neigh_op_lft_4')
// (9, 12, 'neigh_op_bnl_4')

wire n1017;
// (7, 10, 'neigh_op_tnr_5')
// (7, 11, 'neigh_op_rgt_5')
// (7, 12, 'neigh_op_bnr_5')
// (8, 10, 'neigh_op_top_5')
// (8, 11, 'lutff_5/out')
// (8, 11, 'sp4_r_v_b_43')
// (8, 12, 'neigh_op_bot_5')
// (8, 12, 'sp4_r_v_b_30')
// (8, 13, 'sp4_r_v_b_19')
// (8, 14, 'sp4_r_v_b_6')
// (9, 10, 'neigh_op_tnl_5')
// (9, 10, 'sp4_v_t_43')
// (9, 11, 'neigh_op_lft_5')
// (9, 11, 'sp4_v_b_43')
// (9, 12, 'neigh_op_bnl_5')
// (9, 12, 'sp4_v_b_30')
// (9, 13, 'sp4_v_b_19')
// (9, 14, 'local_g0_6')
// (9, 14, 'lutff_1/in_1')
// (9, 14, 'sp4_v_b_6')

reg n1018 = 0;
// (7, 10, 'neigh_op_tnr_6')
// (7, 11, 'neigh_op_rgt_6')
// (7, 12, 'neigh_op_bnr_6')
// (8, 10, 'neigh_op_top_6')
// (8, 11, 'local_g3_6')
// (8, 11, 'lutff_4/in_3')
// (8, 11, 'lutff_6/out')
// (8, 12, 'neigh_op_bot_6')
// (9, 10, 'neigh_op_tnl_6')
// (9, 11, 'neigh_op_lft_6')
// (9, 12, 'neigh_op_bnl_6')

reg n1019 = 0;
// (7, 10, 'sp4_r_v_b_43')
// (7, 11, 'sp4_r_v_b_30')
// (7, 12, 'sp4_r_v_b_19')
// (7, 13, 'local_g1_6')
// (7, 13, 'lutff_0/in_3')
// (7, 13, 'sp4_r_v_b_6')
// (7, 14, 'sp4_r_v_b_36')
// (7, 14, 'sp4_r_v_b_47')
// (7, 15, 'sp4_r_v_b_25')
// (7, 15, 'sp4_r_v_b_34')
// (7, 16, 'sp4_r_v_b_12')
// (7, 16, 'sp4_r_v_b_23')
// (7, 17, 'sp4_r_v_b_1')
// (7, 17, 'sp4_r_v_b_10')
// (7, 18, 'sp4_r_v_b_47')
// (7, 19, 'sp4_r_v_b_34')
// (7, 20, 'neigh_op_tnr_5')
// (7, 20, 'sp4_r_v_b_23')
// (7, 21, 'neigh_op_rgt_5')
// (7, 21, 'sp4_r_v_b_10')
// (7, 22, 'neigh_op_bnr_5')
// (8, 9, 'sp4_v_t_43')
// (8, 10, 'sp4_v_b_43')
// (8, 11, 'sp4_v_b_30')
// (8, 12, 'sp4_v_b_19')
// (8, 13, 'local_g1_1')
// (8, 13, 'lutff_6/in_2')
// (8, 13, 'sp4_h_r_1')
// (8, 13, 'sp4_v_b_6')
// (8, 13, 'sp4_v_t_36')
// (8, 13, 'sp4_v_t_47')
// (8, 14, 'sp4_v_b_36')
// (8, 14, 'sp4_v_b_47')
// (8, 15, 'sp4_v_b_25')
// (8, 15, 'sp4_v_b_34')
// (8, 16, 'local_g1_7')
// (8, 16, 'lutff_5/in_1')
// (8, 16, 'sp4_v_b_12')
// (8, 16, 'sp4_v_b_23')
// (8, 17, 'sp4_v_b_1')
// (8, 17, 'sp4_v_b_10')
// (8, 17, 'sp4_v_t_47')
// (8, 18, 'sp4_v_b_47')
// (8, 19, 'sp4_v_b_34')
// (8, 20, 'neigh_op_top_5')
// (8, 20, 'sp4_r_v_b_38')
// (8, 20, 'sp4_v_b_23')
// (8, 21, 'lutff_5/out')
// (8, 21, 'sp4_r_v_b_27')
// (8, 21, 'sp4_v_b_10')
// (8, 22, 'local_g1_5')
// (8, 22, 'lutff_3/in_1')
// (8, 22, 'neigh_op_bot_5')
// (8, 22, 'sp4_r_v_b_14')
// (8, 23, 'sp4_r_v_b_3')
// (9, 13, 'sp4_h_r_12')
// (9, 19, 'local_g1_3')
// (9, 19, 'lutff_3/in_3')
// (9, 19, 'sp4_h_r_3')
// (9, 19, 'sp4_v_t_38')
// (9, 20, 'local_g2_5')
// (9, 20, 'lutff_3/in_2')
// (9, 20, 'neigh_op_tnl_5')
// (9, 20, 'sp4_v_b_38')
// (9, 21, 'neigh_op_lft_5')
// (9, 21, 'sp4_v_b_27')
// (9, 22, 'local_g3_5')
// (9, 22, 'lutff_0/in_2')
// (9, 22, 'lutff_1/in_3')
// (9, 22, 'neigh_op_bnl_5')
// (9, 22, 'sp4_v_b_14')
// (9, 23, 'sp4_v_b_3')
// (10, 13, 'sp4_h_r_25')
// (10, 19, 'sp4_h_r_14')
// (11, 13, 'sp4_h_r_36')
// (11, 19, 'sp4_h_r_27')
// (12, 13, 'sp4_h_l_36')
// (12, 19, 'sp4_h_r_38')
// (13, 19, 'sp4_h_l_38')

reg n1020 = 0;
// (7, 11, 'local_g2_4')
// (7, 11, 'lutff_0/in_2')
// (7, 11, 'neigh_op_tnr_4')
// (7, 12, 'neigh_op_rgt_4')
// (7, 12, 'sp4_r_v_b_40')
// (7, 13, 'neigh_op_bnr_4')
// (7, 13, 'sp4_r_v_b_29')
// (7, 14, 'sp4_r_v_b_16')
// (7, 15, 'local_g1_5')
// (7, 15, 'lutff_3/in_1')
// (7, 15, 'sp4_r_v_b_5')
// (8, 11, 'neigh_op_top_4')
// (8, 11, 'sp4_v_t_40')
// (8, 12, 'lutff_4/out')
// (8, 12, 'sp4_r_v_b_41')
// (8, 12, 'sp4_v_b_40')
// (8, 13, 'local_g1_4')
// (8, 13, 'lutff_6/in_3')
// (8, 13, 'neigh_op_bot_4')
// (8, 13, 'sp4_r_v_b_28')
// (8, 13, 'sp4_v_b_29')
// (8, 14, 'local_g3_1')
// (8, 14, 'lutff_3/in_3')
// (8, 14, 'sp4_r_v_b_17')
// (8, 14, 'sp4_v_b_16')
// (8, 15, 'local_g1_5')
// (8, 15, 'lutff_3/in_1')
// (8, 15, 'sp4_r_v_b_4')
// (8, 15, 'sp4_v_b_5')
// (9, 11, 'neigh_op_tnl_4')
// (9, 11, 'sp4_v_t_41')
// (9, 12, 'neigh_op_lft_4')
// (9, 12, 'sp4_v_b_41')
// (9, 13, 'neigh_op_bnl_4')
// (9, 13, 'sp4_v_b_28')
// (9, 14, 'sp4_v_b_17')
// (9, 15, 'sp4_v_b_4')

reg n1021 = 0;
// (7, 11, 'neigh_op_tnr_2')
// (7, 12, 'neigh_op_rgt_2')
// (7, 12, 'sp4_r_v_b_36')
// (7, 13, 'neigh_op_bnr_2')
// (7, 13, 'sp4_r_v_b_25')
// (7, 14, 'sp4_r_v_b_12')
// (7, 15, 'local_g1_1')
// (7, 15, 'lutff_7/in_1')
// (7, 15, 'sp4_r_v_b_1')
// (8, 9, 'sp4_r_v_b_40')
// (8, 10, 'sp4_r_v_b_29')
// (8, 11, 'neigh_op_top_2')
// (8, 11, 'sp4_r_v_b_16')
// (8, 11, 'sp4_v_t_36')
// (8, 12, 'lutff_2/out')
// (8, 12, 'sp4_r_v_b_37')
// (8, 12, 'sp4_r_v_b_5')
// (8, 12, 'sp4_v_b_36')
// (8, 13, 'local_g1_2')
// (8, 13, 'lutff_6/in_1')
// (8, 13, 'neigh_op_bot_2')
// (8, 13, 'sp4_r_v_b_24')
// (8, 13, 'sp4_v_b_25')
// (8, 14, 'sp4_r_v_b_13')
// (8, 14, 'sp4_v_b_12')
// (8, 15, 'local_g1_1')
// (8, 15, 'lutff_7/in_1')
// (8, 15, 'sp4_r_v_b_0')
// (8, 15, 'sp4_v_b_1')
// (9, 8, 'sp4_v_t_40')
// (9, 9, 'sp4_v_b_40')
// (9, 10, 'local_g2_5')
// (9, 10, 'lutff_1/in_0')
// (9, 10, 'sp4_v_b_29')
// (9, 11, 'neigh_op_tnl_2')
// (9, 11, 'sp4_v_b_16')
// (9, 11, 'sp4_v_t_37')
// (9, 12, 'neigh_op_lft_2')
// (9, 12, 'sp4_v_b_37')
// (9, 12, 'sp4_v_b_5')
// (9, 13, 'neigh_op_bnl_2')
// (9, 13, 'sp4_v_b_24')
// (9, 14, 'sp4_v_b_13')
// (9, 15, 'local_g1_0')
// (9, 15, 'lutff_4/in_1')
// (9, 15, 'sp4_v_b_0')

reg n1022 = 0;
// (7, 11, 'neigh_op_tnr_7')
// (7, 12, 'neigh_op_rgt_7')
// (7, 12, 'sp4_r_v_b_46')
// (7, 13, 'neigh_op_bnr_7')
// (7, 13, 'sp4_r_v_b_35')
// (7, 14, 'sp4_r_v_b_22')
// (7, 15, 'local_g2_3')
// (7, 15, 'lutff_6/in_1')
// (7, 15, 'sp4_r_v_b_11')
// (8, 10, 'sp4_r_v_b_39')
// (8, 11, 'neigh_op_top_7')
// (8, 11, 'sp4_r_v_b_26')
// (8, 11, 'sp4_r_v_b_42')
// (8, 11, 'sp4_v_t_46')
// (8, 12, 'lutff_7/out')
// (8, 12, 'sp4_r_v_b_15')
// (8, 12, 'sp4_r_v_b_31')
// (8, 12, 'sp4_r_v_b_47')
// (8, 12, 'sp4_v_b_46')
// (8, 13, 'neigh_op_bot_7')
// (8, 13, 'sp4_r_v_b_18')
// (8, 13, 'sp4_r_v_b_2')
// (8, 13, 'sp4_r_v_b_34')
// (8, 13, 'sp4_v_b_35')
// (8, 14, 'local_g1_7')
// (8, 14, 'lutff_6/in_2')
// (8, 14, 'sp4_r_v_b_23')
// (8, 14, 'sp4_r_v_b_7')
// (8, 14, 'sp4_v_b_22')
// (8, 15, 'local_g0_3')
// (8, 15, 'lutff_6/in_1')
// (8, 15, 'sp4_r_v_b_10')
// (8, 15, 'sp4_v_b_11')
// (9, 9, 'sp4_v_t_39')
// (9, 10, 'local_g2_7')
// (9, 10, 'lutff_3/in_0')
// (9, 10, 'sp4_v_b_39')
// (9, 10, 'sp4_v_t_42')
// (9, 11, 'neigh_op_tnl_7')
// (9, 11, 'sp4_v_b_26')
// (9, 11, 'sp4_v_b_42')
// (9, 11, 'sp4_v_t_47')
// (9, 12, 'neigh_op_lft_7')
// (9, 12, 'sp4_v_b_15')
// (9, 12, 'sp4_v_b_31')
// (9, 12, 'sp4_v_b_47')
// (9, 13, 'neigh_op_bnl_7')
// (9, 13, 'sp4_v_b_18')
// (9, 13, 'sp4_v_b_2')
// (9, 13, 'sp4_v_b_34')
// (9, 14, 'sp4_v_b_23')
// (9, 14, 'sp4_v_b_7')
// (9, 15, 'local_g0_2')
// (9, 15, 'lutff_7/in_1')
// (9, 15, 'sp4_v_b_10')

reg n1023 = 0;
// (7, 11, 'sp4_r_v_b_44')
// (7, 12, 'neigh_op_tnr_2')
// (7, 12, 'sp4_r_v_b_33')
// (7, 13, 'neigh_op_rgt_2')
// (7, 13, 'sp4_r_v_b_20')
// (7, 13, 'sp4_r_v_b_36')
// (7, 14, 'neigh_op_bnr_2')
// (7, 14, 'sp4_r_v_b_25')
// (7, 14, 'sp4_r_v_b_9')
// (7, 15, 'local_g2_4')
// (7, 15, 'lutff_5/in_1')
// (7, 15, 'sp4_r_v_b_12')
// (7, 16, 'sp4_r_v_b_1')
// (8, 10, 'local_g0_1')
// (8, 10, 'lutff_4/in_1')
// (8, 10, 'sp4_h_r_9')
// (8, 10, 'sp4_v_t_44')
// (8, 11, 'sp4_v_b_44')
// (8, 12, 'neigh_op_top_2')
// (8, 12, 'sp4_v_b_33')
// (8, 12, 'sp4_v_t_36')
// (8, 13, 'lutff_2/out')
// (8, 13, 'sp4_r_v_b_37')
// (8, 13, 'sp4_v_b_20')
// (8, 13, 'sp4_v_b_36')
// (8, 14, 'local_g1_2')
// (8, 14, 'lutff_5/in_2')
// (8, 14, 'neigh_op_bot_2')
// (8, 14, 'sp4_r_v_b_24')
// (8, 14, 'sp4_v_b_25')
// (8, 14, 'sp4_v_b_9')
// (8, 15, 'local_g0_4')
// (8, 15, 'lutff_5/in_1')
// (8, 15, 'sp4_r_v_b_13')
// (8, 15, 'sp4_v_b_12')
// (8, 16, 'sp4_r_v_b_0')
// (8, 16, 'sp4_v_b_1')
// (9, 10, 'sp4_h_r_20')
// (9, 12, 'neigh_op_tnl_2')
// (9, 12, 'sp4_v_t_37')
// (9, 13, 'neigh_op_lft_2')
// (9, 13, 'sp4_v_b_37')
// (9, 14, 'neigh_op_bnl_2')
// (9, 14, 'sp4_v_b_24')
// (9, 15, 'local_g1_5')
// (9, 15, 'lutff_4/in_2')
// (9, 15, 'sp4_v_b_13')
// (9, 16, 'sp4_v_b_0')
// (10, 10, 'sp4_h_r_33')
// (11, 10, 'sp4_h_r_44')
// (12, 10, 'sp4_h_l_44')

wire n1024;
// (7, 12, 'local_g0_2')
// (7, 12, 'lutff_6/in_2')
// (7, 12, 'sp4_h_r_10')
// (8, 11, 'neigh_op_tnr_1')
// (8, 12, 'neigh_op_rgt_1')
// (8, 12, 'sp4_h_r_23')
// (8, 13, 'neigh_op_bnr_1')
// (9, 11, 'neigh_op_top_1')
// (9, 12, 'lutff_1/out')
// (9, 12, 'sp4_h_r_34')
// (9, 13, 'neigh_op_bot_1')
// (10, 11, 'neigh_op_tnl_1')
// (10, 12, 'neigh_op_lft_1')
// (10, 12, 'sp4_h_r_47')
// (10, 13, 'neigh_op_bnl_1')
// (11, 12, 'sp4_h_l_47')

reg n1025 = 0;
// (7, 12, 'neigh_op_tnr_0')
// (7, 12, 'sp4_r_v_b_45')
// (7, 13, 'local_g2_0')
// (7, 13, 'lutff_1/in_3')
// (7, 13, 'neigh_op_rgt_0')
// (7, 13, 'sp4_r_v_b_32')
// (7, 14, 'neigh_op_bnr_0')
// (7, 14, 'sp4_r_v_b_21')
// (7, 15, 'local_g2_0')
// (7, 15, 'lutff_4/in_2')
// (7, 15, 'sp4_r_v_b_8')
// (8, 11, 'sp4_v_t_45')
// (8, 12, 'neigh_op_top_0')
// (8, 12, 'sp4_v_b_45')
// (8, 13, 'lutff_0/out')
// (8, 13, 'sp4_v_b_32')
// (8, 14, 'local_g0_0')
// (8, 14, 'local_g1_0')
// (8, 14, 'lutff_1/in_2')
// (8, 14, 'lutff_5/in_1')
// (8, 14, 'neigh_op_bot_0')
// (8, 14, 'sp4_v_b_21')
// (8, 15, 'local_g1_0')
// (8, 15, 'lutff_4/in_1')
// (8, 15, 'sp4_v_b_8')
// (9, 12, 'neigh_op_tnl_0')
// (9, 13, 'neigh_op_lft_0')
// (9, 14, 'neigh_op_bnl_0')

reg n1026 = 0;
// (7, 12, 'neigh_op_tnr_3')
// (7, 13, 'neigh_op_rgt_3')
// (7, 13, 'sp4_r_v_b_38')
// (7, 14, 'neigh_op_bnr_3')
// (7, 14, 'sp4_r_v_b_27')
// (7, 15, 'local_g2_6')
// (7, 15, 'lutff_2/in_2')
// (7, 15, 'sp4_r_v_b_14')
// (7, 16, 'sp4_r_v_b_3')
// (8, 10, 'sp4_r_v_b_42')
// (8, 11, 'local_g0_7')
// (8, 11, 'lutff_3/in_2')
// (8, 11, 'sp4_r_v_b_31')
// (8, 12, 'neigh_op_top_3')
// (8, 12, 'sp4_r_v_b_18')
// (8, 12, 'sp4_v_t_38')
// (8, 13, 'lutff_3/out')
// (8, 13, 'sp4_r_v_b_7')
// (8, 13, 'sp4_v_b_38')
// (8, 14, 'local_g0_3')
// (8, 14, 'lutff_0/in_1')
// (8, 14, 'lutff_3/in_2')
// (8, 14, 'neigh_op_bot_3')
// (8, 14, 'sp4_v_b_27')
// (8, 15, 'local_g1_6')
// (8, 15, 'lutff_2/in_1')
// (8, 15, 'sp4_v_b_14')
// (8, 16, 'sp4_v_b_3')
// (9, 9, 'sp4_v_t_42')
// (9, 10, 'sp4_v_b_42')
// (9, 11, 'sp4_v_b_31')
// (9, 12, 'neigh_op_tnl_3')
// (9, 12, 'sp4_v_b_18')
// (9, 13, 'neigh_op_lft_3')
// (9, 13, 'sp4_v_b_7')
// (9, 14, 'neigh_op_bnl_3')

wire n1027;
// (7, 12, 'neigh_op_tnr_4')
// (7, 13, 'neigh_op_rgt_4')
// (7, 14, 'neigh_op_bnr_4')
// (8, 12, 'neigh_op_top_4')
// (8, 13, 'lutff_4/out')
// (8, 13, 'sp4_h_r_8')
// (8, 14, 'neigh_op_bot_4')
// (9, 12, 'neigh_op_tnl_4')
// (9, 13, 'neigh_op_lft_4')
// (9, 13, 'sp4_h_r_21')
// (9, 14, 'neigh_op_bnl_4')
// (10, 13, 'local_g3_0')
// (10, 13, 'lutff_0/in_1')
// (10, 13, 'sp4_h_r_32')
// (11, 13, 'sp4_h_r_45')
// (12, 13, 'sp4_h_l_45')

reg n1028 = 0;
// (7, 12, 'neigh_op_tnr_5')
// (7, 13, 'neigh_op_rgt_5')
// (7, 13, 'sp4_r_v_b_42')
// (7, 14, 'neigh_op_bnr_5')
// (7, 14, 'sp4_r_v_b_31')
// (7, 15, 'local_g3_2')
// (7, 15, 'lutff_0/in_1')
// (7, 15, 'sp4_r_v_b_18')
// (7, 16, 'sp4_r_v_b_7')
// (8, 12, 'neigh_op_top_5')
// (8, 12, 'sp4_v_t_42')
// (8, 13, 'lutff_5/out')
// (8, 13, 'sp4_r_v_b_43')
// (8, 13, 'sp4_v_b_42')
// (8, 14, 'local_g0_5')
// (8, 14, 'lutff_0/in_3')
// (8, 14, 'neigh_op_bot_5')
// (8, 14, 'sp4_r_v_b_30')
// (8, 14, 'sp4_v_b_31')
// (8, 15, 'local_g3_3')
// (8, 15, 'lutff_0/in_2')
// (8, 15, 'sp4_r_v_b_19')
// (8, 15, 'sp4_v_b_18')
// (8, 16, 'sp4_r_v_b_6')
// (8, 16, 'sp4_v_b_7')
// (9, 12, 'neigh_op_tnl_5')
// (9, 12, 'sp4_v_t_43')
// (9, 13, 'local_g0_5')
// (9, 13, 'lutff_7/in_0')
// (9, 13, 'neigh_op_lft_5')
// (9, 13, 'sp4_v_b_43')
// (9, 14, 'neigh_op_bnl_5')
// (9, 14, 'sp4_v_b_30')
// (9, 15, 'local_g0_3')
// (9, 15, 'lutff_7/in_2')
// (9, 15, 'sp4_v_b_19')
// (9, 16, 'sp4_v_b_6')

wire n1029;
// (7, 12, 'neigh_op_tnr_6')
// (7, 13, 'neigh_op_rgt_6')
// (7, 14, 'neigh_op_bnr_6')
// (8, 12, 'neigh_op_top_6')
// (8, 13, 'lutff_6/out')
// (8, 14, 'local_g1_6')
// (8, 14, 'lutff_6/in_1')
// (8, 14, 'neigh_op_bot_6')
// (9, 12, 'neigh_op_tnl_6')
// (9, 13, 'neigh_op_lft_6')
// (9, 14, 'neigh_op_bnl_6')

wire n1030;
// (7, 12, 'neigh_op_tnr_7')
// (7, 13, 'neigh_op_rgt_7')
// (7, 14, 'neigh_op_bnr_7')
// (8, 12, 'neigh_op_top_7')
// (8, 13, 'local_g3_7')
// (8, 13, 'lutff_4/in_0')
// (8, 13, 'lutff_7/out')
// (8, 14, 'neigh_op_bot_7')
// (9, 12, 'neigh_op_tnl_7')
// (9, 13, 'neigh_op_lft_7')
// (9, 14, 'neigh_op_bnl_7')

wire n1031;
// (7, 12, 'sp12_h_r_0')
// (7, 12, 'sp12_v_t_23')
// (7, 13, 'sp12_v_b_23')
// (7, 14, 'sp12_v_b_20')
// (7, 15, 'sp12_v_b_19')
// (7, 16, 'sp12_v_b_16')
// (7, 17, 'sp12_v_b_15')
// (7, 18, 'sp12_v_b_12')
// (7, 19, 'sp12_v_b_11')
// (7, 20, 'sp12_v_b_8')
// (7, 21, 'local_g3_7')
// (7, 21, 'lutff_3/in_1')
// (7, 21, 'lutff_6/in_0')
// (7, 21, 'lutff_7/in_1')
// (7, 21, 'sp12_v_b_7')
// (7, 22, 'sp12_v_b_4')
// (7, 23, 'sp12_v_b_3')
// (7, 24, 'sp12_v_b_0')
// (8, 10, 'sp4_r_v_b_36')
// (8, 11, 'neigh_op_tnr_6')
// (8, 11, 'sp4_r_v_b_25')
// (8, 11, 'sp4_r_v_b_41')
// (8, 12, 'neigh_op_rgt_6')
// (8, 12, 'sp12_h_r_3')
// (8, 12, 'sp4_r_v_b_12')
// (8, 12, 'sp4_r_v_b_28')
// (8, 13, 'neigh_op_bnr_6')
// (8, 13, 'sp4_r_v_b_1')
// (8, 13, 'sp4_r_v_b_17')
// (8, 14, 'sp4_r_v_b_36')
// (8, 14, 'sp4_r_v_b_4')
// (8, 15, 'sp4_r_v_b_25')
// (8, 15, 'sp4_r_v_b_41')
// (8, 16, 'sp4_r_v_b_12')
// (8, 16, 'sp4_r_v_b_28')
// (8, 17, 'sp4_r_v_b_1')
// (8, 17, 'sp4_r_v_b_17')
// (8, 18, 'sp4_r_v_b_36')
// (8, 18, 'sp4_r_v_b_4')
// (8, 18, 'sp4_r_v_b_44')
// (8, 19, 'sp4_r_v_b_25')
// (8, 19, 'sp4_r_v_b_33')
// (8, 19, 'sp4_r_v_b_41')
// (8, 20, 'local_g2_4')
// (8, 20, 'local_g3_4')
// (8, 20, 'lutff_2/in_0')
// (8, 20, 'lutff_5/in_3')
// (8, 20, 'lutff_7/in_2')
// (8, 20, 'sp4_r_v_b_12')
// (8, 20, 'sp4_r_v_b_20')
// (8, 20, 'sp4_r_v_b_28')
// (8, 21, 'sp4_r_v_b_1')
// (8, 21, 'sp4_r_v_b_17')
// (8, 21, 'sp4_r_v_b_9')
// (8, 22, 'sp4_r_v_b_4')
// (9, 9, 'sp4_v_t_36')
// (9, 10, 'sp4_v_b_36')
// (9, 10, 'sp4_v_t_41')
// (9, 11, 'neigh_op_top_6')
// (9, 11, 'sp4_v_b_25')
// (9, 11, 'sp4_v_b_41')
// (9, 12, 'lutff_6/out')
// (9, 12, 'sp12_h_r_4')
// (9, 12, 'sp4_r_v_b_45')
// (9, 12, 'sp4_v_b_12')
// (9, 12, 'sp4_v_b_28')
// (9, 13, 'neigh_op_bot_6')
// (9, 13, 'sp4_r_v_b_32')
// (9, 13, 'sp4_v_b_1')
// (9, 13, 'sp4_v_b_17')
// (9, 13, 'sp4_v_t_36')
// (9, 14, 'sp4_r_v_b_21')
// (9, 14, 'sp4_v_b_36')
// (9, 14, 'sp4_v_b_4')
// (9, 14, 'sp4_v_t_41')
// (9, 15, 'sp4_r_v_b_8')
// (9, 15, 'sp4_v_b_25')
// (9, 15, 'sp4_v_b_41')
// (9, 16, 'sp4_r_v_b_45')
// (9, 16, 'sp4_v_b_12')
// (9, 16, 'sp4_v_b_28')
// (9, 17, 'sp4_r_v_b_32')
// (9, 17, 'sp4_v_b_1')
// (9, 17, 'sp4_v_b_17')
// (9, 17, 'sp4_v_t_36')
// (9, 17, 'sp4_v_t_44')
// (9, 18, 'sp4_r_v_b_21')
// (9, 18, 'sp4_v_b_36')
// (9, 18, 'sp4_v_b_4')
// (9, 18, 'sp4_v_b_44')
// (9, 18, 'sp4_v_t_41')
// (9, 19, 'sp4_r_v_b_8')
// (9, 19, 'sp4_v_b_25')
// (9, 19, 'sp4_v_b_33')
// (9, 19, 'sp4_v_b_41')
// (9, 20, 'sp4_v_b_12')
// (9, 20, 'sp4_v_b_20')
// (9, 20, 'sp4_v_b_28')
// (9, 21, 'local_g0_1')
// (9, 21, 'lutff_5/in_2')
// (9, 21, 'lutff_7/in_0')
// (9, 21, 'sp4_v_b_1')
// (9, 21, 'sp4_v_b_17')
// (9, 21, 'sp4_v_b_9')
// (9, 22, 'sp4_v_b_4')
// (10, 11, 'neigh_op_tnl_6')
// (10, 11, 'sp4_v_t_45')
// (10, 12, 'neigh_op_lft_6')
// (10, 12, 'sp12_h_r_7')
// (10, 12, 'sp4_v_b_45')
// (10, 13, 'neigh_op_bnl_6')
// (10, 13, 'sp4_v_b_32')
// (10, 14, 'sp4_v_b_21')
// (10, 15, 'sp4_v_b_8')
// (10, 15, 'sp4_v_t_45')
// (10, 16, 'sp4_v_b_45')
// (10, 17, 'sp4_v_b_32')
// (10, 18, 'sp4_v_b_21')
// (10, 19, 'local_g1_0')
// (10, 19, 'lutff_1/in_0')
// (10, 19, 'lutff_2/in_1')
// (10, 19, 'sp4_v_b_8')
// (11, 12, 'sp12_h_r_8')
// (12, 12, 'sp12_h_r_11')
// (13, 12, 'sp12_h_r_12')
// (14, 12, 'sp12_h_r_15')
// (15, 12, 'sp12_h_r_16')
// (16, 12, 'sp12_h_r_19')
// (17, 12, 'sp12_h_r_20')
// (18, 12, 'sp12_h_r_23')
// (19, 12, 'sp12_h_l_23')

reg n1032 = 0;
// (7, 12, 'sp4_h_r_0')
// (8, 12, 'sp4_h_r_13')
// (9, 12, 'local_g2_0')
// (9, 12, 'lutff_5/in_3')
// (9, 12, 'sp4_h_r_24')
// (10, 5, 'sp4_r_v_b_46')
// (10, 6, 'neigh_op_tnr_3')
// (10, 6, 'sp4_r_v_b_35')
// (10, 7, 'neigh_op_rgt_3')
// (10, 7, 'sp4_r_v_b_22')
// (10, 8, 'neigh_op_bnr_3')
// (10, 8, 'sp4_r_v_b_11')
// (10, 9, 'sp4_r_v_b_42')
// (10, 10, 'sp4_r_v_b_31')
// (10, 11, 'sp4_r_v_b_18')
// (10, 12, 'sp4_h_r_37')
// (10, 12, 'sp4_r_v_b_7')
// (11, 4, 'sp4_v_t_46')
// (11, 5, 'sp4_v_b_46')
// (11, 6, 'neigh_op_top_3')
// (11, 6, 'sp4_v_b_35')
// (11, 7, 'lutff_3/out')
// (11, 7, 'sp4_v_b_22')
// (11, 8, 'neigh_op_bot_3')
// (11, 8, 'sp4_v_b_11')
// (11, 8, 'sp4_v_t_42')
// (11, 9, 'sp4_v_b_42')
// (11, 10, 'sp4_v_b_31')
// (11, 11, 'sp4_v_b_18')
// (11, 12, 'sp4_h_l_37')
// (11, 12, 'sp4_v_b_7')
// (12, 6, 'neigh_op_tnl_3')
// (12, 7, 'neigh_op_lft_3')
// (12, 8, 'neigh_op_bnl_3')

wire n1033;
// (7, 12, 'sp4_r_v_b_42')
// (7, 13, 'sp4_r_v_b_31')
// (7, 14, 'local_g3_2')
// (7, 14, 'lutff_2/in_3')
// (7, 14, 'sp4_r_v_b_18')
// (7, 15, 'sp4_r_v_b_7')
// (8, 11, 'sp4_v_t_42')
// (8, 12, 'sp4_v_b_42')
// (8, 13, 'sp4_v_b_31')
// (8, 14, 'sp4_v_b_18')
// (8, 15, 'sp4_h_r_7')
// (8, 15, 'sp4_v_b_7')
// (9, 15, 'sp4_h_r_18')
// (10, 15, 'sp4_h_r_31')
// (11, 15, 'local_g2_2')
// (11, 15, 'lutff_0/in_2')
// (11, 15, 'lutff_6/in_0')
// (11, 15, 'neigh_op_tnr_2')
// (11, 15, 'sp4_h_r_42')
// (11, 16, 'neigh_op_rgt_2')
// (11, 16, 'sp4_r_v_b_36')
// (11, 17, 'neigh_op_bnr_2')
// (11, 17, 'sp4_r_v_b_25')
// (11, 18, 'sp4_r_v_b_12')
// (11, 19, 'sp4_r_v_b_1')
// (12, 15, 'neigh_op_top_2')
// (12, 15, 'sp4_h_l_42')
// (12, 15, 'sp4_v_t_36')
// (12, 16, 'lutff_2/out')
// (12, 16, 'sp4_v_b_36')
// (12, 17, 'local_g0_2')
// (12, 17, 'lutff_3/in_3')
// (12, 17, 'lutff_4/in_0')
// (12, 17, 'neigh_op_bot_2')
// (12, 17, 'sp4_v_b_25')
// (12, 18, 'sp4_v_b_12')
// (12, 19, 'sp4_v_b_1')
// (13, 15, 'neigh_op_tnl_2')
// (13, 16, 'neigh_op_lft_2')
// (13, 17, 'neigh_op_bnl_2')

wire n1034;
// (7, 12, 'sp4_r_v_b_44')
// (7, 13, 'sp4_r_v_b_33')
// (7, 14, 'sp4_r_v_b_20')
// (7, 15, 'sp4_r_v_b_9')
// (7, 16, 'sp4_r_v_b_36')
// (7, 17, 'neigh_op_tnr_6')
// (7, 17, 'sp4_r_v_b_25')
// (7, 18, 'local_g2_6')
// (7, 18, 'lutff_0/in_2')
// (7, 18, 'neigh_op_rgt_6')
// (7, 18, 'sp4_r_v_b_12')
// (7, 19, 'neigh_op_bnr_6')
// (7, 19, 'sp4_r_v_b_1')
// (8, 11, 'sp4_v_t_44')
// (8, 12, 'sp4_v_b_44')
// (8, 13, 'sp4_v_b_33')
// (8, 14, 'sp4_v_b_20')
// (8, 15, 'local_g0_1')
// (8, 15, 'lutff_0/in_1')
// (8, 15, 'sp4_v_b_9')
// (8, 15, 'sp4_v_t_36')
// (8, 16, 'sp4_v_b_36')
// (8, 17, 'local_g0_6')
// (8, 17, 'lutff_0/in_2')
// (8, 17, 'neigh_op_top_6')
// (8, 17, 'sp4_v_b_25')
// (8, 18, 'lutff_6/out')
// (8, 18, 'sp4_v_b_12')
// (8, 19, 'neigh_op_bot_6')
// (8, 19, 'sp4_v_b_1')
// (9, 17, 'neigh_op_tnl_6')
// (9, 18, 'local_g0_6')
// (9, 18, 'lutff_0/in_2')
// (9, 18, 'neigh_op_lft_6')
// (9, 19, 'neigh_op_bnl_6')

wire n1035;
// (7, 13, 'neigh_op_tnr_0')
// (7, 14, 'neigh_op_rgt_0')
// (7, 15, 'neigh_op_bnr_0')
// (8, 13, 'neigh_op_top_0')
// (8, 14, 'local_g3_0')
// (8, 14, 'lutff_0/out')
// (8, 14, 'lutff_6/in_3')
// (8, 15, 'neigh_op_bot_0')
// (9, 13, 'neigh_op_tnl_0')
// (9, 14, 'neigh_op_lft_0')
// (9, 15, 'neigh_op_bnl_0')

wire n1036;
// (7, 13, 'neigh_op_tnr_1')
// (7, 14, 'neigh_op_rgt_1')
// (7, 15, 'neigh_op_bnr_1')
// (8, 13, 'neigh_op_top_1')
// (8, 14, 'lutff_1/out')
// (8, 15, 'neigh_op_bot_1')
// (9, 13, 'neigh_op_tnl_1')
// (9, 14, 'neigh_op_lft_1')
// (9, 15, 'local_g2_1')
// (9, 15, 'lutff_0/in_1')
// (9, 15, 'neigh_op_bnl_1')

reg n1037 = 0;
// (7, 13, 'neigh_op_tnr_2')
// (7, 14, 'neigh_op_rgt_2')
// (7, 15, 'neigh_op_bnr_2')
// (8, 11, 'sp4_r_v_b_40')
// (8, 12, 'sp4_r_v_b_29')
// (8, 12, 'sp4_r_v_b_45')
// (8, 13, 'neigh_op_top_2')
// (8, 13, 'sp4_r_v_b_16')
// (8, 13, 'sp4_r_v_b_32')
// (8, 14, 'lutff_2/out')
// (8, 14, 'sp4_h_r_4')
// (8, 14, 'sp4_r_v_b_21')
// (8, 14, 'sp4_r_v_b_37')
// (8, 14, 'sp4_r_v_b_5')
// (8, 15, 'neigh_op_bot_2')
// (8, 15, 'sp4_r_v_b_24')
// (8, 15, 'sp4_r_v_b_8')
// (8, 16, 'sp4_r_v_b_13')
// (8, 17, 'sp4_r_v_b_0')
// (9, 10, 'sp4_h_r_10')
// (9, 10, 'sp4_h_r_5')
// (9, 10, 'sp4_v_t_40')
// (9, 11, 'sp4_v_b_40')
// (9, 11, 'sp4_v_t_45')
// (9, 12, 'sp4_v_b_29')
// (9, 12, 'sp4_v_b_45')
// (9, 13, 'neigh_op_tnl_2')
// (9, 13, 'sp4_h_r_5')
// (9, 13, 'sp4_v_b_16')
// (9, 13, 'sp4_v_b_32')
// (9, 13, 'sp4_v_t_37')
// (9, 14, 'neigh_op_lft_2')
// (9, 14, 'sp4_h_r_17')
// (9, 14, 'sp4_v_b_21')
// (9, 14, 'sp4_v_b_37')
// (9, 14, 'sp4_v_b_5')
// (9, 15, 'neigh_op_bnl_2')
// (9, 15, 'sp4_h_r_2')
// (9, 15, 'sp4_v_b_24')
// (9, 15, 'sp4_v_b_8')
// (9, 16, 'sp4_v_b_13')
// (9, 17, 'sp4_v_b_0')
// (10, 10, 'sp4_h_r_16')
// (10, 10, 'sp4_h_r_23')
// (10, 13, 'sp4_h_r_16')
// (10, 14, 'sp4_h_r_28')
// (10, 15, 'sp4_h_r_15')
// (11, 10, 'sp4_h_r_29')
// (11, 10, 'sp4_h_r_34')
// (11, 13, 'sp4_h_r_29')
// (11, 14, 'sp4_h_r_41')
// (11, 15, 'sp4_h_r_26')
// (12, 7, 'sp4_r_v_b_40')
// (12, 7, 'sp4_r_v_b_41')
// (12, 8, 'sp4_r_v_b_28')
// (12, 8, 'sp4_r_v_b_29')
// (12, 9, 'sp4_r_v_b_16')
// (12, 9, 'sp4_r_v_b_17')
// (12, 10, 'sp4_h_r_40')
// (12, 10, 'sp4_h_r_47')
// (12, 10, 'sp4_r_v_b_4')
// (12, 10, 'sp4_r_v_b_40')
// (12, 10, 'sp4_r_v_b_5')
// (12, 11, 'sp4_r_v_b_29')
// (12, 12, 'sp4_r_v_b_16')
// (12, 13, 'sp4_h_r_40')
// (12, 13, 'sp4_r_v_b_5')
// (12, 14, 'sp4_h_l_41')
// (12, 14, 'sp4_h_r_4')
// (12, 15, 'sp4_h_r_39')
// (13, 6, 'local_g0_4')
// (13, 6, 'lutff_1/in_1')
// (13, 6, 'lutff_2/in_0')
// (13, 6, 'sp4_h_r_4')
// (13, 6, 'sp4_v_t_40')
// (13, 6, 'sp4_v_t_41')
// (13, 7, 'local_g3_0')
// (13, 7, 'lutff_4/in_3')
// (13, 7, 'lutff_6/in_3')
// (13, 7, 'sp4_v_b_40')
// (13, 7, 'sp4_v_b_41')
// (13, 8, 'local_g2_4')
// (13, 8, 'lutff_1/in_3')
// (13, 8, 'sp4_v_b_28')
// (13, 8, 'sp4_v_b_29')
// (13, 9, 'sp4_v_b_16')
// (13, 9, 'sp4_v_b_17')
// (13, 9, 'sp4_v_t_40')
// (13, 10, 'sp4_h_l_40')
// (13, 10, 'sp4_h_l_47')
// (13, 10, 'sp4_v_b_4')
// (13, 10, 'sp4_v_b_40')
// (13, 10, 'sp4_v_b_5')
// (13, 11, 'sp4_v_b_29')
// (13, 12, 'local_g0_0')
// (13, 12, 'lutff_6/in_0')
// (13, 12, 'sp4_v_b_16')
// (13, 13, 'sp4_h_l_40')
// (13, 13, 'sp4_v_b_5')
// (13, 14, 'sp4_h_r_17')
// (13, 15, 'sp4_h_l_39')
// (13, 15, 'sp4_h_r_10')
// (14, 6, 'sp4_h_r_17')
// (14, 14, 'sp4_h_r_28')
// (14, 15, 'sp4_h_r_23')
// (15, 6, 'sp4_h_r_28')
// (15, 14, 'sp4_h_r_41')
// (15, 15, 'local_g3_2')
// (15, 15, 'lutff_5/in_2')
// (15, 15, 'sp4_h_r_34')
// (16, 6, 'sp4_h_r_41')
// (16, 14, 'local_g0_0')
// (16, 14, 'local_g1_0')
// (16, 14, 'lutff_6/in_3')
// (16, 14, 'lutff_7/in_1')
// (16, 14, 'sp4_h_l_41')
// (16, 14, 'sp4_h_r_0')
// (16, 15, 'sp4_h_r_47')
// (17, 6, 'sp4_h_l_41')
// (17, 14, 'sp4_h_r_13')
// (17, 15, 'sp4_h_l_47')
// (18, 14, 'sp4_h_r_24')
// (19, 14, 'sp4_h_r_37')
// (20, 14, 'sp4_h_l_37')

wire n1038;
// (7, 13, 'neigh_op_tnr_3')
// (7, 14, 'neigh_op_rgt_3')
// (7, 15, 'neigh_op_bnr_3')
// (8, 13, 'neigh_op_top_3')
// (8, 14, 'lutff_3/out')
// (8, 15, 'neigh_op_bot_3')
// (9, 13, 'neigh_op_tnl_3')
// (9, 14, 'neigh_op_lft_3')
// (9, 15, 'local_g3_3')
// (9, 15, 'lutff_0/in_0')
// (9, 15, 'neigh_op_bnl_3')

wire n1039;
// (7, 13, 'neigh_op_tnr_4')
// (7, 14, 'neigh_op_rgt_4')
// (7, 15, 'neigh_op_bnr_4')
// (8, 13, 'neigh_op_top_4')
// (8, 14, 'local_g3_4')
// (8, 14, 'lutff_4/out')
// (8, 14, 'lutff_7/in_2')
// (8, 15, 'neigh_op_bot_4')
// (9, 13, 'neigh_op_tnl_4')
// (9, 14, 'neigh_op_lft_4')
// (9, 15, 'neigh_op_bnl_4')

wire n1040;
// (7, 13, 'neigh_op_tnr_5')
// (7, 14, 'neigh_op_rgt_5')
// (7, 15, 'neigh_op_bnr_5')
// (8, 13, 'neigh_op_top_5')
// (8, 14, 'local_g1_5')
// (8, 14, 'lutff_4/in_0')
// (8, 14, 'lutff_5/out')
// (8, 15, 'neigh_op_bot_5')
// (9, 13, 'neigh_op_tnl_5')
// (9, 14, 'neigh_op_lft_5')
// (9, 15, 'neigh_op_bnl_5')

wire n1041;
// (7, 13, 'neigh_op_tnr_6')
// (7, 14, 'neigh_op_rgt_6')
// (7, 15, 'neigh_op_bnr_6')
// (8, 13, 'neigh_op_top_6')
// (8, 14, 'local_g2_6')
// (8, 14, 'lutff_6/out')
// (8, 14, 'lutff_7/in_3')
// (8, 15, 'neigh_op_bot_6')
// (9, 13, 'neigh_op_tnl_6')
// (9, 14, 'neigh_op_lft_6')
// (9, 15, 'neigh_op_bnl_6')

wire n1042;
// (7, 13, 'neigh_op_tnr_7')
// (7, 14, 'neigh_op_rgt_7')
// (7, 15, 'neigh_op_bnr_7')
// (8, 13, 'neigh_op_top_7')
// (8, 14, 'lutff_7/out')
// (8, 14, 'sp4_r_v_b_47')
// (8, 15, 'neigh_op_bot_7')
// (8, 15, 'sp4_r_v_b_34')
// (8, 16, 'local_g3_7')
// (8, 16, 'lutff_1/in_1')
// (8, 16, 'sp4_r_v_b_23')
// (8, 17, 'sp4_r_v_b_10')
// (9, 13, 'neigh_op_tnl_7')
// (9, 13, 'sp4_v_t_47')
// (9, 14, 'neigh_op_lft_7')
// (9, 14, 'sp4_v_b_47')
// (9, 15, 'neigh_op_bnl_7')
// (9, 15, 'sp4_v_b_34')
// (9, 16, 'sp4_v_b_23')
// (9, 17, 'sp4_v_b_10')

reg n1043 = 0;
// (7, 13, 'sp4_r_v_b_41')
// (7, 14, 'sp4_r_v_b_28')
// (7, 15, 'sp4_r_v_b_17')
// (7, 16, 'sp4_r_v_b_4')
// (7, 17, 'sp4_r_v_b_45')
// (7, 18, 'sp4_r_v_b_32')
// (7, 19, 'neigh_op_tnr_4')
// (7, 19, 'sp4_r_v_b_21')
// (7, 20, 'neigh_op_rgt_4')
// (7, 20, 'sp4_r_v_b_8')
// (7, 21, 'neigh_op_bnr_4')
// (8, 12, 'sp4_r_v_b_38')
// (8, 12, 'sp4_v_t_41')
// (8, 13, 'sp4_r_v_b_27')
// (8, 13, 'sp4_v_b_41')
// (8, 14, 'local_g2_4')
// (8, 14, 'lutff_0/in_2')
// (8, 14, 'sp4_r_v_b_14')
// (8, 14, 'sp4_v_b_28')
// (8, 15, 'sp4_r_v_b_3')
// (8, 15, 'sp4_v_b_17')
// (8, 16, 'local_g1_1')
// (8, 16, 'lutff_2/in_0')
// (8, 16, 'sp4_h_r_1')
// (8, 16, 'sp4_r_v_b_42')
// (8, 16, 'sp4_v_b_4')
// (8, 16, 'sp4_v_t_45')
// (8, 17, 'sp4_r_v_b_31')
// (8, 17, 'sp4_v_b_45')
// (8, 18, 'sp4_r_v_b_18')
// (8, 18, 'sp4_v_b_32')
// (8, 19, 'neigh_op_top_4')
// (8, 19, 'sp4_r_v_b_7')
// (8, 19, 'sp4_v_b_21')
// (8, 20, 'local_g0_4')
// (8, 20, 'lutff_4/in_2')
// (8, 20, 'lutff_4/out')
// (8, 20, 'lutff_6/in_0')
// (8, 20, 'sp4_r_v_b_41')
// (8, 20, 'sp4_v_b_8')
// (8, 21, 'neigh_op_bot_4')
// (8, 21, 'sp4_r_v_b_28')
// (8, 22, 'sp4_r_v_b_17')
// (8, 23, 'sp4_r_v_b_4')
// (9, 11, 'sp4_v_t_38')
// (9, 12, 'sp4_v_b_38')
// (9, 13, 'local_g3_3')
// (9, 13, 'lutff_4/in_0')
// (9, 13, 'sp4_v_b_27')
// (9, 14, 'sp4_v_b_14')
// (9, 15, 'sp4_v_b_3')
// (9, 15, 'sp4_v_t_42')
// (9, 16, 'sp4_h_r_12')
// (9, 16, 'sp4_v_b_42')
// (9, 17, 'sp4_v_b_31')
// (9, 18, 'sp4_v_b_18')
// (9, 19, 'local_g3_4')
// (9, 19, 'lutff_3/in_0')
// (9, 19, 'neigh_op_tnl_4')
// (9, 19, 'sp4_v_b_7')
// (9, 19, 'sp4_v_t_41')
// (9, 20, 'local_g1_4')
// (9, 20, 'lutff_0/in_1')
// (9, 20, 'neigh_op_lft_4')
// (9, 20, 'sp4_v_b_41')
// (9, 21, 'neigh_op_bnl_4')
// (9, 21, 'sp4_v_b_28')
// (9, 22, 'sp4_v_b_17')
// (9, 23, 'sp4_v_b_4')
// (10, 16, 'sp4_h_r_25')
// (11, 16, 'sp4_h_r_36')
// (12, 16, 'sp4_h_l_36')

reg n1044 = 0;
// (7, 13, 'sp4_r_v_b_43')
// (7, 14, 'sp4_r_v_b_30')
// (7, 15, 'sp4_r_v_b_19')
// (7, 16, 'sp4_r_v_b_6')
// (7, 17, 'sp4_r_v_b_47')
// (7, 18, 'sp4_r_v_b_34')
// (7, 19, 'neigh_op_tnr_5')
// (7, 19, 'sp4_r_v_b_23')
// (7, 20, 'neigh_op_rgt_5')
// (7, 20, 'sp4_r_v_b_10')
// (7, 21, 'neigh_op_bnr_5')
// (8, 12, 'sp4_v_t_43')
// (8, 13, 'sp4_r_v_b_46')
// (8, 13, 'sp4_v_b_43')
// (8, 14, 'local_g3_6')
// (8, 14, 'lutff_4/in_3')
// (8, 14, 'sp4_r_v_b_35')
// (8, 14, 'sp4_v_b_30')
// (8, 15, 'sp4_r_v_b_22')
// (8, 15, 'sp4_v_b_19')
// (8, 16, 'local_g0_3')
// (8, 16, 'lutff_4/in_1')
// (8, 16, 'sp4_h_r_3')
// (8, 16, 'sp4_r_v_b_11')
// (8, 16, 'sp4_v_b_6')
// (8, 16, 'sp4_v_t_47')
// (8, 17, 'sp4_r_v_b_46')
// (8, 17, 'sp4_v_b_47')
// (8, 18, 'sp4_r_v_b_35')
// (8, 18, 'sp4_v_b_34')
// (8, 19, 'neigh_op_top_5')
// (8, 19, 'sp4_r_v_b_22')
// (8, 19, 'sp4_v_b_23')
// (8, 20, 'local_g2_5')
// (8, 20, 'lutff_5/out')
// (8, 20, 'lutff_6/in_3')
// (8, 20, 'sp4_r_v_b_11')
// (8, 20, 'sp4_v_b_10')
// (8, 21, 'neigh_op_bot_5')
// (9, 12, 'sp4_v_t_46')
// (9, 13, 'local_g2_6')
// (9, 13, 'lutff_1/in_3')
// (9, 13, 'sp4_v_b_46')
// (9, 14, 'sp4_v_b_35')
// (9, 15, 'sp4_v_b_22')
// (9, 16, 'sp4_h_r_14')
// (9, 16, 'sp4_v_b_11')
// (9, 16, 'sp4_v_t_46')
// (9, 17, 'sp4_v_b_46')
// (9, 18, 'sp4_v_b_35')
// (9, 19, 'local_g3_5')
// (9, 19, 'lutff_3/in_1')
// (9, 19, 'neigh_op_tnl_5')
// (9, 19, 'sp4_v_b_22')
// (9, 20, 'local_g1_5')
// (9, 20, 'lutff_1/in_1')
// (9, 20, 'neigh_op_lft_5')
// (9, 20, 'sp4_v_b_11')
// (9, 21, 'neigh_op_bnl_5')
// (10, 16, 'sp4_h_r_27')
// (11, 16, 'sp4_h_r_38')
// (12, 16, 'sp4_h_l_38')

wire n1045;
// (7, 13, 'sp4_r_v_b_45')
// (7, 14, 'sp4_r_v_b_32')
// (7, 15, 'local_g3_4')
// (7, 15, 'lutff_1/in_2')
// (7, 15, 'neigh_op_tnr_4')
// (7, 15, 'sp4_r_v_b_21')
// (7, 16, 'neigh_op_rgt_4')
// (7, 16, 'sp4_r_v_b_40')
// (7, 16, 'sp4_r_v_b_8')
// (7, 17, 'neigh_op_bnr_4')
// (7, 17, 'sp4_r_v_b_29')
// (7, 17, 'sp4_r_v_b_46')
// (7, 18, 'sp4_r_v_b_16')
// (7, 18, 'sp4_r_v_b_35')
// (7, 19, 'sp4_r_v_b_22')
// (7, 19, 'sp4_r_v_b_5')
// (7, 20, 'local_g2_3')
// (7, 20, 'lutff_1/in_2')
// (7, 20, 'sp4_r_v_b_11')
// (8, 12, 'sp4_v_t_45')
// (8, 13, 'sp4_v_b_45')
// (8, 14, 'sp4_v_b_32')
// (8, 15, 'neigh_op_top_4')
// (8, 15, 'sp4_v_b_21')
// (8, 15, 'sp4_v_t_40')
// (8, 16, 'lutff_4/out')
// (8, 16, 'sp4_v_b_40')
// (8, 16, 'sp4_v_b_8')
// (8, 16, 'sp4_v_t_46')
// (8, 17, 'neigh_op_bot_4')
// (8, 17, 'sp4_v_b_29')
// (8, 17, 'sp4_v_b_46')
// (8, 18, 'sp4_v_b_16')
// (8, 18, 'sp4_v_b_35')
// (8, 19, 'local_g1_5')
// (8, 19, 'lutff_1/in_1')
// (8, 19, 'sp4_v_b_22')
// (8, 19, 'sp4_v_b_5')
// (8, 20, 'sp4_v_b_11')
// (9, 15, 'neigh_op_tnl_4')
// (9, 16, 'local_g1_4')
// (9, 16, 'lutff_1/in_2')
// (9, 16, 'neigh_op_lft_4')
// (9, 17, 'neigh_op_bnl_4')

reg n1046 = 0;
// (7, 14, 'local_g0_0')
// (7, 14, 'lutff_2/in_0')
// (7, 14, 'sp4_h_r_0')
// (8, 13, 'neigh_op_tnr_4')
// (8, 14, 'neigh_op_rgt_4')
// (8, 14, 'sp4_h_r_13')
// (8, 15, 'neigh_op_bnr_4')
// (9, 13, 'local_g0_4')
// (9, 13, 'lutff_2/in_2')
// (9, 13, 'neigh_op_top_4')
// (9, 14, 'lutff_4/out')
// (9, 14, 'sp4_h_r_24')
// (9, 15, 'neigh_op_bot_4')
// (10, 13, 'neigh_op_tnl_4')
// (10, 14, 'neigh_op_lft_4')
// (10, 14, 'sp4_h_r_37')
// (10, 15, 'neigh_op_bnl_4')
// (11, 14, 'sp4_h_l_37')

wire n1047;
// (7, 15, 'local_g2_5')
// (7, 15, 'lutff_3/in_2')
// (7, 15, 'neigh_op_tnr_5')
// (7, 16, 'neigh_op_rgt_5')
// (7, 16, 'sp4_r_v_b_42')
// (7, 17, 'neigh_op_bnr_5')
// (7, 17, 'sp4_r_v_b_31')
// (7, 17, 'sp4_r_v_b_41')
// (7, 18, 'sp4_r_v_b_18')
// (7, 18, 'sp4_r_v_b_28')
// (7, 19, 'sp4_r_v_b_17')
// (7, 19, 'sp4_r_v_b_7')
// (7, 20, 'local_g1_4')
// (7, 20, 'lutff_3/in_2')
// (7, 20, 'sp4_r_v_b_4')
// (8, 15, 'neigh_op_top_5')
// (8, 15, 'sp4_v_t_42')
// (8, 16, 'lutff_5/out')
// (8, 16, 'sp4_h_r_10')
// (8, 16, 'sp4_v_b_42')
// (8, 16, 'sp4_v_t_41')
// (8, 17, 'neigh_op_bot_5')
// (8, 17, 'sp4_v_b_31')
// (8, 17, 'sp4_v_b_41')
// (8, 18, 'sp4_v_b_18')
// (8, 18, 'sp4_v_b_28')
// (8, 19, 'local_g0_7')
// (8, 19, 'lutff_3/in_2')
// (8, 19, 'sp4_v_b_17')
// (8, 19, 'sp4_v_b_7')
// (8, 20, 'sp4_v_b_4')
// (9, 15, 'neigh_op_tnl_5')
// (9, 16, 'local_g1_5')
// (9, 16, 'lutff_3/in_1')
// (9, 16, 'neigh_op_lft_5')
// (9, 16, 'sp4_h_r_23')
// (9, 17, 'neigh_op_bnl_5')
// (10, 16, 'sp4_h_r_34')
// (11, 16, 'sp4_h_r_47')
// (12, 16, 'sp4_h_l_47')

wire n1048;
// (7, 15, 'lutff_7/cout')
// (7, 16, 'carry_in')
// (7, 16, 'carry_in_mux')

wire n1049;
// (7, 15, 'neigh_op_tnr_1')
// (7, 16, 'neigh_op_rgt_1')
// (7, 17, 'neigh_op_bnr_1')
// (8, 15, 'neigh_op_top_1')
// (8, 16, 'lutff_1/out')
// (8, 17, 'neigh_op_bot_1')
// (9, 15, 'neigh_op_tnl_1')
// (9, 16, 'neigh_op_lft_1')
// (9, 17, 'local_g3_1')
// (9, 17, 'lutff_3/in_1')
// (9, 17, 'neigh_op_bnl_1')

reg n1050 = 0;
// (7, 15, 'sp4_r_v_b_43')
// (7, 16, 'sp4_r_v_b_30')
// (7, 17, 'sp4_r_v_b_19')
// (7, 18, 'sp4_r_v_b_6')
// (7, 19, 'sp4_r_v_b_38')
// (7, 20, 'neigh_op_tnr_7')
// (7, 20, 'sp4_r_v_b_27')
// (7, 21, 'neigh_op_rgt_7')
// (7, 21, 'sp4_r_v_b_14')
// (7, 22, 'neigh_op_bnr_7')
// (7, 22, 'sp4_r_v_b_3')
// (8, 11, 'sp4_r_v_b_36')
// (8, 12, 'sp4_r_v_b_25')
// (8, 13, 'sp4_r_v_b_12')
// (8, 14, 'local_g0_6')
// (8, 14, 'lutff_5/in_3')
// (8, 14, 'sp4_h_r_6')
// (8, 14, 'sp4_r_v_b_1')
// (8, 14, 'sp4_v_t_43')
// (8, 15, 'sp4_r_v_b_47')
// (8, 15, 'sp4_v_b_43')
// (8, 16, 'local_g3_6')
// (8, 16, 'lutff_7/in_2')
// (8, 16, 'sp4_r_v_b_34')
// (8, 16, 'sp4_v_b_30')
// (8, 17, 'sp4_r_v_b_23')
// (8, 17, 'sp4_v_b_19')
// (8, 18, 'sp4_r_v_b_10')
// (8, 18, 'sp4_v_b_6')
// (8, 18, 'sp4_v_t_38')
// (8, 19, 'sp4_r_v_b_39')
// (8, 19, 'sp4_v_b_38')
// (8, 20, 'neigh_op_top_7')
// (8, 20, 'sp4_r_v_b_26')
// (8, 20, 'sp4_r_v_b_42')
// (8, 20, 'sp4_v_b_27')
// (8, 21, 'lutff_7/out')
// (8, 21, 'sp4_r_v_b_15')
// (8, 21, 'sp4_r_v_b_31')
// (8, 21, 'sp4_v_b_14')
// (8, 22, 'neigh_op_bot_7')
// (8, 22, 'sp4_r_v_b_18')
// (8, 22, 'sp4_r_v_b_2')
// (8, 22, 'sp4_v_b_3')
// (8, 23, 'sp4_r_v_b_7')
// (9, 10, 'sp4_v_t_36')
// (9, 11, 'sp4_v_b_36')
// (9, 12, 'sp4_v_b_25')
// (9, 13, 'local_g1_4')
// (9, 13, 'lutff_3/in_2')
// (9, 13, 'sp4_v_b_12')
// (9, 14, 'sp4_h_r_19')
// (9, 14, 'sp4_v_b_1')
// (9, 14, 'sp4_v_t_47')
// (9, 15, 'sp4_v_b_47')
// (9, 16, 'sp4_v_b_34')
// (9, 17, 'sp4_v_b_23')
// (9, 18, 'sp4_v_b_10')
// (9, 18, 'sp4_v_t_39')
// (9, 19, 'local_g2_7')
// (9, 19, 'lutff_5/in_0')
// (9, 19, 'lutff_7/in_2')
// (9, 19, 'sp4_h_r_7')
// (9, 19, 'sp4_v_b_39')
// (9, 19, 'sp4_v_t_42')
// (9, 20, 'local_g2_7')
// (9, 20, 'lutff_4/in_1')
// (9, 20, 'neigh_op_tnl_7')
// (9, 20, 'sp4_v_b_26')
// (9, 20, 'sp4_v_b_42')
// (9, 21, 'neigh_op_lft_7')
// (9, 21, 'sp4_v_b_15')
// (9, 21, 'sp4_v_b_31')
// (9, 22, 'local_g3_7')
// (9, 22, 'lutff_1/in_1')
// (9, 22, 'neigh_op_bnl_7')
// (9, 22, 'sp4_v_b_18')
// (9, 22, 'sp4_v_b_2')
// (9, 23, 'sp4_v_b_7')
// (10, 14, 'sp4_h_r_30')
// (10, 19, 'local_g1_2')
// (10, 19, 'lutff_7/in_0')
// (10, 19, 'sp4_h_r_18')
// (11, 14, 'sp4_h_r_43')
// (11, 19, 'sp4_h_r_31')
// (12, 14, 'sp4_h_l_43')
// (12, 19, 'sp4_h_r_42')
// (13, 19, 'sp4_h_l_42')

wire n1051;
// (7, 16, 'lutff_0/cout')
// (7, 16, 'lutff_1/in_3')

wire n1052;
// (7, 17, 'neigh_op_tnr_1')
// (7, 18, 'neigh_op_rgt_1')
// (7, 19, 'neigh_op_bnr_1')
// (8, 17, 'neigh_op_top_1')
// (8, 18, 'local_g0_1')
// (8, 18, 'lutff_1/out')
// (8, 18, 'lutff_5/in_2')
// (8, 19, 'neigh_op_bot_1')
// (9, 17, 'neigh_op_tnl_1')
// (9, 18, 'neigh_op_lft_1')
// (9, 19, 'neigh_op_bnl_1')

wire n1053;
// (7, 17, 'neigh_op_tnr_2')
// (7, 18, 'local_g2_2')
// (7, 18, 'lutff_1/in_1')
// (7, 18, 'neigh_op_rgt_2')
// (7, 19, 'neigh_op_bnr_2')
// (8, 15, 'local_g3_0')
// (8, 15, 'lutff_1/in_2')
// (8, 15, 'sp4_r_v_b_40')
// (8, 16, 'sp4_r_v_b_29')
// (8, 17, 'local_g0_2')
// (8, 17, 'lutff_1/in_1')
// (8, 17, 'neigh_op_top_2')
// (8, 17, 'sp4_r_v_b_16')
// (8, 18, 'lutff_2/out')
// (8, 18, 'sp4_r_v_b_5')
// (8, 19, 'neigh_op_bot_2')
// (9, 14, 'sp4_v_t_40')
// (9, 15, 'sp4_v_b_40')
// (9, 16, 'sp4_v_b_29')
// (9, 17, 'neigh_op_tnl_2')
// (9, 17, 'sp4_v_b_16')
// (9, 18, 'local_g1_2')
// (9, 18, 'lutff_1/in_2')
// (9, 18, 'neigh_op_lft_2')
// (9, 18, 'sp4_v_b_5')
// (9, 19, 'neigh_op_bnl_2')

wire n1054;
// (7, 17, 'neigh_op_tnr_3')
// (7, 18, 'neigh_op_rgt_3')
// (7, 19, 'neigh_op_bnr_3')
// (8, 16, 'sp4_r_v_b_47')
// (8, 17, 'neigh_op_top_3')
// (8, 17, 'sp4_r_v_b_34')
// (8, 18, 'lutff_3/out')
// (8, 18, 'sp4_r_v_b_23')
// (8, 19, 'neigh_op_bot_3')
// (8, 19, 'sp4_r_v_b_10')
// (9, 15, 'sp4_v_t_47')
// (9, 16, 'sp4_v_b_47')
// (9, 17, 'neigh_op_tnl_3')
// (9, 17, 'sp4_v_b_34')
// (9, 18, 'neigh_op_lft_3')
// (9, 18, 'sp4_v_b_23')
// (9, 19, 'local_g2_3')
// (9, 19, 'lutff_6/in_3')
// (9, 19, 'neigh_op_bnl_3')
// (9, 19, 'sp4_h_r_10')
// (9, 19, 'sp4_v_b_10')
// (10, 19, 'local_g1_7')
// (10, 19, 'lutff_5/in_1')
// (10, 19, 'sp4_h_r_23')
// (11, 19, 'sp4_h_r_34')
// (12, 19, 'sp4_h_r_47')
// (13, 19, 'sp4_h_l_47')

wire n1055;
// (7, 17, 'neigh_op_tnr_4')
// (7, 18, 'neigh_op_rgt_4')
// (7, 19, 'neigh_op_bnr_4')
// (8, 17, 'neigh_op_top_4')
// (8, 18, 'local_g0_4')
// (8, 18, 'lutff_4/out')
// (8, 18, 'lutff_5/in_1')
// (8, 19, 'neigh_op_bot_4')
// (9, 17, 'neigh_op_tnl_4')
// (9, 18, 'neigh_op_lft_4')
// (9, 19, 'neigh_op_bnl_4')

wire n1056;
// (7, 17, 'neigh_op_tnr_5')
// (7, 18, 'neigh_op_rgt_5')
// (7, 19, 'neigh_op_bnr_5')
// (8, 17, 'neigh_op_top_5')
// (8, 18, 'lutff_5/out')
// (8, 19, 'neigh_op_bot_5')
// (9, 17, 'local_g2_5')
// (9, 17, 'lutff_3/in_0')
// (9, 17, 'neigh_op_tnl_5')
// (9, 18, 'neigh_op_lft_5')
// (9, 19, 'neigh_op_bnl_5')

wire n1057;
// (7, 17, 'neigh_op_tnr_7')
// (7, 18, 'neigh_op_rgt_7')
// (7, 19, 'neigh_op_bnr_7')
// (8, 17, 'neigh_op_top_7')
// (8, 18, 'local_g0_7')
// (8, 18, 'lutff_3/in_0')
// (8, 18, 'lutff_4/in_3')
// (8, 18, 'lutff_7/out')
// (8, 19, 'neigh_op_bot_7')
// (9, 17, 'neigh_op_tnl_7')
// (9, 18, 'neigh_op_lft_7')
// (9, 19, 'neigh_op_bnl_7')

wire n1058;
// (7, 18, 'lutff_7/cout')
// (7, 19, 'carry_in')
// (7, 19, 'carry_in_mux')

wire n1059;
// (7, 19, 'lutff_0/cout')
// (7, 19, 'lutff_1/in_3')

wire n1060;
// (7, 19, 'neigh_op_tnr_1')
// (7, 20, 'neigh_op_rgt_1')
// (7, 21, 'local_g1_1')
// (7, 21, 'lutff_4/in_2')
// (7, 21, 'neigh_op_bnr_1')
// (8, 19, 'neigh_op_top_1')
// (8, 20, 'lutff_1/out')
// (8, 21, 'neigh_op_bot_1')
// (9, 19, 'neigh_op_tnl_1')
// (9, 20, 'neigh_op_lft_1')
// (9, 21, 'neigh_op_bnl_1')

reg n1061 = 0;
// (7, 19, 'neigh_op_tnr_2')
// (7, 20, 'neigh_op_rgt_2')
// (7, 21, 'neigh_op_bnr_2')
// (8, 9, 'sp4_r_v_b_45')
// (8, 10, 'sp4_r_v_b_32')
// (8, 11, 'local_g3_5')
// (8, 11, 'lutff_6/in_2')
// (8, 11, 'sp4_r_v_b_21')
// (8, 12, 'sp4_r_v_b_8')
// (8, 13, 'sp4_r_v_b_45')
// (8, 14, 'local_g2_0')
// (8, 14, 'lutff_0/in_0')
// (8, 14, 'sp4_r_v_b_32')
// (8, 15, 'sp4_r_v_b_21')
// (8, 16, 'local_g2_0')
// (8, 16, 'lutff_6/in_2')
// (8, 16, 'sp4_r_v_b_8')
// (8, 17, 'sp4_r_v_b_40')
// (8, 18, 'sp4_r_v_b_29')
// (8, 19, 'neigh_op_top_2')
// (8, 19, 'sp4_r_v_b_16')
// (8, 20, 'lutff_2/out')
// (8, 20, 'sp4_r_v_b_5')
// (8, 21, 'neigh_op_bot_2')
// (9, 8, 'sp4_v_t_45')
// (9, 9, 'sp4_v_b_45')
// (9, 10, 'sp4_v_b_32')
// (9, 11, 'sp4_v_b_21')
// (9, 12, 'sp4_v_b_8')
// (9, 12, 'sp4_v_t_45')
// (9, 13, 'sp4_v_b_45')
// (9, 14, 'sp4_v_b_32')
// (9, 15, 'sp4_v_b_21')
// (9, 16, 'sp4_v_b_8')
// (9, 16, 'sp4_v_t_40')
// (9, 17, 'sp4_v_b_40')
// (9, 18, 'sp4_v_b_29')
// (9, 19, 'local_g3_2')
// (9, 19, 'lutff_3/in_2')
// (9, 19, 'neigh_op_tnl_2')
// (9, 19, 'sp4_v_b_16')
// (9, 20, 'local_g0_2')
// (9, 20, 'lutff_2/in_2')
// (9, 20, 'neigh_op_lft_2')
// (9, 20, 'sp4_v_b_5')
// (9, 21, 'neigh_op_bnl_2')

wire n1062;
// (7, 19, 'neigh_op_tnr_3')
// (7, 20, 'neigh_op_rgt_3')
// (7, 21, 'neigh_op_bnr_3')
// (8, 19, 'neigh_op_top_3')
// (8, 20, 'local_g3_3')
// (8, 20, 'lutff_3/out')
// (8, 20, 'lutff_global/cen')
// (8, 21, 'neigh_op_bot_3')
// (9, 19, 'neigh_op_tnl_3')
// (9, 20, 'neigh_op_lft_3')
// (9, 21, 'neigh_op_bnl_3')

wire n1063;
// (7, 19, 'neigh_op_tnr_6')
// (7, 20, 'neigh_op_rgt_6')
// (7, 21, 'neigh_op_bnr_6')
// (8, 19, 'neigh_op_top_6')
// (8, 20, 'local_g3_6')
// (8, 20, 'lutff_5/in_2')
// (8, 20, 'lutff_6/out')
// (8, 21, 'neigh_op_bot_6')
// (9, 19, 'neigh_op_tnl_6')
// (9, 20, 'neigh_op_lft_6')
// (9, 21, 'neigh_op_bnl_6')

wire n1064;
// (7, 19, 'neigh_op_tnr_7')
// (7, 20, 'neigh_op_rgt_7')
// (7, 21, 'neigh_op_bnr_7')
// (8, 19, 'neigh_op_top_7')
// (8, 20, 'local_g0_7')
// (8, 20, 'lutff_3/in_0')
// (8, 20, 'lutff_4/in_1')
// (8, 20, 'lutff_6/in_1')
// (8, 20, 'lutff_7/out')
// (8, 21, 'local_g0_7')
// (8, 21, 'lutff_1/in_2')
// (8, 21, 'lutff_3/in_2')
// (8, 21, 'lutff_5/in_0')
// (8, 21, 'lutff_6/in_1')
// (8, 21, 'lutff_7/in_2')
// (8, 21, 'neigh_op_bot_7')
// (9, 19, 'neigh_op_tnl_7')
// (9, 20, 'local_g1_7')
// (9, 20, 'lutff_2/in_0')
// (9, 20, 'neigh_op_lft_7')
// (9, 21, 'local_g2_7')
// (9, 21, 'lutff_1/in_0')
// (9, 21, 'lutff_4/in_3')
// (9, 21, 'neigh_op_bnl_7')

wire n1065;
// (7, 20, 'lutff_7/cout')
// (7, 21, 'carry_in')
// (7, 21, 'carry_in_mux')

wire n1066;
// (7, 20, 'neigh_op_tnr_0')
// (7, 21, 'neigh_op_rgt_0')
// (7, 22, 'neigh_op_bnr_0')
// (8, 20, 'neigh_op_top_0')
// (8, 21, 'local_g0_0')
// (8, 21, 'lutff_0/out')
// (8, 21, 'lutff_7/in_1')
// (8, 22, 'neigh_op_bot_0')
// (9, 20, 'neigh_op_tnl_0')
// (9, 21, 'neigh_op_lft_0')
// (9, 22, 'neigh_op_bnl_0')

wire n1067;
// (7, 20, 'neigh_op_tnr_2')
// (7, 21, 'neigh_op_rgt_2')
// (7, 22, 'neigh_op_bnr_2')
// (8, 20, 'neigh_op_top_2')
// (8, 21, 'local_g2_2')
// (8, 21, 'lutff_2/out')
// (8, 21, 'lutff_5/in_3')
// (8, 22, 'neigh_op_bot_2')
// (9, 20, 'neigh_op_tnl_2')
// (9, 21, 'neigh_op_lft_2')
// (9, 22, 'neigh_op_bnl_2')

wire n1068;
// (7, 20, 'neigh_op_tnr_3')
// (7, 21, 'neigh_op_rgt_3')
// (7, 22, 'neigh_op_bnr_3')
// (8, 20, 'neigh_op_top_3')
// (8, 21, 'local_g3_3')
// (8, 21, 'lutff_3/out')
// (8, 21, 'lutff_global/cen')
// (8, 22, 'neigh_op_bot_3')
// (9, 20, 'neigh_op_tnl_3')
// (9, 21, 'local_g1_3')
// (9, 21, 'lutff_global/cen')
// (9, 21, 'neigh_op_lft_3')
// (9, 22, 'neigh_op_bnl_3')

wire n1069;
// (7, 20, 'neigh_op_tnr_4')
// (7, 21, 'local_g3_4')
// (7, 21, 'lutff_2/in_1')
// (7, 21, 'neigh_op_rgt_4')
// (7, 22, 'neigh_op_bnr_4')
// (8, 20, 'neigh_op_top_4')
// (8, 21, 'local_g3_4')
// (8, 21, 'lutff_0/in_3')
// (8, 21, 'lutff_2/in_1')
// (8, 21, 'lutff_4/out')
// (8, 21, 'sp4_h_r_8')
// (8, 22, 'local_g0_4')
// (8, 22, 'lutff_0/in_2')
// (8, 22, 'lutff_2/in_2')
// (8, 22, 'lutff_3/in_3')
// (8, 22, 'lutff_7/in_3')
// (8, 22, 'neigh_op_bot_4')
// (9, 20, 'neigh_op_tnl_4')
// (9, 21, 'local_g1_4')
// (9, 21, 'lutff_2/in_1')
// (9, 21, 'lutff_3/in_2')
// (9, 21, 'lutff_6/in_3')
// (9, 21, 'neigh_op_lft_4')
// (9, 21, 'sp4_h_r_21')
// (9, 22, 'local_g3_4')
// (9, 22, 'lutff_6/in_3')
// (9, 22, 'lutff_7/in_0')
// (9, 22, 'neigh_op_bnl_4')
// (10, 21, 'local_g3_0')
// (10, 21, 'lutff_7/in_0')
// (10, 21, 'sp4_h_r_32')
// (11, 21, 'local_g2_5')
// (11, 21, 'lutff_3/in_2')
// (11, 21, 'sp4_h_r_45')
// (12, 21, 'sp4_h_l_45')

wire n1070;
// (7, 21, 'lutff_0/cout')
// (7, 21, 'lutff_1/in_3')

wire n1071;
// (7, 21, 'lutff_1/cout')
// (7, 21, 'lutff_2/in_3')

wire n1072;
// (7, 21, 'neigh_op_tnr_0')
// (7, 22, 'neigh_op_rgt_0')
// (7, 23, 'neigh_op_bnr_0')
// (8, 21, 'local_g1_0')
// (8, 21, 'lutff_7/in_0')
// (8, 21, 'neigh_op_top_0')
// (8, 22, 'lutff_0/out')
// (8, 23, 'neigh_op_bot_0')
// (9, 21, 'neigh_op_tnl_0')
// (9, 22, 'neigh_op_lft_0')
// (9, 23, 'neigh_op_bnl_0')

reg n1073 = 0;
// (7, 21, 'neigh_op_tnr_2')
// (7, 22, 'neigh_op_rgt_2')
// (7, 22, 'sp4_h_r_9')
// (7, 23, 'neigh_op_bnr_2')
// (8, 21, 'neigh_op_top_2')
// (8, 22, 'lutff_2/out')
// (8, 22, 'sp4_h_r_20')
// (8, 23, 'neigh_op_bot_2')
// (9, 21, 'neigh_op_tnl_2')
// (9, 22, 'neigh_op_lft_2')
// (9, 22, 'sp4_h_r_33')
// (9, 23, 'neigh_op_bnl_2')
// (10, 19, 'sp4_r_v_b_38')
// (10, 20, 'sp4_r_v_b_27')
// (10, 21, 'local_g2_6')
// (10, 21, 'lutff_7/in_3')
// (10, 21, 'sp4_r_v_b_14')
// (10, 22, 'sp4_h_r_44')
// (10, 22, 'sp4_r_v_b_3')
// (11, 18, 'sp4_v_t_38')
// (11, 19, 'sp4_v_b_38')
// (11, 20, 'sp4_v_b_27')
// (11, 21, 'sp4_v_b_14')
// (11, 22, 'sp4_h_l_44')
// (11, 22, 'sp4_v_b_3')

wire n1074;
// (7, 21, 'neigh_op_tnr_3')
// (7, 22, 'neigh_op_rgt_3')
// (7, 23, 'neigh_op_bnr_3')
// (8, 21, 'local_g1_3')
// (8, 21, 'lutff_5/in_1')
// (8, 21, 'neigh_op_top_3')
// (8, 22, 'lutff_3/out')
// (8, 23, 'neigh_op_bot_3')
// (9, 21, 'neigh_op_tnl_3')
// (9, 22, 'neigh_op_lft_3')
// (9, 23, 'neigh_op_bnl_3')

wire n1075;
// (7, 21, 'neigh_op_tnr_7')
// (7, 22, 'neigh_op_rgt_7')
// (7, 23, 'neigh_op_bnr_7')
// (8, 21, 'local_g1_7')
// (8, 21, 'lutff_1/in_3')
// (8, 21, 'neigh_op_top_7')
// (8, 22, 'lutff_7/out')
// (8, 23, 'neigh_op_bot_7')
// (9, 21, 'neigh_op_tnl_7')
// (9, 22, 'neigh_op_lft_7')
// (9, 23, 'neigh_op_bnl_7')

wire n1076;
// (8, 0, 'logic_op_tnr_0')
// (8, 1, 'neigh_op_rgt_0')
// (8, 2, 'local_g0_0')
// (8, 2, 'lutff_0/in_0')
// (8, 2, 'neigh_op_bnr_0')
// (9, 0, 'logic_op_top_0')
// (9, 1, 'lutff_0/out')
// (9, 2, 'neigh_op_bot_0')
// (10, 0, 'logic_op_tnl_0')
// (10, 1, 'neigh_op_lft_0')
// (10, 2, 'neigh_op_bnl_0')

wire n1077;
// (8, 0, 'logic_op_tnr_1')
// (8, 1, 'neigh_op_rgt_1')
// (8, 2, 'neigh_op_bnr_1')
// (9, 0, 'logic_op_top_1')
// (9, 1, 'lutff_1/out')
// (9, 2, 'neigh_op_bot_1')
// (10, 0, 'logic_op_tnl_1')
// (10, 1, 'neigh_op_lft_1')
// (10, 2, 'local_g2_1')
// (10, 2, 'lutff_1/in_0')
// (10, 2, 'neigh_op_bnl_1')

reg n1078 = 0;
// (8, 0, 'logic_op_tnr_3')
// (8, 1, 'neigh_op_rgt_3')
// (8, 2, 'neigh_op_bnr_3')
// (9, 0, 'logic_op_top_3')
// (9, 1, 'lutff_3/out')
// (9, 1, 'sp4_r_v_b_39')
// (9, 2, 'local_g0_3')
// (9, 2, 'lutff_5/in_0')
// (9, 2, 'neigh_op_bot_3')
// (9, 2, 'sp4_r_v_b_26')
// (9, 3, 'sp4_r_v_b_15')
// (9, 4, 'sp4_r_v_b_2')
// (10, 0, 'logic_op_tnl_3')
// (10, 0, 'span4_vert_39')
// (10, 1, 'neigh_op_lft_3')
// (10, 1, 'sp4_v_b_39')
// (10, 2, 'neigh_op_bnl_3')
// (10, 2, 'sp4_v_b_26')
// (10, 3, 'sp4_v_b_15')
// (10, 4, 'local_g1_2')
// (10, 4, 'lutff_6/in_3')
// (10, 4, 'sp4_v_b_2')

wire n1079;
// (8, 0, 'logic_op_tnr_4')
// (8, 1, 'neigh_op_rgt_4')
// (8, 2, 'local_g1_4')
// (8, 2, 'lutff_3/in_2')
// (8, 2, 'neigh_op_bnr_4')
// (9, 0, 'logic_op_top_4')
// (9, 1, 'lutff_4/out')
// (9, 2, 'neigh_op_bot_4')
// (10, 0, 'logic_op_tnl_4')
// (10, 1, 'neigh_op_lft_4')
// (10, 2, 'neigh_op_bnl_4')

reg n1080 = 0;
// (8, 0, 'logic_op_tnr_5')
// (8, 1, 'neigh_op_rgt_5')
// (8, 1, 'sp4_r_v_b_42')
// (8, 2, 'neigh_op_bnr_5')
// (8, 2, 'sp4_r_v_b_31')
// (8, 3, 'sp4_r_v_b_18')
// (8, 4, 'sp4_r_v_b_7')
// (9, 0, 'logic_op_top_5')
// (9, 0, 'span4_vert_42')
// (9, 1, 'lutff_5/out')
// (9, 1, 'sp4_v_b_42')
// (9, 2, 'local_g2_7')
// (9, 2, 'lutff_0/in_3')
// (9, 2, 'neigh_op_bot_5')
// (9, 2, 'sp4_v_b_31')
// (9, 3, 'sp4_v_b_18')
// (9, 4, 'sp4_v_b_7')
// (10, 0, 'logic_op_tnl_5')
// (10, 1, 'neigh_op_lft_5')
// (10, 2, 'local_g3_5')
// (10, 2, 'lutff_1/in_1')
// (10, 2, 'neigh_op_bnl_5')

wire n1081;
// (8, 0, 'logic_op_tnr_6')
// (8, 1, 'local_g2_6')
// (8, 1, 'lutff_3/in_1')
// (8, 1, 'lutff_7/in_3')
// (8, 1, 'neigh_op_rgt_6')
// (8, 2, 'neigh_op_bnr_6')
// (9, 0, 'logic_op_top_6')
// (9, 1, 'lutff_6/out')
// (9, 2, 'neigh_op_bot_6')
// (10, 0, 'logic_op_tnl_6')
// (10, 1, 'neigh_op_lft_6')
// (10, 2, 'neigh_op_bnl_6')

reg n1082 = 0;
// (8, 0, 'logic_op_tnr_7')
// (8, 1, 'neigh_op_rgt_7')
// (8, 2, 'neigh_op_bnr_7')
// (9, 0, 'logic_op_top_7')
// (9, 1, 'lutff_7/out')
// (9, 1, 'sp4_r_v_b_47')
// (9, 2, 'local_g1_7')
// (9, 2, 'lutff_5/in_1')
// (9, 2, 'neigh_op_bot_7')
// (9, 2, 'sp4_r_v_b_34')
// (9, 3, 'sp4_r_v_b_23')
// (9, 4, 'local_g2_2')
// (9, 4, 'lutff_3/in_1')
// (9, 4, 'sp4_r_v_b_10')
// (10, 0, 'logic_op_tnl_7')
// (10, 0, 'span4_vert_47')
// (10, 1, 'neigh_op_lft_7')
// (10, 1, 'sp4_v_b_47')
// (10, 2, 'neigh_op_bnl_7')
// (10, 2, 'sp4_v_b_34')
// (10, 3, 'sp4_v_b_23')
// (10, 4, 'sp4_v_b_10')

wire n1083;
// (8, 1, 'local_g2_1')
// (8, 1, 'lutff_3/in_0')
// (8, 1, 'lutff_7/in_2')
// (8, 1, 'neigh_op_tnr_1')
// (8, 2, 'neigh_op_rgt_1')
// (8, 3, 'neigh_op_bnr_1')
// (9, 1, 'neigh_op_top_1')
// (9, 2, 'lutff_1/out')
// (9, 3, 'neigh_op_bot_1')
// (10, 1, 'neigh_op_tnl_1')
// (10, 2, 'neigh_op_lft_1')
// (10, 3, 'neigh_op_bnl_1')

wire n1084;
// (8, 1, 'neigh_op_tnr_0')
// (8, 2, 'neigh_op_rgt_0')
// (8, 3, 'local_g1_0')
// (8, 3, 'lutff_7/in_2')
// (8, 3, 'neigh_op_bnr_0')
// (9, 1, 'neigh_op_top_0')
// (9, 2, 'lutff_0/out')
// (9, 3, 'neigh_op_bot_0')
// (10, 1, 'neigh_op_tnl_0')
// (10, 2, 'neigh_op_lft_0')
// (10, 3, 'neigh_op_bnl_0')

wire n1085;
// (8, 1, 'neigh_op_tnr_2')
// (8, 2, 'local_g2_2')
// (8, 2, 'lutff_0/in_2')
// (8, 2, 'neigh_op_rgt_2')
// (8, 3, 'neigh_op_bnr_2')
// (9, 1, 'neigh_op_top_2')
// (9, 2, 'lutff_2/out')
// (9, 3, 'local_g0_2')
// (9, 3, 'lutff_6/in_0')
// (9, 3, 'neigh_op_bot_2')
// (10, 1, 'neigh_op_tnl_2')
// (10, 2, 'neigh_op_lft_2')
// (10, 3, 'neigh_op_bnl_2')

wire n1086;
// (8, 1, 'neigh_op_tnr_3')
// (8, 2, 'neigh_op_rgt_3')
// (8, 3, 'local_g0_3')
// (8, 3, 'lutff_0/in_3')
// (8, 3, 'neigh_op_bnr_3')
// (9, 1, 'neigh_op_top_3')
// (9, 2, 'lutff_3/out')
// (9, 3, 'neigh_op_bot_3')
// (10, 1, 'neigh_op_tnl_3')
// (10, 2, 'neigh_op_lft_3')
// (10, 3, 'neigh_op_bnl_3')

wire n1087;
// (8, 1, 'neigh_op_tnr_4')
// (8, 2, 'neigh_op_rgt_4')
// (8, 2, 'sp4_r_v_b_40')
// (8, 3, 'neigh_op_bnr_4')
// (8, 3, 'sp4_r_v_b_29')
// (8, 4, 'local_g3_0')
// (8, 4, 'lutff_5/in_0')
// (8, 4, 'sp4_r_v_b_16')
// (8, 5, 'sp4_r_v_b_5')
// (9, 1, 'neigh_op_top_4')
// (9, 1, 'sp4_v_t_40')
// (9, 2, 'lutff_4/out')
// (9, 2, 'sp4_v_b_40')
// (9, 3, 'neigh_op_bot_4')
// (9, 3, 'sp4_v_b_29')
// (9, 4, 'sp4_v_b_16')
// (9, 5, 'sp4_v_b_5')
// (10, 1, 'neigh_op_tnl_4')
// (10, 2, 'neigh_op_lft_4')
// (10, 3, 'neigh_op_bnl_4')

wire n1088;
// (8, 1, 'neigh_op_tnr_5')
// (8, 2, 'neigh_op_rgt_5')
// (8, 3, 'neigh_op_bnr_5')
// (9, 1, 'neigh_op_top_5')
// (9, 2, 'local_g3_5')
// (9, 2, 'lutff_5/out')
// (9, 2, 'lutff_7/in_1')
// (9, 3, 'neigh_op_bot_5')
// (10, 1, 'neigh_op_tnl_5')
// (10, 2, 'neigh_op_lft_5')
// (10, 3, 'neigh_op_bnl_5')

wire n1089;
// (8, 1, 'neigh_op_tnr_6')
// (8, 2, 'neigh_op_rgt_6')
// (8, 3, 'local_g0_6')
// (8, 3, 'lutff_0/in_2')
// (8, 3, 'neigh_op_bnr_6')
// (9, 1, 'neigh_op_top_6')
// (9, 2, 'lutff_6/out')
// (9, 3, 'neigh_op_bot_6')
// (10, 1, 'neigh_op_tnl_6')
// (10, 2, 'neigh_op_lft_6')
// (10, 3, 'neigh_op_bnl_6')

wire n1090;
// (8, 1, 'neigh_op_tnr_7')
// (8, 2, 'neigh_op_rgt_7')
// (8, 3, 'neigh_op_bnr_7')
// (9, 1, 'local_g1_7')
// (9, 1, 'lutff_0/in_2')
// (9, 1, 'neigh_op_top_7')
// (9, 2, 'lutff_7/out')
// (9, 3, 'local_g1_7')
// (9, 3, 'lutff_3/in_3')
// (9, 3, 'neigh_op_bot_7')
// (10, 1, 'neigh_op_tnl_7')
// (10, 2, 'neigh_op_lft_7')
// (10, 3, 'neigh_op_bnl_7')

reg n1091 = 0;
// (8, 1, 'sp4_r_v_b_24')
// (8, 2, 'neigh_op_tnr_0')
// (8, 2, 'sp4_r_v_b_13')
// (8, 3, 'neigh_op_rgt_0')
// (8, 3, 'sp4_r_v_b_0')
// (8, 4, 'neigh_op_bnr_0')
// (9, 0, 'span4_vert_24')
// (9, 1, 'local_g2_0')
// (9, 1, 'lutff_1/in_3')
// (9, 1, 'sp4_v_b_24')
// (9, 2, 'neigh_op_top_0')
// (9, 2, 'sp4_v_b_13')
// (9, 3, 'lutff_0/out')
// (9, 3, 'sp4_v_b_0')
// (9, 4, 'neigh_op_bot_0')
// (10, 2, 'neigh_op_tnl_0')
// (10, 3, 'local_g1_0')
// (10, 3, 'lutff_3/in_2')
// (10, 3, 'neigh_op_lft_0')
// (10, 4, 'neigh_op_bnl_0')

wire n1092;
// (8, 2, 'local_g2_1')
// (8, 2, 'lutff_0/in_1')
// (8, 2, 'neigh_op_tnr_1')
// (8, 3, 'neigh_op_rgt_1')
// (8, 4, 'neigh_op_bnr_1')
// (9, 2, 'neigh_op_top_1')
// (9, 3, 'local_g2_1')
// (9, 3, 'lutff_1/out')
// (9, 3, 'lutff_6/in_3')
// (9, 4, 'neigh_op_bot_1')
// (10, 2, 'neigh_op_tnl_1')
// (10, 3, 'neigh_op_lft_1')
// (10, 4, 'neigh_op_bnl_1')

wire n1093;
// (8, 2, 'local_g2_3')
// (8, 2, 'lutff_6/in_1')
// (8, 2, 'neigh_op_tnr_3')
// (8, 3, 'neigh_op_rgt_3')
// (8, 4, 'neigh_op_bnr_3')
// (9, 2, 'neigh_op_top_3')
// (9, 3, 'lutff_3/out')
// (9, 4, 'neigh_op_bot_3')
// (10, 2, 'neigh_op_tnl_3')
// (10, 3, 'neigh_op_lft_3')
// (10, 4, 'neigh_op_bnl_3')

wire n1094;
// (8, 2, 'local_g2_6')
// (8, 2, 'lutff_6/in_2')
// (8, 2, 'neigh_op_tnr_6')
// (8, 3, 'neigh_op_rgt_6')
// (8, 4, 'neigh_op_bnr_6')
// (9, 2, 'neigh_op_top_6')
// (9, 3, 'lutff_6/out')
// (9, 4, 'neigh_op_bot_6')
// (10, 2, 'neigh_op_tnl_6')
// (10, 3, 'neigh_op_lft_6')
// (10, 4, 'neigh_op_bnl_6')

reg n1095 = 0;
// (8, 2, 'neigh_op_tnr_2')
// (8, 3, 'neigh_op_rgt_2')
// (8, 4, 'neigh_op_bnr_2')
// (9, 2, 'neigh_op_top_2')
// (9, 3, 'local_g3_2')
// (9, 3, 'lutff_2/out')
// (9, 3, 'lutff_5/in_2')
// (9, 3, 'lutff_7/in_2')
// (9, 4, 'neigh_op_bot_2')
// (10, 2, 'neigh_op_tnl_2')
// (10, 3, 'neigh_op_lft_2')
// (10, 4, 'neigh_op_bnl_2')

wire n1096;
// (8, 2, 'neigh_op_tnr_5')
// (8, 3, 'neigh_op_rgt_5')
// (8, 4, 'neigh_op_bnr_5')
// (9, 2, 'local_g0_5')
// (9, 2, 'lutff_7/in_0')
// (9, 2, 'neigh_op_top_5')
// (9, 3, 'lutff_5/out')
// (9, 4, 'neigh_op_bot_5')
// (10, 2, 'neigh_op_tnl_5')
// (10, 3, 'neigh_op_lft_5')
// (10, 4, 'neigh_op_bnl_5')

wire n1097;
// (8, 2, 'neigh_op_tnr_7')
// (8, 3, 'neigh_op_rgt_7')
// (8, 4, 'neigh_op_bnr_7')
// (9, 2, 'neigh_op_top_7')
// (9, 3, 'lutff_7/out')
// (9, 4, 'local_g1_7')
// (9, 4, 'lutff_2/in_0')
// (9, 4, 'neigh_op_bot_7')
// (10, 2, 'neigh_op_tnl_7')
// (10, 3, 'neigh_op_lft_7')
// (10, 4, 'neigh_op_bnl_7')

wire n1098;
// (8, 2, 'sp4_h_r_4')
// (9, 1, 'neigh_op_tnr_6')
// (9, 2, 'local_g0_1')
// (9, 2, 'lutff_2/in_1')
// (9, 2, 'neigh_op_rgt_6')
// (9, 2, 'sp4_h_r_17')
// (9, 3, 'neigh_op_bnr_6')
// (10, 1, 'neigh_op_top_6')
// (10, 2, 'lutff_6/out')
// (10, 2, 'sp4_h_r_28')
// (10, 3, 'neigh_op_bot_6')
// (11, 1, 'neigh_op_tnl_6')
// (11, 2, 'neigh_op_lft_6')
// (11, 2, 'sp4_h_r_41')
// (11, 3, 'neigh_op_bnl_6')
// (12, 2, 'sp4_h_l_41')

wire n1099;
// (8, 3, 'local_g2_5')
// (8, 3, 'lutff_1/in_2')
// (8, 3, 'neigh_op_tnr_5')
// (8, 4, 'neigh_op_rgt_5')
// (8, 5, 'neigh_op_bnr_5')
// (9, 3, 'neigh_op_top_5')
// (9, 4, 'lutff_5/out')
// (9, 5, 'neigh_op_bot_5')
// (10, 3, 'neigh_op_tnl_5')
// (10, 4, 'neigh_op_lft_5')
// (10, 5, 'neigh_op_bnl_5')

wire n1100;
// (8, 3, 'local_g2_7')
// (8, 3, 'lutff_1/in_0')
// (8, 3, 'neigh_op_tnr_7')
// (8, 4, 'neigh_op_rgt_7')
// (8, 5, 'neigh_op_bnr_7')
// (9, 3, 'neigh_op_top_7')
// (9, 4, 'lutff_7/out')
// (9, 5, 'neigh_op_bot_7')
// (10, 3, 'neigh_op_tnl_7')
// (10, 4, 'neigh_op_lft_7')
// (10, 5, 'neigh_op_bnl_7')

wire n1101;
// (8, 3, 'neigh_op_tnr_1')
// (8, 4, 'local_g2_1')
// (8, 4, 'lutff_2/in_1')
// (8, 4, 'neigh_op_rgt_1')
// (8, 5, 'neigh_op_bnr_1')
// (9, 3, 'neigh_op_top_1')
// (9, 4, 'lutff_1/out')
// (9, 5, 'neigh_op_bot_1')
// (10, 3, 'neigh_op_tnl_1')
// (10, 4, 'neigh_op_lft_1')
// (10, 5, 'neigh_op_bnl_1')

wire n1102;
// (8, 3, 'neigh_op_tnr_2')
// (8, 4, 'local_g3_2')
// (8, 4, 'lutff_6/in_1')
// (8, 4, 'neigh_op_rgt_2')
// (8, 5, 'neigh_op_bnr_2')
// (9, 3, 'neigh_op_top_2')
// (9, 4, 'lutff_2/out')
// (9, 5, 'neigh_op_bot_2')
// (10, 3, 'neigh_op_tnl_2')
// (10, 4, 'neigh_op_lft_2')
// (10, 5, 'neigh_op_bnl_2')

wire n1103;
// (8, 3, 'neigh_op_tnr_3')
// (8, 4, 'neigh_op_rgt_3')
// (8, 5, 'neigh_op_bnr_3')
// (9, 3, 'neigh_op_top_3')
// (9, 4, 'local_g2_3')
// (9, 4, 'lutff_1/in_2')
// (9, 4, 'lutff_3/out')
// (9, 5, 'neigh_op_bot_3')
// (10, 3, 'neigh_op_tnl_3')
// (10, 4, 'neigh_op_lft_3')
// (10, 5, 'neigh_op_bnl_3')

reg n1104 = 0;
// (8, 3, 'neigh_op_tnr_4')
// (8, 4, 'neigh_op_rgt_4')
// (8, 5, 'neigh_op_bnr_4')
// (9, 3, 'neigh_op_top_4')
// (9, 4, 'local_g2_4')
// (9, 4, 'local_g3_4')
// (9, 4, 'lutff_1/in_3')
// (9, 4, 'lutff_4/out')
// (9, 4, 'lutff_5/in_0')
// (9, 5, 'neigh_op_bot_4')
// (10, 3, 'neigh_op_tnl_4')
// (10, 4, 'neigh_op_lft_4')
// (10, 5, 'neigh_op_bnl_4')

reg n1105 = 0;
// (8, 3, 'neigh_op_tnr_6')
// (8, 4, 'neigh_op_rgt_6')
// (8, 5, 'neigh_op_bnr_6')
// (9, 3, 'neigh_op_top_6')
// (9, 4, 'local_g2_6')
// (9, 4, 'local_g3_6')
// (9, 4, 'lutff_2/in_1')
// (9, 4, 'lutff_5/in_1')
// (9, 4, 'lutff_6/out')
// (9, 5, 'neigh_op_bot_6')
// (10, 3, 'neigh_op_tnl_6')
// (10, 4, 'neigh_op_lft_6')
// (10, 5, 'neigh_op_bnl_6')

wire n1106;
// (8, 3, 'sp4_r_v_b_47')
// (8, 4, 'sp4_r_v_b_34')
// (8, 5, 'local_g3_7')
// (8, 5, 'lutff_2/in_0')
// (8, 5, 'sp4_r_v_b_23')
// (8, 6, 'local_g2_2')
// (8, 6, 'lutff_1/in_3')
// (8, 6, 'lutff_2/in_0')
// (8, 6, 'lutff_5/in_1')
// (8, 6, 'lutff_7/in_1')
// (8, 6, 'sp4_r_v_b_10')
// (9, 2, 'sp4_v_t_47')
// (9, 3, 'sp4_v_b_47')
// (9, 4, 'sp4_v_b_34')
// (9, 5, 'sp4_v_b_23')
// (9, 6, 'sp4_h_r_10')
// (9, 6, 'sp4_v_b_10')
// (10, 3, 'sp4_r_v_b_39')
// (10, 4, 'sp4_r_v_b_26')
// (10, 4, 'sp4_r_v_b_42')
// (10, 5, 'neigh_op_tnr_1')
// (10, 5, 'sp4_r_v_b_15')
// (10, 5, 'sp4_r_v_b_31')
// (10, 6, 'neigh_op_rgt_1')
// (10, 6, 'sp4_h_r_23')
// (10, 6, 'sp4_r_v_b_18')
// (10, 6, 'sp4_r_v_b_2')
// (10, 7, 'neigh_op_bnr_1')
// (10, 7, 'sp4_r_v_b_7')
// (11, 2, 'sp4_v_t_39')
// (11, 3, 'sp4_h_r_7')
// (11, 3, 'sp4_v_b_39')
// (11, 3, 'sp4_v_t_42')
// (11, 4, 'local_g3_2')
// (11, 4, 'lutff_0/in_1')
// (11, 4, 'sp4_v_b_26')
// (11, 4, 'sp4_v_b_42')
// (11, 5, 'local_g1_1')
// (11, 5, 'lutff_0/in_2')
// (11, 5, 'lutff_4/in_0')
// (11, 5, 'neigh_op_top_1')
// (11, 5, 'sp4_v_b_15')
// (11, 5, 'sp4_v_b_31')
// (11, 6, 'lutff_1/out')
// (11, 6, 'sp4_h_r_34')
// (11, 6, 'sp4_v_b_18')
// (11, 6, 'sp4_v_b_2')
// (11, 7, 'neigh_op_bot_1')
// (11, 7, 'sp4_v_b_7')
// (12, 3, 'sp4_h_r_18')
// (12, 5, 'neigh_op_tnl_1')
// (12, 6, 'neigh_op_lft_1')
// (12, 6, 'sp4_h_r_47')
// (12, 7, 'neigh_op_bnl_1')
// (13, 3, 'local_g2_7')
// (13, 3, 'lutff_5/in_0')
// (13, 3, 'sp4_h_r_31')
// (13, 6, 'sp4_h_l_47')
// (14, 3, 'sp4_h_r_42')
// (15, 3, 'sp4_h_l_42')

wire n1107;
// (8, 4, 'local_g1_2')
// (8, 4, 'lutff_5/in_2')
// (8, 4, 'sp4_h_r_10')
// (9, 2, 'local_g3_2')
// (9, 2, 'lutff_0/in_1')
// (9, 2, 'sp4_r_v_b_42')
// (9, 3, 'local_g3_1')
// (9, 3, 'lutff_7/in_3')
// (9, 3, 'neigh_op_tnr_1')
// (9, 3, 'sp4_r_v_b_31')
// (9, 4, 'local_g3_1')
// (9, 4, 'lutff_3/in_3')
// (9, 4, 'neigh_op_rgt_1')
// (9, 4, 'sp4_h_r_23')
// (9, 4, 'sp4_r_v_b_18')
// (9, 5, 'neigh_op_bnr_1')
// (9, 5, 'sp4_r_v_b_7')
// (10, 1, 'sp4_v_t_42')
// (10, 2, 'sp4_v_b_42')
// (10, 3, 'local_g1_1')
// (10, 3, 'lutff_3/in_1')
// (10, 3, 'neigh_op_top_1')
// (10, 3, 'sp4_v_b_31')
// (10, 4, 'local_g2_1')
// (10, 4, 'local_g3_1')
// (10, 4, 'lutff_1/out')
// (10, 4, 'lutff_5/in_0')
// (10, 4, 'lutff_6/in_0')
// (10, 4, 'sp4_h_r_34')
// (10, 4, 'sp4_v_b_18')
// (10, 5, 'neigh_op_bot_1')
// (10, 5, 'sp4_v_b_7')
// (11, 3, 'neigh_op_tnl_1')
// (11, 4, 'neigh_op_lft_1')
// (11, 4, 'sp4_h_r_47')
// (11, 5, 'neigh_op_bnl_1')
// (12, 4, 'sp4_h_l_47')

wire n1108;
// (8, 4, 'neigh_op_tnr_0')
// (8, 5, 'local_g2_0')
// (8, 5, 'lutff_4/in_2')
// (8, 5, 'neigh_op_rgt_0')
// (8, 6, 'neigh_op_bnr_0')
// (9, 4, 'neigh_op_top_0')
// (9, 5, 'lutff_0/out')
// (9, 6, 'neigh_op_bot_0')
// (10, 4, 'neigh_op_tnl_0')
// (10, 5, 'neigh_op_lft_0')
// (10, 6, 'neigh_op_bnl_0')

wire n1109;
// (8, 4, 'neigh_op_tnr_2')
// (8, 5, 'local_g2_2')
// (8, 5, 'lutff_6/in_2')
// (8, 5, 'neigh_op_rgt_2')
// (8, 6, 'neigh_op_bnr_2')
// (9, 4, 'neigh_op_top_2')
// (9, 5, 'lutff_2/out')
// (9, 6, 'neigh_op_bot_2')
// (10, 4, 'neigh_op_tnl_2')
// (10, 5, 'neigh_op_lft_2')
// (10, 6, 'neigh_op_bnl_2')

reg n1110 = 0;
// (8, 4, 'neigh_op_tnr_3')
// (8, 5, 'neigh_op_rgt_3')
// (8, 6, 'neigh_op_bnr_3')
// (9, 4, 'local_g1_3')
// (9, 4, 'lutff_7/in_3')
// (9, 4, 'neigh_op_top_3')
// (9, 5, 'local_g0_3')
// (9, 5, 'lutff_2/in_3')
// (9, 5, 'lutff_3/out')
// (9, 6, 'neigh_op_bot_3')
// (10, 4, 'neigh_op_tnl_3')
// (10, 5, 'neigh_op_lft_3')
// (10, 6, 'neigh_op_bnl_3')

wire n1111;
// (8, 4, 'neigh_op_tnr_4')
// (8, 5, 'neigh_op_rgt_4')
// (8, 6, 'neigh_op_bnr_4')
// (9, 4, 'neigh_op_top_4')
// (9, 5, 'local_g1_4')
// (9, 5, 'lutff_4/out')
// (9, 5, 'lutff_7/in_0')
// (9, 6, 'neigh_op_bot_4')
// (10, 4, 'neigh_op_tnl_4')
// (10, 5, 'neigh_op_lft_4')
// (10, 6, 'neigh_op_bnl_4')

wire n1112;
// (8, 4, 'neigh_op_tnr_5')
// (8, 5, 'neigh_op_rgt_5')
// (8, 6, 'neigh_op_bnr_5')
// (9, 4, 'local_g0_5')
// (9, 4, 'lutff_1/in_0')
// (9, 4, 'lutff_2/in_3')
// (9, 4, 'neigh_op_top_5')
// (9, 5, 'local_g3_5')
// (9, 5, 'lutff_2/in_2')
// (9, 5, 'lutff_5/out')
// (9, 6, 'neigh_op_bot_5')
// (10, 4, 'neigh_op_tnl_5')
// (10, 5, 'neigh_op_lft_5')
// (10, 6, 'neigh_op_bnl_5')

reg n1113 = 0;
// (8, 4, 'neigh_op_tnr_6')
// (8, 5, 'neigh_op_rgt_6')
// (8, 6, 'neigh_op_bnr_6')
// (9, 4, 'local_g0_6')
// (9, 4, 'lutff_7/in_1')
// (9, 4, 'neigh_op_top_6')
// (9, 5, 'local_g2_6')
// (9, 5, 'lutff_6/out')
// (9, 5, 'lutff_7/in_1')
// (9, 6, 'neigh_op_bot_6')
// (10, 4, 'neigh_op_tnl_6')
// (10, 5, 'neigh_op_lft_6')
// (10, 6, 'neigh_op_bnl_6')

wire n1114;
// (8, 4, 'neigh_op_tnr_7')
// (8, 5, 'neigh_op_rgt_7')
// (8, 6, 'neigh_op_bnr_7')
// (9, 4, 'neigh_op_top_7')
// (9, 5, 'local_g0_7')
// (9, 5, 'lutff_0/in_3')
// (9, 5, 'lutff_7/out')
// (9, 6, 'neigh_op_bot_7')
// (10, 4, 'neigh_op_tnl_7')
// (10, 5, 'neigh_op_lft_7')
// (10, 6, 'neigh_op_bnl_7')

wire n1115;
// (8, 5, 'local_g1_3')
// (8, 5, 'lutff_3/in_1')
// (8, 5, 'sp4_h_r_3')
// (9, 5, 'sp4_h_r_14')
// (10, 5, 'sp4_h_r_27')
// (10, 5, 'sp4_r_v_b_40')
// (10, 6, 'local_g1_5')
// (10, 6, 'lutff_2/in_2')
// (10, 6, 'sp4_r_v_b_29')
// (10, 7, 'sp4_r_v_b_16')
// (10, 8, 'sp4_r_v_b_5')
// (11, 4, 'sp4_v_t_40')
// (11, 5, 'sp4_h_r_38')
// (11, 5, 'sp4_v_b_40')
// (11, 6, 'local_g2_4')
// (11, 6, 'lutff_0/in_0')
// (11, 6, 'sp4_r_v_b_36')
// (11, 6, 'sp4_v_b_29')
// (11, 7, 'sp4_r_v_b_25')
// (11, 7, 'sp4_v_b_16')
// (11, 8, 'sp4_h_r_0')
// (11, 8, 'sp4_r_v_b_12')
// (11, 8, 'sp4_v_b_5')
// (11, 9, 'sp4_r_v_b_1')
// (12, 5, 'sp4_h_l_38')
// (12, 5, 'sp4_h_r_7')
// (12, 5, 'sp4_v_t_36')
// (12, 6, 'sp4_v_b_36')
// (12, 7, 'sp4_v_b_25')
// (12, 8, 'sp4_h_r_13')
// (12, 8, 'sp4_v_b_12')
// (12, 9, 'sp4_v_b_1')
// (13, 5, 'sp4_h_r_18')
// (13, 8, 'sp4_h_r_24')
// (14, 4, 'local_g2_5')
// (14, 4, 'lutff_0/in_3')
// (14, 4, 'neigh_op_tnr_5')
// (14, 5, 'neigh_op_rgt_5')
// (14, 5, 'sp4_h_r_31')
// (14, 5, 'sp4_r_v_b_42')
// (14, 6, 'neigh_op_bnr_5')
// (14, 6, 'sp4_r_v_b_31')
// (14, 7, 'sp4_r_v_b_18')
// (14, 8, 'sp4_h_r_37')
// (14, 8, 'sp4_r_v_b_7')
// (15, 4, 'neigh_op_top_5')
// (15, 4, 'sp4_v_t_42')
// (15, 5, 'lutff_5/out')
// (15, 5, 'sp4_h_r_42')
// (15, 5, 'sp4_v_b_42')
// (15, 6, 'neigh_op_bot_5')
// (15, 6, 'sp4_v_b_31')
// (15, 7, 'sp4_v_b_18')
// (15, 8, 'sp4_h_l_37')
// (15, 8, 'sp4_v_b_7')
// (16, 4, 'neigh_op_tnl_5')
// (16, 5, 'neigh_op_lft_5')
// (16, 5, 'sp4_h_l_42')
// (16, 6, 'neigh_op_bnl_5')

wire n1116;
// (8, 5, 'local_g2_5')
// (8, 5, 'lutff_3/in_0')
// (8, 5, 'neigh_op_tnr_5')
// (8, 6, 'neigh_op_rgt_5')
// (8, 7, 'neigh_op_bnr_5')
// (9, 5, 'neigh_op_top_5')
// (9, 6, 'local_g3_5')
// (9, 6, 'lutff_4/in_0')
// (9, 6, 'lutff_5/out')
// (9, 7, 'local_g1_5')
// (9, 7, 'lutff_7/in_1')
// (9, 7, 'neigh_op_bot_5')
// (10, 5, 'neigh_op_tnl_5')
// (10, 6, 'neigh_op_lft_5')
// (10, 7, 'neigh_op_bnl_5')

reg n1117 = 0;
// (8, 5, 'neigh_op_tnr_1')
// (8, 6, 'neigh_op_rgt_1')
// (8, 7, 'neigh_op_bnr_1')
// (9, 5, 'neigh_op_top_1')
// (9, 6, 'local_g3_1')
// (9, 6, 'lutff_1/out')
// (9, 6, 'lutff_3/in_1')
// (9, 7, 'neigh_op_bot_1')
// (10, 5, 'neigh_op_tnl_1')
// (10, 6, 'neigh_op_lft_1')
// (10, 7, 'neigh_op_bnl_1')

wire n1118;
// (8, 5, 'neigh_op_tnr_3')
// (8, 6, 'neigh_op_rgt_3')
// (8, 7, 'neigh_op_bnr_3')
// (9, 5, 'neigh_op_top_3')
// (9, 6, 'lutff_3/out')
// (9, 6, 'sp4_r_v_b_39')
// (9, 7, 'neigh_op_bot_3')
// (9, 7, 'sp4_r_v_b_26')
// (9, 8, 'sp4_r_v_b_15')
// (9, 9, 'sp4_r_v_b_2')
// (10, 5, 'neigh_op_tnl_3')
// (10, 5, 'sp4_v_t_39')
// (10, 6, 'neigh_op_lft_3')
// (10, 6, 'sp4_v_b_39')
// (10, 7, 'neigh_op_bnl_3')
// (10, 7, 'sp4_v_b_26')
// (10, 8, 'local_g1_7')
// (10, 8, 'lutff_0/in_0')
// (10, 8, 'sp4_v_b_15')
// (10, 9, 'sp4_v_b_2')

reg n1119 = 0;
// (8, 5, 'neigh_op_tnr_6')
// (8, 6, 'neigh_op_rgt_6')
// (8, 7, 'neigh_op_bnr_6')
// (9, 0, 'span12_vert_23')
// (9, 1, 'sp12_v_b_23')
// (9, 2, 'sp12_v_b_20')
// (9, 3, 'sp12_v_b_19')
// (9, 4, 'sp12_v_b_16')
// (9, 5, 'neigh_op_top_6')
// (9, 5, 'sp12_v_b_15')
// (9, 6, 'lutff_6/out')
// (9, 6, 'sp12_v_b_12')
// (9, 7, 'neigh_op_bot_6')
// (9, 7, 'sp12_v_b_11')
// (9, 8, 'sp12_v_b_8')
// (9, 9, 'sp12_v_b_7')
// (9, 10, 'local_g3_4')
// (9, 10, 'lutff_7/in_0')
// (9, 10, 'sp12_v_b_4')
// (9, 11, 'sp12_v_b_3')
// (9, 12, 'sp12_v_b_0')
// (10, 5, 'neigh_op_tnl_6')
// (10, 6, 'neigh_op_lft_6')
// (10, 7, 'neigh_op_bnl_6')

wire n1120;
// (8, 5, 'sp4_h_r_5')
// (9, 5, 'sp4_h_r_16')
// (10, 1, 'local_g1_3')
// (10, 1, 'lutff_global/cen')
// (10, 1, 'sp4_r_v_b_27')
// (10, 2, 'sp4_r_v_b_14')
// (10, 3, 'sp4_r_v_b_3')
// (10, 4, 'neigh_op_tnr_4')
// (10, 4, 'sp4_r_v_b_37')
// (10, 5, 'neigh_op_rgt_4')
// (10, 5, 'sp4_h_r_29')
// (10, 5, 'sp4_r_v_b_24')
// (10, 6, 'neigh_op_bnr_4')
// (10, 6, 'sp4_r_v_b_13')
// (10, 7, 'sp4_r_v_b_0')
// (11, 0, 'span4_vert_27')
// (11, 1, 'sp4_v_b_27')
// (11, 2, 'local_g3_3')
// (11, 2, 'lutff_global/cen')
// (11, 2, 'sp4_r_v_b_43')
// (11, 2, 'sp4_v_b_14')
// (11, 3, 'sp4_r_v_b_30')
// (11, 3, 'sp4_v_b_3')
// (11, 3, 'sp4_v_t_37')
// (11, 4, 'neigh_op_top_4')
// (11, 4, 'sp4_r_v_b_19')
// (11, 4, 'sp4_v_b_37')
// (11, 5, 'lutff_4/out')
// (11, 5, 'sp4_h_r_40')
// (11, 5, 'sp4_r_v_b_6')
// (11, 5, 'sp4_v_b_24')
// (11, 6, 'neigh_op_bot_4')
// (11, 6, 'sp4_v_b_13')
// (11, 7, 'sp4_v_b_0')
// (12, 1, 'sp4_v_t_43')
// (12, 2, 'sp4_v_b_43')
// (12, 3, 'sp4_v_b_30')
// (12, 4, 'neigh_op_tnl_4')
// (12, 4, 'sp4_v_b_19')
// (12, 5, 'neigh_op_lft_4')
// (12, 5, 'sp4_h_l_40')
// (12, 5, 'sp4_h_r_1')
// (12, 5, 'sp4_v_b_6')
// (12, 6, 'neigh_op_bnl_4')
// (13, 5, 'sp4_h_r_12')
// (14, 5, 'sp4_h_r_25')
// (15, 5, 'sp4_h_r_36')
// (16, 5, 'sp4_h_l_36')

reg n1121 = 0;
// (8, 5, 'sp4_r_v_b_39')
// (8, 6, 'sp4_r_v_b_26')
// (8, 7, 'neigh_op_tnr_1')
// (8, 7, 'sp4_r_v_b_15')
// (8, 8, 'neigh_op_rgt_1')
// (8, 8, 'sp4_r_v_b_2')
// (8, 9, 'neigh_op_bnr_1')
// (9, 4, 'sp4_v_t_39')
// (9, 5, 'sp4_v_b_39')
// (9, 6, 'local_g2_2')
// (9, 6, 'lutff_3/in_3')
// (9, 6, 'sp4_v_b_26')
// (9, 7, 'neigh_op_top_1')
// (9, 7, 'sp4_v_b_15')
// (9, 8, 'lutff_1/out')
// (9, 8, 'sp4_v_b_2')
// (9, 9, 'neigh_op_bot_1')
// (10, 7, 'neigh_op_tnl_1')
// (10, 8, 'neigh_op_lft_1')
// (10, 9, 'neigh_op_bnl_1')

wire n1122;
// (8, 6, 'local_g0_5')
// (8, 6, 'lutff_2/in_3')
// (8, 6, 'lutff_3/in_2')
// (8, 6, 'lutff_5/in_2')
// (8, 6, 'sp4_h_r_5')
// (9, 6, 'sp4_h_r_16')
// (10, 5, 'neigh_op_tnr_4')
// (10, 6, 'neigh_op_rgt_4')
// (10, 6, 'sp4_h_r_29')
// (10, 7, 'neigh_op_bnr_4')
// (11, 5, 'neigh_op_top_4')
// (11, 6, 'local_g0_4')
// (11, 6, 'lutff_0/in_2')
// (11, 6, 'lutff_4/out')
// (11, 6, 'sp4_h_r_40')
// (11, 7, 'local_g0_4')
// (11, 7, 'lutff_5/in_1')
// (11, 7, 'neigh_op_bot_4')
// (12, 5, 'neigh_op_tnl_4')
// (12, 6, 'neigh_op_lft_4')
// (12, 6, 'sp4_h_l_40')
// (12, 7, 'neigh_op_bnl_4')

wire n1123;
// (8, 6, 'neigh_op_tnr_0')
// (8, 7, 'neigh_op_rgt_0')
// (8, 8, 'neigh_op_bnr_0')
// (9, 6, 'local_g0_0')
// (9, 6, 'lutff_1/in_1')
// (9, 6, 'lutff_6/in_2')
// (9, 6, 'neigh_op_top_0')
// (9, 7, 'lutff_0/out')
// (9, 8, 'neigh_op_bot_0')
// (10, 6, 'neigh_op_tnl_0')
// (10, 7, 'neigh_op_lft_0')
// (10, 8, 'neigh_op_bnl_0')

wire n1124;
// (8, 6, 'neigh_op_tnr_7')
// (8, 7, 'neigh_op_rgt_7')
// (8, 8, 'neigh_op_bnr_7')
// (9, 6, 'neigh_op_top_7')
// (9, 7, 'lutff_7/out')
// (9, 8, 'local_g1_7')
// (9, 8, 'lutff_7/in_3')
// (9, 8, 'neigh_op_bot_7')
// (10, 6, 'neigh_op_tnl_7')
// (10, 7, 'neigh_op_lft_7')
// (10, 8, 'neigh_op_bnl_7')

reg n1125 = 0;
// (8, 6, 'sp4_h_r_1')
// (8, 7, 'sp4_r_v_b_38')
// (8, 8, 'sp4_r_v_b_27')
// (8, 9, 'sp4_r_v_b_14')
// (8, 10, 'sp4_r_v_b_3')
// (9, 6, 'local_g0_4')
// (9, 6, 'local_g1_0')
// (9, 6, 'lutff_2/in_2')
// (9, 6, 'lutff_5/in_0')
// (9, 6, 'lutff_7/in_1')
// (9, 6, 'sp4_h_r_12')
// (9, 6, 'sp4_h_r_3')
// (9, 6, 'sp4_h_r_8')
// (9, 6, 'sp4_v_t_38')
// (9, 7, 'local_g2_6')
// (9, 7, 'lutff_1/in_3')
// (9, 7, 'lutff_2/in_0')
// (9, 7, 'sp4_v_b_38')
// (9, 8, 'sp4_v_b_27')
// (9, 9, 'sp4_v_b_14')
// (9, 10, 'sp4_v_b_3')
// (10, 6, 'local_g0_5')
// (10, 6, 'lutff_1/in_2')
// (10, 6, 'sp4_h_r_14')
// (10, 6, 'sp4_h_r_21')
// (10, 6, 'sp4_h_r_25')
// (11, 2, 'sp4_h_r_8')
// (11, 4, 'local_g0_0')
// (11, 4, 'lutff_3/in_1')
// (11, 4, 'sp4_h_r_0')
// (11, 5, 'local_g1_3')
// (11, 5, 'lutff_1/in_3')
// (11, 5, 'lutff_2/in_0')
// (11, 5, 'lutff_7/in_1')
// (11, 5, 'sp4_h_r_11')
// (11, 6, 'local_g0_0')
// (11, 6, 'lutff_5/in_1')
// (11, 6, 'sp4_h_r_27')
// (11, 6, 'sp4_h_r_32')
// (11, 6, 'sp4_h_r_36')
// (11, 6, 'sp4_h_r_8')
// (12, 2, 'local_g0_5')
// (12, 2, 'lutff_6/in_3')
// (12, 2, 'sp4_h_r_21')
// (12, 3, 'sp4_r_v_b_40')
// (12, 4, 'local_g0_5')
// (12, 4, 'lutff_1/in_0')
// (12, 4, 'sp4_h_r_13')
// (12, 4, 'sp4_r_v_b_29')
// (12, 5, 'sp4_h_r_22')
// (12, 5, 'sp4_r_v_b_16')
// (12, 6, 'sp4_h_l_36')
// (12, 6, 'sp4_h_r_21')
// (12, 6, 'sp4_h_r_38')
// (12, 6, 'sp4_h_r_45')
// (12, 6, 'sp4_h_r_5')
// (12, 6, 'sp4_r_v_b_5')
// (12, 7, 'sp4_r_v_b_43')
// (12, 8, 'sp4_r_v_b_30')
// (12, 9, 'sp4_r_v_b_19')
// (12, 10, 'sp4_r_v_b_6')
// (12, 11, 'sp4_r_v_b_39')
// (12, 12, 'sp4_r_v_b_26')
// (12, 13, 'sp4_r_v_b_15')
// (12, 14, 'sp4_r_v_b_2')
// (12, 15, 'sp4_r_v_b_47')
// (12, 16, 'sp4_r_v_b_34')
// (12, 17, 'sp4_r_v_b_23')
// (12, 18, 'sp4_r_v_b_10')
// (13, 2, 'sp4_h_r_32')
// (13, 2, 'sp4_v_t_40')
// (13, 3, 'sp4_v_b_40')
// (13, 4, 'sp4_h_r_24')
// (13, 4, 'sp4_v_b_29')
// (13, 5, 'sp4_h_r_35')
// (13, 5, 'sp4_v_b_16')
// (13, 6, 'sp4_h_l_38')
// (13, 6, 'sp4_h_l_45')
// (13, 6, 'sp4_h_r_0')
// (13, 6, 'sp4_h_r_16')
// (13, 6, 'sp4_h_r_32')
// (13, 6, 'sp4_v_b_5')
// (13, 6, 'sp4_v_t_43')
// (13, 7, 'sp4_v_b_43')
// (13, 8, 'sp4_v_b_30')
// (13, 9, 'sp4_v_b_19')
// (13, 10, 'sp4_v_b_6')
// (13, 10, 'sp4_v_t_39')
// (13, 11, 'sp4_v_b_39')
// (13, 12, 'sp4_v_b_26')
// (13, 13, 'sp4_v_b_15')
// (13, 14, 'sp4_v_b_2')
// (13, 14, 'sp4_v_t_47')
// (13, 15, 'sp4_v_b_47')
// (13, 16, 'local_g2_2')
// (13, 16, 'lutff_6/in_0')
// (13, 16, 'lutff_7/in_1')
// (13, 16, 'sp4_v_b_34')
// (13, 17, 'sp4_v_b_23')
// (13, 18, 'sp4_v_b_10')
// (14, 1, 'sp4_r_v_b_17')
// (14, 2, 'local_g1_4')
// (14, 2, 'lutff_0/in_3')
// (14, 2, 'sp4_h_r_45')
// (14, 2, 'sp4_r_v_b_4')
// (14, 3, 'sp4_r_v_b_45')
// (14, 4, 'sp4_h_r_37')
// (14, 4, 'sp4_r_v_b_32')
// (14, 5, 'local_g2_4')
// (14, 5, 'lutff_2/in_0')
// (14, 5, 'lutff_5/in_1')
// (14, 5, 'neigh_op_tnr_4')
// (14, 5, 'sp4_h_r_46')
// (14, 5, 'sp4_r_v_b_21')
// (14, 5, 'sp4_r_v_b_37')
// (14, 6, 'neigh_op_rgt_4')
// (14, 6, 'sp4_h_r_13')
// (14, 6, 'sp4_h_r_29')
// (14, 6, 'sp4_h_r_45')
// (14, 6, 'sp4_r_v_b_24')
// (14, 6, 'sp4_r_v_b_40')
// (14, 6, 'sp4_r_v_b_8')
// (14, 7, 'neigh_op_bnr_4')
// (14, 7, 'sp4_r_v_b_13')
// (14, 7, 'sp4_r_v_b_29')
// (14, 8, 'sp4_r_v_b_0')
// (14, 8, 'sp4_r_v_b_16')
// (14, 9, 'sp4_r_v_b_5')
// (15, 0, 'span4_vert_17')
// (15, 1, 'sp4_v_b_17')
// (15, 2, 'sp4_h_l_45')
// (15, 2, 'sp4_v_b_4')
// (15, 2, 'sp4_v_t_45')
// (15, 3, 'sp4_v_b_45')
// (15, 4, 'sp4_h_l_37')
// (15, 4, 'sp4_v_b_32')
// (15, 4, 'sp4_v_t_37')
// (15, 5, 'local_g1_4')
// (15, 5, 'lutff_5/in_2')
// (15, 5, 'lutff_7/in_0')
// (15, 5, 'neigh_op_top_4')
// (15, 5, 'sp4_h_l_46')
// (15, 5, 'sp4_v_b_21')
// (15, 5, 'sp4_v_b_37')
// (15, 5, 'sp4_v_t_40')
// (15, 6, 'local_g0_4')
// (15, 6, 'lutff_4/in_0')
// (15, 6, 'lutff_4/out')
// (15, 6, 'sp4_h_l_45')
// (15, 6, 'sp4_h_r_24')
// (15, 6, 'sp4_h_r_40')
// (15, 6, 'sp4_h_r_8')
// (15, 6, 'sp4_v_b_24')
// (15, 6, 'sp4_v_b_40')
// (15, 6, 'sp4_v_b_8')
// (15, 7, 'neigh_op_bot_4')
// (15, 7, 'sp4_v_b_13')
// (15, 7, 'sp4_v_b_29')
// (15, 8, 'sp4_v_b_0')
// (15, 8, 'sp4_v_b_16')
// (15, 9, 'sp4_v_b_5')
// (16, 5, 'neigh_op_tnl_4')
// (16, 6, 'neigh_op_lft_4')
// (16, 6, 'sp4_h_l_40')
// (16, 6, 'sp4_h_r_21')
// (16, 6, 'sp4_h_r_37')
// (16, 7, 'neigh_op_bnl_4')
// (17, 6, 'local_g2_0')
// (17, 6, 'lutff_4/in_2')
// (17, 6, 'sp4_h_l_37')
// (17, 6, 'sp4_h_r_32')
// (18, 6, 'sp4_h_r_45')
// (19, 6, 'sp4_h_l_45')

reg n1126 = 0;
// (8, 6, 'sp4_h_r_11')
// (9, 6, 'local_g0_6')
// (9, 6, 'lutff_2/in_0')
// (9, 6, 'lutff_5/in_1')
// (9, 6, 'lutff_7/in_3')
// (9, 6, 'sp4_h_r_22')
// (9, 7, 'local_g2_7')
// (9, 7, 'lutff_1/in_0')
// (9, 7, 'lutff_2/in_1')
// (9, 7, 'sp4_r_v_b_39')
// (9, 8, 'sp4_r_v_b_26')
// (9, 9, 'sp4_r_v_b_15')
// (9, 10, 'sp4_r_v_b_2')
// (10, 6, 'local_g0_2')
// (10, 6, 'lutff_1/in_3')
// (10, 6, 'sp4_h_r_2')
// (10, 6, 'sp4_h_r_35')
// (10, 6, 'sp4_v_t_39')
// (10, 7, 'sp4_v_b_39')
// (10, 8, 'sp4_v_b_26')
// (10, 9, 'sp4_v_b_15')
// (10, 10, 'sp4_v_b_2')
// (11, 3, 'sp4_r_v_b_38')
// (11, 3, 'sp4_r_v_b_40')
// (11, 4, 'local_g1_3')
// (11, 4, 'lutff_3/in_3')
// (11, 4, 'sp4_r_v_b_27')
// (11, 4, 'sp4_r_v_b_29')
// (11, 5, 'local_g2_6')
// (11, 5, 'lutff_1/in_1')
// (11, 5, 'lutff_2/in_2')
// (11, 5, 'lutff_7/in_3')
// (11, 5, 'sp4_r_v_b_14')
// (11, 5, 'sp4_r_v_b_16')
// (11, 6, 'local_g3_6')
// (11, 6, 'lutff_5/in_0')
// (11, 6, 'sp4_h_r_15')
// (11, 6, 'sp4_h_r_46')
// (11, 6, 'sp4_r_v_b_3')
// (11, 6, 'sp4_r_v_b_5')
// (11, 16, 'sp4_h_r_3')
// (12, 2, 'local_g0_3')
// (12, 2, 'lutff_7/in_0')
// (12, 2, 'sp4_h_r_3')
// (12, 2, 'sp4_v_t_38')
// (12, 2, 'sp4_v_t_40')
// (12, 3, 'sp4_v_b_38')
// (12, 3, 'sp4_v_b_40')
// (12, 4, 'local_g3_5')
// (12, 4, 'lutff_1/in_3')
// (12, 4, 'sp4_v_b_27')
// (12, 4, 'sp4_v_b_29')
// (12, 5, 'sp4_v_b_14')
// (12, 5, 'sp4_v_b_16')
// (12, 6, 'sp4_h_l_46')
// (12, 6, 'sp4_h_r_26')
// (12, 6, 'sp4_h_r_3')
// (12, 6, 'sp4_v_b_3')
// (12, 6, 'sp4_v_b_5')
// (12, 16, 'sp4_h_r_14')
// (13, 2, 'sp4_h_r_14')
// (13, 6, 'sp4_h_r_14')
// (13, 6, 'sp4_h_r_39')
// (13, 16, 'local_g2_3')
// (13, 16, 'lutff_0/in_1')
// (13, 16, 'lutff_1/in_0')
// (13, 16, 'sp4_h_r_27')
// (14, 1, 'sp4_r_v_b_15')
// (14, 2, 'local_g1_2')
// (14, 2, 'lutff_0/in_1')
// (14, 2, 'sp4_h_r_27')
// (14, 2, 'sp4_r_v_b_2')
// (14, 3, 'sp4_r_v_b_43')
// (14, 4, 'sp4_r_v_b_30')
// (14, 5, 'local_g3_3')
// (14, 5, 'lutff_2/in_2')
// (14, 5, 'lutff_5/in_3')
// (14, 5, 'neigh_op_tnr_3')
// (14, 5, 'sp4_r_v_b_19')
// (14, 6, 'neigh_op_rgt_3')
// (14, 6, 'sp4_h_l_39')
// (14, 6, 'sp4_h_r_11')
// (14, 6, 'sp4_h_r_27')
// (14, 6, 'sp4_r_v_b_6')
// (14, 7, 'neigh_op_bnr_3')
// (14, 13, 'sp4_r_v_b_38')
// (14, 14, 'sp4_r_v_b_27')
// (14, 15, 'sp4_r_v_b_14')
// (14, 16, 'sp4_h_r_38')
// (14, 16, 'sp4_r_v_b_3')
// (15, 0, 'span4_vert_15')
// (15, 1, 'sp4_v_b_15')
// (15, 2, 'sp4_h_r_38')
// (15, 2, 'sp4_v_b_2')
// (15, 2, 'sp4_v_t_43')
// (15, 3, 'sp4_v_b_43')
// (15, 4, 'sp4_v_b_30')
// (15, 5, 'local_g0_3')
// (15, 5, 'lutff_5/in_0')
// (15, 5, 'lutff_7/in_2')
// (15, 5, 'neigh_op_top_3')
// (15, 5, 'sp12_v_t_22')
// (15, 5, 'sp4_v_b_19')
// (15, 6, 'local_g1_3')
// (15, 6, 'lutff_3/in_1')
// (15, 6, 'lutff_3/out')
// (15, 6, 'sp12_v_b_22')
// (15, 6, 'sp4_h_r_22')
// (15, 6, 'sp4_h_r_38')
// (15, 6, 'sp4_v_b_6')
// (15, 7, 'neigh_op_bot_3')
// (15, 7, 'sp12_v_b_21')
// (15, 8, 'sp12_v_b_18')
// (15, 9, 'sp12_v_b_17')
// (15, 10, 'sp12_v_b_14')
// (15, 11, 'sp12_v_b_13')
// (15, 12, 'sp12_v_b_10')
// (15, 12, 'sp4_v_t_38')
// (15, 13, 'sp12_v_b_9')
// (15, 13, 'sp4_v_b_38')
// (15, 14, 'sp12_v_b_6')
// (15, 14, 'sp4_v_b_27')
// (15, 15, 'sp12_v_b_5')
// (15, 15, 'sp4_v_b_14')
// (15, 16, 'sp12_v_b_2')
// (15, 16, 'sp4_h_l_38')
// (15, 16, 'sp4_v_b_3')
// (15, 17, 'sp12_v_b_1')
// (16, 2, 'sp4_h_l_38')
// (16, 5, 'neigh_op_tnl_3')
// (16, 6, 'neigh_op_lft_3')
// (16, 6, 'sp4_h_l_38')
// (16, 6, 'sp4_h_r_35')
// (16, 7, 'neigh_op_bnl_3')
// (17, 6, 'local_g2_6')
// (17, 6, 'lutff_6/in_2')
// (17, 6, 'sp4_h_r_46')
// (18, 6, 'sp4_h_l_46')

wire n1127;
// (8, 7, 'lutff_5/cout')
// (8, 7, 'lutff_6/in_3')

wire n1128;
// (8, 7, 'neigh_op_tnr_0')
// (8, 8, 'neigh_op_rgt_0')
// (8, 9, 'neigh_op_bnr_0')
// (9, 7, 'neigh_op_top_0')
// (9, 8, 'local_g0_0')
// (9, 8, 'lutff_0/out')
// (9, 8, 'lutff_2/in_0')
// (9, 8, 'lutff_4/in_2')
// (9, 9, 'neigh_op_bot_0')
// (10, 7, 'neigh_op_tnl_0')
// (10, 8, 'neigh_op_lft_0')
// (10, 9, 'neigh_op_bnl_0')

reg n1129 = 0;
// (8, 7, 'neigh_op_tnr_2')
// (8, 8, 'neigh_op_rgt_2')
// (8, 9, 'neigh_op_bnr_2')
// (9, 7, 'neigh_op_top_2')
// (9, 8, 'lutff_2/out')
// (9, 9, 'local_g0_2')
// (9, 9, 'lutff_5/in_1')
// (9, 9, 'neigh_op_bot_2')
// (10, 7, 'neigh_op_tnl_2')
// (10, 8, 'neigh_op_lft_2')
// (10, 9, 'neigh_op_bnl_2')

reg n1130 = 0;
// (8, 7, 'neigh_op_tnr_3')
// (8, 8, 'neigh_op_rgt_3')
// (8, 9, 'neigh_op_bnr_3')
// (9, 7, 'neigh_op_top_3')
// (9, 8, 'lutff_3/out')
// (9, 9, 'neigh_op_bot_3')
// (10, 7, 'neigh_op_tnl_3')
// (10, 8, 'local_g1_3')
// (10, 8, 'lutff_1/in_3')
// (10, 8, 'neigh_op_lft_3')
// (10, 9, 'neigh_op_bnl_3')

reg n1131 = 0;
// (8, 7, 'neigh_op_tnr_4')
// (8, 8, 'neigh_op_rgt_4')
// (8, 9, 'neigh_op_bnr_4')
// (9, 7, 'neigh_op_top_4')
// (9, 8, 'lutff_4/out')
// (9, 9, 'neigh_op_bot_4')
// (10, 7, 'neigh_op_tnl_4')
// (10, 8, 'neigh_op_lft_4')
// (10, 9, 'local_g3_4')
// (10, 9, 'lutff_7/in_0')
// (10, 9, 'neigh_op_bnl_4')

wire n1132;
// (8, 7, 'neigh_op_tnr_5')
// (8, 8, 'neigh_op_rgt_5')
// (8, 9, 'neigh_op_bnr_5')
// (9, 7, 'neigh_op_top_5')
// (9, 8, 'lutff_5/out')
// (9, 9, 'neigh_op_bot_5')
// (10, 7, 'neigh_op_tnl_5')
// (10, 8, 'local_g0_5')
// (10, 8, 'lutff_5/in_0')
// (10, 8, 'neigh_op_lft_5')
// (10, 9, 'neigh_op_bnl_5')

reg n1133 = 0;
// (8, 7, 'neigh_op_tnr_6')
// (8, 8, 'neigh_op_rgt_6')
// (8, 9, 'neigh_op_bnr_6')
// (9, 7, 'neigh_op_top_6')
// (9, 8, 'local_g3_6')
// (9, 8, 'lutff_5/in_2')
// (9, 8, 'lutff_6/out')
// (9, 9, 'neigh_op_bot_6')
// (10, 7, 'neigh_op_tnl_6')
// (10, 8, 'neigh_op_lft_6')
// (10, 9, 'neigh_op_bnl_6')

reg n1134 = 0;
// (8, 7, 'neigh_op_tnr_7')
// (8, 7, 'sp4_r_v_b_43')
// (8, 8, 'neigh_op_rgt_7')
// (8, 8, 'sp4_r_v_b_30')
// (8, 9, 'neigh_op_bnr_7')
// (8, 9, 'sp4_r_v_b_19')
// (8, 10, 'local_g1_6')
// (8, 10, 'lutff_6/in_1')
// (8, 10, 'sp4_r_v_b_6')
// (9, 6, 'sp4_v_t_43')
// (9, 7, 'neigh_op_top_7')
// (9, 7, 'sp4_v_b_43')
// (9, 8, 'lutff_7/out')
// (9, 8, 'sp4_v_b_30')
// (9, 9, 'neigh_op_bot_7')
// (9, 9, 'sp4_v_b_19')
// (9, 10, 'sp4_v_b_6')
// (10, 7, 'neigh_op_tnl_7')
// (10, 8, 'neigh_op_lft_7')
// (10, 9, 'neigh_op_bnl_7')

reg n1135 = 0;
// (8, 7, 'sp4_h_r_3')
// (9, 7, 'sp4_h_r_14')
// (10, 7, 'local_g2_3')
// (10, 7, 'lutff_2/in_1')
// (10, 7, 'sp4_h_r_27')
// (11, 5, 'sp4_r_v_b_39')
// (11, 6, 'sp4_r_v_b_26')
// (11, 7, 'sp4_h_r_38')
// (11, 7, 'sp4_r_v_b_15')
// (11, 8, 'sp4_r_v_b_2')
// (11, 8, 'sp4_r_v_b_38')
// (11, 9, 'local_g3_7')
// (11, 9, 'lutff_4/in_2')
// (11, 9, 'neigh_op_tnr_7')
// (11, 9, 'sp4_r_v_b_27')
// (11, 9, 'sp4_r_v_b_43')
// (11, 10, 'neigh_op_rgt_7')
// (11, 10, 'sp4_r_v_b_14')
// (11, 10, 'sp4_r_v_b_30')
// (11, 11, 'neigh_op_bnr_7')
// (11, 11, 'sp4_r_v_b_19')
// (11, 11, 'sp4_r_v_b_3')
// (11, 12, 'sp4_r_v_b_6')
// (12, 4, 'sp4_v_t_39')
// (12, 5, 'sp4_v_b_39')
// (12, 6, 'sp4_v_b_26')
// (12, 7, 'local_g0_7')
// (12, 7, 'lutff_1/in_0')
// (12, 7, 'sp4_h_l_38')
// (12, 7, 'sp4_v_b_15')
// (12, 7, 'sp4_v_t_38')
// (12, 8, 'sp4_v_b_2')
// (12, 8, 'sp4_v_b_38')
// (12, 8, 'sp4_v_t_43')
// (12, 9, 'local_g0_7')
// (12, 9, 'lutff_5/in_2')
// (12, 9, 'neigh_op_top_7')
// (12, 9, 'sp4_v_b_27')
// (12, 9, 'sp4_v_b_43')
// (12, 10, 'lutff_7/out')
// (12, 10, 'sp4_v_b_14')
// (12, 10, 'sp4_v_b_30')
// (12, 11, 'neigh_op_bot_7')
// (12, 11, 'sp4_v_b_19')
// (12, 11, 'sp4_v_b_3')
// (12, 12, 'sp4_v_b_6')
// (13, 9, 'neigh_op_tnl_7')
// (13, 10, 'neigh_op_lft_7')
// (13, 11, 'neigh_op_bnl_7')

wire n1136;
// (8, 8, 'neigh_op_tnr_0')
// (8, 9, 'neigh_op_rgt_0')
// (8, 10, 'neigh_op_bnr_0')
// (9, 8, 'neigh_op_top_0')
// (9, 9, 'local_g3_0')
// (9, 9, 'lutff_0/out')
// (9, 9, 'lutff_7/in_0')
// (9, 10, 'neigh_op_bot_0')
// (10, 8, 'neigh_op_tnl_0')
// (10, 9, 'neigh_op_lft_0')
// (10, 10, 'neigh_op_bnl_0')

reg n1137 = 0;
// (8, 8, 'neigh_op_tnr_1')
// (8, 9, 'neigh_op_rgt_1')
// (8, 10, 'neigh_op_bnr_1')
// (9, 6, 'sp12_v_t_22')
// (9, 7, 'sp12_v_b_22')
// (9, 8, 'neigh_op_top_1')
// (9, 8, 'sp12_v_b_21')
// (9, 9, 'lutff_1/out')
// (9, 9, 'sp12_v_b_18')
// (9, 10, 'neigh_op_bot_1')
// (9, 10, 'sp12_v_b_17')
// (9, 11, 'sp12_v_b_14')
// (9, 12, 'sp12_v_b_13')
// (9, 13, 'sp12_v_b_10')
// (9, 14, 'sp12_v_b_9')
// (9, 15, 'local_g2_6')
// (9, 15, 'lutff_2/in_0')
// (9, 15, 'sp12_v_b_6')
// (9, 16, 'sp12_v_b_5')
// (9, 17, 'sp12_v_b_2')
// (9, 18, 'sp12_v_b_1')
// (10, 8, 'neigh_op_tnl_1')
// (10, 9, 'neigh_op_lft_1')
// (10, 10, 'neigh_op_bnl_1')

wire n1138;
// (8, 8, 'neigh_op_tnr_2')
// (8, 9, 'neigh_op_rgt_2')
// (8, 10, 'neigh_op_bnr_2')
// (9, 8, 'neigh_op_top_2')
// (9, 9, 'lutff_2/out')
// (9, 10, 'local_g1_2')
// (9, 10, 'lutff_7/in_2')
// (9, 10, 'neigh_op_bot_2')
// (10, 8, 'neigh_op_tnl_2')
// (10, 9, 'neigh_op_lft_2')
// (10, 10, 'neigh_op_bnl_2')

reg n1139 = 0;
// (8, 8, 'neigh_op_tnr_3')
// (8, 9, 'neigh_op_rgt_3')
// (8, 10, 'neigh_op_bnr_3')
// (9, 8, 'neigh_op_top_3')
// (9, 9, 'local_g0_3')
// (9, 9, 'lutff_2/in_1')
// (9, 9, 'lutff_3/out')
// (9, 10, 'neigh_op_bot_3')
// (10, 8, 'neigh_op_tnl_3')
// (10, 9, 'neigh_op_lft_3')
// (10, 10, 'neigh_op_bnl_3')

reg n1140 = 0;
// (8, 8, 'neigh_op_tnr_4')
// (8, 9, 'neigh_op_rgt_4')
// (8, 10, 'neigh_op_bnr_4')
// (9, 8, 'neigh_op_top_4')
// (9, 9, 'local_g2_4')
// (9, 9, 'lutff_2/in_2')
// (9, 9, 'lutff_4/out')
// (9, 10, 'neigh_op_bot_4')
// (10, 8, 'neigh_op_tnl_4')
// (10, 9, 'neigh_op_lft_4')
// (10, 10, 'neigh_op_bnl_4')

wire n1141;
// (8, 8, 'neigh_op_tnr_5')
// (8, 9, 'neigh_op_rgt_5')
// (8, 9, 'sp4_r_v_b_42')
// (8, 10, 'neigh_op_bnr_5')
// (8, 10, 'sp4_r_v_b_31')
// (8, 11, 'sp4_r_v_b_18')
// (8, 12, 'sp4_r_v_b_7')
// (9, 8, 'neigh_op_top_5')
// (9, 8, 'sp4_v_t_42')
// (9, 9, 'lutff_5/out')
// (9, 9, 'sp4_v_b_42')
// (9, 10, 'neigh_op_bot_5')
// (9, 10, 'sp4_v_b_31')
// (9, 11, 'sp4_v_b_18')
// (9, 12, 'local_g0_7')
// (9, 12, 'lutff_3/in_2')
// (9, 12, 'sp4_v_b_7')
// (10, 8, 'neigh_op_tnl_5')
// (10, 9, 'neigh_op_lft_5')
// (10, 10, 'neigh_op_bnl_5')

reg n1142 = 0;
// (8, 8, 'neigh_op_tnr_6')
// (8, 9, 'neigh_op_rgt_6')
// (8, 10, 'neigh_op_bnr_6')
// (9, 3, 'sp12_v_t_23')
// (9, 4, 'sp12_v_b_23')
// (9, 5, 'sp12_v_b_20')
// (9, 6, 'sp12_v_b_19')
// (9, 7, 'sp12_v_b_16')
// (9, 8, 'neigh_op_top_6')
// (9, 8, 'sp12_v_b_15')
// (9, 9, 'lutff_6/out')
// (9, 9, 'sp12_v_b_12')
// (9, 10, 'neigh_op_bot_6')
// (9, 10, 'sp12_v_b_11')
// (9, 11, 'sp12_v_b_8')
// (9, 12, 'sp12_v_b_7')
// (9, 13, 'sp12_v_b_4')
// (9, 14, 'local_g3_3')
// (9, 14, 'lutff_1/in_3')
// (9, 14, 'sp12_v_b_3')
// (9, 15, 'sp12_v_b_0')
// (10, 8, 'neigh_op_tnl_6')
// (10, 9, 'neigh_op_lft_6')
// (10, 10, 'neigh_op_bnl_6')

reg n1143 = 0;
// (8, 8, 'neigh_op_tnr_7')
// (8, 9, 'neigh_op_rgt_7')
// (8, 10, 'neigh_op_bnr_7')
// (9, 8, 'neigh_op_top_7')
// (9, 9, 'lutff_7/out')
// (9, 10, 'local_g0_7')
// (9, 10, 'lutff_2/in_3')
// (9, 10, 'neigh_op_bot_7')
// (10, 8, 'neigh_op_tnl_7')
// (10, 9, 'neigh_op_lft_7')
// (10, 10, 'neigh_op_bnl_7')

reg n1144 = 0;
// (8, 8, 'sp4_r_v_b_44')
// (8, 9, 'sp4_r_v_b_33')
// (8, 10, 'sp4_r_v_b_20')
// (8, 11, 'sp4_r_v_b_9')
// (8, 12, 'sp4_r_v_b_44')
// (8, 13, 'neigh_op_tnr_2')
// (8, 13, 'sp4_r_v_b_33')
// (8, 14, 'neigh_op_rgt_2')
// (8, 14, 'sp4_r_v_b_20')
// (8, 15, 'neigh_op_bnr_2')
// (8, 15, 'sp4_r_v_b_9')
// (9, 7, 'sp4_v_t_44')
// (9, 8, 'sp4_v_b_44')
// (9, 9, 'sp4_v_b_33')
// (9, 10, 'local_g1_4')
// (9, 10, 'lutff_6/in_3')
// (9, 10, 'sp4_v_b_20')
// (9, 11, 'sp4_v_b_9')
// (9, 11, 'sp4_v_t_44')
// (9, 12, 'sp4_v_b_44')
// (9, 13, 'neigh_op_top_2')
// (9, 13, 'sp4_v_b_33')
// (9, 14, 'lutff_2/out')
// (9, 14, 'sp4_v_b_20')
// (9, 15, 'local_g1_2')
// (9, 15, 'lutff_6/in_1')
// (9, 15, 'neigh_op_bot_2')
// (9, 15, 'sp4_v_b_9')
// (10, 13, 'neigh_op_tnl_2')
// (10, 14, 'neigh_op_lft_2')
// (10, 15, 'neigh_op_bnl_2')

reg n1145 = 0;
// (8, 8, 'sp4_r_v_b_45')
// (8, 9, 'sp4_r_v_b_32')
// (8, 10, 'sp4_r_v_b_21')
// (8, 11, 'local_g2_0')
// (8, 11, 'lutff_4/in_2')
// (8, 11, 'sp4_r_v_b_8')
// (9, 7, 'sp4_h_r_8')
// (9, 7, 'sp4_v_t_45')
// (9, 8, 'sp4_v_b_45')
// (9, 9, 'sp4_v_b_32')
// (9, 10, 'sp4_v_b_21')
// (9, 11, 'sp4_v_b_8')
// (10, 6, 'neigh_op_tnr_0')
// (10, 7, 'neigh_op_rgt_0')
// (10, 7, 'sp4_h_r_21')
// (10, 8, 'neigh_op_bnr_0')
// (11, 6, 'neigh_op_top_0')
// (11, 7, 'lutff_0/out')
// (11, 7, 'sp4_h_r_32')
// (11, 8, 'neigh_op_bot_0')
// (12, 6, 'neigh_op_tnl_0')
// (12, 7, 'neigh_op_lft_0')
// (12, 7, 'sp4_h_r_45')
// (12, 8, 'neigh_op_bnl_0')
// (13, 7, 'sp4_h_l_45')

wire n1146;
// (8, 8, 'sp4_r_v_b_47')
// (8, 9, 'sp4_r_v_b_34')
// (8, 10, 'sp4_r_v_b_23')
// (8, 11, 'sp4_r_v_b_10')
// (8, 12, 'sp4_r_v_b_43')
// (8, 13, 'sp4_r_v_b_30')
// (8, 14, 'sp4_r_v_b_19')
// (8, 15, 'sp4_r_v_b_6')
// (9, 7, 'sp4_h_r_4')
// (9, 7, 'sp4_v_t_47')
// (9, 8, 'sp4_r_v_b_36')
// (9, 8, 'sp4_v_b_47')
// (9, 9, 'local_g1_1')
// (9, 9, 'local_g3_2')
// (9, 9, 'lutff_1/in_2')
// (9, 9, 'lutff_6/in_0')
// (9, 9, 'sp4_r_v_b_25')
// (9, 9, 'sp4_v_b_34')
// (9, 10, 'local_g1_7')
// (9, 10, 'lutff_5/in_3')
// (9, 10, 'lutff_6/in_2')
// (9, 10, 'sp4_r_v_b_12')
// (9, 10, 'sp4_v_b_23')
// (9, 11, 'local_g0_2')
// (9, 11, 'lutff_7/in_1')
// (9, 11, 'sp4_r_v_b_1')
// (9, 11, 'sp4_v_b_10')
// (9, 11, 'sp4_v_t_43')
// (9, 12, 'sp4_v_b_43')
// (9, 13, 'local_g3_6')
// (9, 13, 'lutff_2/in_3')
// (9, 13, 'sp4_v_b_30')
// (9, 14, 'sp4_v_b_19')
// (9, 15, 'local_g1_6')
// (9, 15, 'lutff_3/in_0')
// (9, 15, 'lutff_5/in_2')
// (9, 15, 'sp4_v_b_6')
// (10, 6, 'neigh_op_tnr_6')
// (10, 6, 'sp4_r_v_b_41')
// (10, 7, 'local_g3_6')
// (10, 7, 'lutff_1/in_2')
// (10, 7, 'lutff_5/in_0')
// (10, 7, 'lutff_6/in_1')
// (10, 7, 'neigh_op_rgt_6')
// (10, 7, 'sp4_h_r_1')
// (10, 7, 'sp4_h_r_17')
// (10, 7, 'sp4_r_v_b_28')
// (10, 7, 'sp4_r_v_b_44')
// (10, 7, 'sp4_v_t_36')
// (10, 8, 'local_g1_6')
// (10, 8, 'lutff_3/in_0')
// (10, 8, 'lutff_4/in_1')
// (10, 8, 'neigh_op_bnr_6')
// (10, 8, 'sp4_r_v_b_17')
// (10, 8, 'sp4_r_v_b_33')
// (10, 8, 'sp4_v_b_36')
// (10, 9, 'local_g1_4')
// (10, 9, 'lutff_5/in_0')
// (10, 9, 'sp4_r_v_b_20')
// (10, 9, 'sp4_r_v_b_4')
// (10, 9, 'sp4_v_b_25')
// (10, 10, 'local_g2_1')
// (10, 10, 'lutff_1/in_0')
// (10, 10, 'lutff_2/in_1')
// (10, 10, 'sp4_r_v_b_9')
// (10, 10, 'sp4_v_b_12')
// (10, 11, 'sp4_r_v_b_44')
// (10, 11, 'sp4_v_b_1')
// (10, 12, 'sp4_r_v_b_33')
// (10, 13, 'local_g3_4')
// (10, 13, 'lutff_2/in_1')
// (10, 13, 'lutff_7/in_2')
// (10, 13, 'sp4_r_v_b_20')
// (10, 14, 'sp4_r_v_b_9')
// (11, 5, 'sp4_v_t_41')
// (11, 6, 'neigh_op_top_6')
// (11, 6, 'sp4_v_b_41')
// (11, 6, 'sp4_v_t_44')
// (11, 7, 'local_g1_6')
// (11, 7, 'lutff_4/in_3')
// (11, 7, 'lutff_6/out')
// (11, 7, 'sp4_h_r_12')
// (11, 7, 'sp4_h_r_28')
// (11, 7, 'sp4_v_b_28')
// (11, 7, 'sp4_v_b_44')
// (11, 8, 'local_g0_6')
// (11, 8, 'lutff_2/in_2')
// (11, 8, 'lutff_3/in_3')
// (11, 8, 'lutff_4/in_0')
// (11, 8, 'lutff_5/in_3')
// (11, 8, 'lutff_6/in_0')
// (11, 8, 'lutff_7/in_1')
// (11, 8, 'neigh_op_bot_6')
// (11, 8, 'sp4_v_b_17')
// (11, 8, 'sp4_v_b_33')
// (11, 9, 'local_g1_4')
// (11, 9, 'lutff_1/in_0')
// (11, 9, 'lutff_4/in_1')
// (11, 9, 'sp4_v_b_20')
// (11, 9, 'sp4_v_b_4')
// (11, 10, 'local_g1_1')
// (11, 10, 'lutff_0/in_2')
// (11, 10, 'sp4_v_b_9')
// (11, 10, 'sp4_v_t_44')
// (11, 11, 'sp4_v_b_44')
// (11, 12, 'sp4_v_b_33')
// (11, 13, 'sp4_v_b_20')
// (11, 14, 'local_g1_1')
// (11, 14, 'lutff_2/in_0')
// (11, 14, 'sp4_v_b_9')
// (12, 6, 'neigh_op_tnl_6')
// (12, 7, 'neigh_op_lft_6')
// (12, 7, 'sp4_h_r_25')
// (12, 7, 'sp4_h_r_41')
// (12, 8, 'neigh_op_bnl_6')
// (13, 7, 'sp4_h_l_41')
// (13, 7, 'sp4_h_r_36')
// (14, 7, 'sp4_h_l_36')

wire n1147;
// (8, 9, 'lutff_1/cout')
// (8, 9, 'lutff_2/in_3')

wire n1148;
// (8, 9, 'lutff_2/cout')
// (8, 9, 'lutff_3/in_3')

wire n1149;
// (8, 9, 'lutff_3/cout')
// (8, 9, 'lutff_4/in_3')

wire n1150;
// (8, 9, 'lutff_4/cout')
// (8, 9, 'lutff_5/in_3')

reg n1151 = 0;
// (8, 9, 'neigh_op_tnr_0')
// (8, 10, 'neigh_op_rgt_0')
// (8, 11, 'neigh_op_bnr_0')
// (9, 9, 'neigh_op_top_0')
// (9, 10, 'lutff_0/out')
// (9, 11, 'local_g1_0')
// (9, 11, 'lutff_3/in_2')
// (9, 11, 'neigh_op_bot_0')
// (10, 9, 'neigh_op_tnl_0')
// (10, 10, 'neigh_op_lft_0')
// (10, 11, 'neigh_op_bnl_0')

reg n1152 = 0;
// (8, 9, 'neigh_op_tnr_1')
// (8, 10, 'neigh_op_rgt_1')
// (8, 11, 'neigh_op_bnr_1')
// (9, 9, 'neigh_op_top_1')
// (9, 10, 'local_g3_1')
// (9, 10, 'lutff_1/out')
// (9, 10, 'lutff_2/in_0')
// (9, 11, 'neigh_op_bot_1')
// (10, 9, 'neigh_op_tnl_1')
// (10, 10, 'neigh_op_lft_1')
// (10, 11, 'neigh_op_bnl_1')

wire n1153;
// (8, 9, 'neigh_op_tnr_2')
// (8, 10, 'neigh_op_rgt_2')
// (8, 11, 'neigh_op_bnr_2')
// (9, 9, 'local_g1_2')
// (9, 9, 'lutff_2/in_3')
// (9, 9, 'neigh_op_top_2')
// (9, 10, 'lutff_2/out')
// (9, 11, 'neigh_op_bot_2')
// (10, 9, 'neigh_op_tnl_2')
// (10, 10, 'neigh_op_lft_2')
// (10, 11, 'neigh_op_bnl_2')

reg n1154 = 0;
// (8, 9, 'neigh_op_tnr_3')
// (8, 10, 'neigh_op_rgt_3')
// (8, 11, 'neigh_op_bnr_3')
// (9, 9, 'neigh_op_top_3')
// (9, 10, 'local_g2_3')
// (9, 10, 'lutff_3/out')
// (9, 10, 'lutff_4/in_1')
// (9, 11, 'neigh_op_bot_3')
// (10, 9, 'neigh_op_tnl_3')
// (10, 10, 'neigh_op_lft_3')
// (10, 11, 'neigh_op_bnl_3')

wire n1155;
// (8, 9, 'neigh_op_tnr_4')
// (8, 10, 'neigh_op_rgt_4')
// (8, 11, 'neigh_op_bnr_4')
// (9, 9, 'local_g1_4')
// (9, 9, 'lutff_5/in_0')
// (9, 9, 'neigh_op_top_4')
// (9, 10, 'lutff_4/out')
// (9, 11, 'neigh_op_bot_4')
// (10, 9, 'neigh_op_tnl_4')
// (10, 10, 'neigh_op_lft_4')
// (10, 11, 'neigh_op_bnl_4')

reg n1156 = 0;
// (8, 9, 'neigh_op_tnr_5')
// (8, 10, 'neigh_op_rgt_5')
// (8, 11, 'neigh_op_bnr_5')
// (9, 9, 'neigh_op_top_5')
// (9, 10, 'lutff_5/out')
// (9, 11, 'local_g0_5')
// (9, 11, 'lutff_5/in_0')
// (9, 11, 'neigh_op_bot_5')
// (10, 9, 'neigh_op_tnl_5')
// (10, 10, 'neigh_op_lft_5')
// (10, 11, 'neigh_op_bnl_5')

reg n1157 = 0;
// (8, 9, 'neigh_op_tnr_6')
// (8, 10, 'neigh_op_rgt_6')
// (8, 11, 'neigh_op_bnr_6')
// (9, 9, 'neigh_op_top_6')
// (9, 10, 'local_g2_6')
// (9, 10, 'lutff_6/out')
// (9, 10, 'lutff_7/in_1')
// (9, 11, 'neigh_op_bot_6')
// (10, 9, 'neigh_op_tnl_6')
// (10, 10, 'neigh_op_lft_6')
// (10, 11, 'neigh_op_bnl_6')

wire n1158;
// (8, 9, 'neigh_op_tnr_7')
// (8, 10, 'neigh_op_rgt_7')
// (8, 11, 'neigh_op_bnr_7')
// (9, 9, 'neigh_op_top_7')
// (9, 10, 'lutff_7/out')
// (9, 11, 'neigh_op_bot_7')
// (10, 9, 'neigh_op_tnl_7')
// (10, 10, 'local_g0_7')
// (10, 10, 'lutff_5/in_2')
// (10, 10, 'neigh_op_lft_7')
// (10, 11, 'neigh_op_bnl_7')

reg n1159 = 0;
// (8, 10, 'neigh_op_tnr_1')
// (8, 11, 'neigh_op_rgt_1')
// (8, 12, 'neigh_op_bnr_1')
// (9, 10, 'neigh_op_top_1')
// (9, 11, 'local_g1_1')
// (9, 11, 'lutff_1/out')
// (9, 11, 'lutff_5/in_1')
// (9, 12, 'neigh_op_bot_1')
// (10, 10, 'neigh_op_tnl_1')
// (10, 11, 'neigh_op_lft_1')
// (10, 12, 'neigh_op_bnl_1')

reg n1160 = 0;
// (8, 10, 'neigh_op_tnr_2')
// (8, 11, 'neigh_op_rgt_2')
// (8, 12, 'neigh_op_bnr_2')
// (9, 10, 'neigh_op_top_2')
// (9, 11, 'local_g3_2')
// (9, 11, 'lutff_2/out')
// (9, 11, 'lutff_3/in_0')
// (9, 12, 'neigh_op_bot_2')
// (10, 10, 'neigh_op_tnl_2')
// (10, 11, 'neigh_op_lft_2')
// (10, 12, 'neigh_op_bnl_2')

wire n1161;
// (8, 10, 'neigh_op_tnr_3')
// (8, 11, 'neigh_op_rgt_3')
// (8, 12, 'neigh_op_bnr_3')
// (9, 10, 'neigh_op_top_3')
// (9, 11, 'lutff_3/out')
// (9, 12, 'neigh_op_bot_3')
// (10, 10, 'neigh_op_tnl_3')
// (10, 11, 'neigh_op_lft_3')
// (10, 12, 'local_g2_3')
// (10, 12, 'lutff_4/in_3')
// (10, 12, 'neigh_op_bnl_3')

reg n1162 = 0;
// (8, 10, 'neigh_op_tnr_4')
// (8, 11, 'neigh_op_rgt_4')
// (8, 12, 'neigh_op_bnr_4')
// (9, 10, 'neigh_op_top_4')
// (9, 11, 'local_g0_4')
// (9, 11, 'lutff_3/in_1')
// (9, 11, 'lutff_4/out')
// (9, 12, 'neigh_op_bot_4')
// (10, 10, 'neigh_op_tnl_4')
// (10, 11, 'neigh_op_lft_4')
// (10, 12, 'neigh_op_bnl_4')

wire n1163;
// (8, 10, 'neigh_op_tnr_5')
// (8, 11, 'neigh_op_rgt_5')
// (8, 12, 'neigh_op_bnr_5')
// (9, 10, 'neigh_op_top_5')
// (9, 11, 'lutff_5/out')
// (9, 12, 'neigh_op_bot_5')
// (10, 10, 'neigh_op_tnl_5')
// (10, 11, 'local_g0_5')
// (10, 11, 'lutff_4/in_3')
// (10, 11, 'neigh_op_lft_5')
// (10, 12, 'neigh_op_bnl_5')

wire n1164;
// (8, 10, 'neigh_op_tnr_6')
// (8, 11, 'neigh_op_rgt_6')
// (8, 12, 'neigh_op_bnr_6')
// (9, 10, 'neigh_op_top_6')
// (9, 10, 'sp4_r_v_b_40')
// (9, 11, 'lutff_6/out')
// (9, 11, 'sp4_r_v_b_29')
// (9, 12, 'neigh_op_bot_6')
// (9, 12, 'sp4_r_v_b_16')
// (9, 13, 'sp4_r_v_b_5')
// (10, 9, 'sp4_h_r_10')
// (10, 9, 'sp4_v_t_40')
// (10, 10, 'neigh_op_tnl_6')
// (10, 10, 'sp4_v_b_40')
// (10, 11, 'neigh_op_lft_6')
// (10, 11, 'sp4_v_b_29')
// (10, 12, 'neigh_op_bnl_6')
// (10, 12, 'sp4_v_b_16')
// (10, 13, 'sp4_v_b_5')
// (11, 9, 'sp4_h_r_23')
// (12, 9, 'local_g2_2')
// (12, 9, 'lutff_global/cen')
// (12, 9, 'sp4_h_r_34')
// (13, 9, 'sp4_h_r_47')
// (14, 9, 'sp4_h_l_47')

reg n1165 = 0;
// (8, 10, 'neigh_op_tnr_7')
// (8, 11, 'neigh_op_rgt_7')
// (8, 12, 'neigh_op_bnr_7')
// (9, 10, 'neigh_op_top_7')
// (9, 11, 'local_g2_7')
// (9, 11, 'lutff_5/in_2')
// (9, 11, 'lutff_7/out')
// (9, 12, 'neigh_op_bot_7')
// (10, 10, 'neigh_op_tnl_7')
// (10, 11, 'neigh_op_lft_7')
// (10, 12, 'neigh_op_bnl_7')

wire n1166;
// (8, 10, 'sp4_r_v_b_38')
// (8, 11, 'neigh_op_tnr_7')
// (8, 11, 'sp4_r_v_b_27')
// (8, 12, 'local_g1_3')
// (8, 12, 'lutff_global/cen')
// (8, 12, 'neigh_op_rgt_7')
// (8, 12, 'sp4_h_r_3')
// (8, 12, 'sp4_r_v_b_14')
// (8, 13, 'local_g1_3')
// (8, 13, 'lutff_global/cen')
// (8, 13, 'neigh_op_bnr_7')
// (8, 13, 'sp4_r_v_b_3')
// (9, 9, 'sp4_v_t_38')
// (9, 10, 'sp4_v_b_38')
// (9, 11, 'neigh_op_top_7')
// (9, 11, 'sp4_v_b_27')
// (9, 12, 'lutff_7/out')
// (9, 12, 'sp4_h_r_14')
// (9, 12, 'sp4_v_b_14')
// (9, 13, 'neigh_op_bot_7')
// (9, 13, 'sp4_v_b_3')
// (10, 11, 'neigh_op_tnl_7')
// (10, 12, 'neigh_op_lft_7')
// (10, 12, 'sp4_h_r_27')
// (10, 13, 'neigh_op_bnl_7')
// (11, 12, 'sp4_h_r_38')
// (12, 12, 'sp4_h_l_38')

reg n1167 = 0;
// (8, 10, 'sp4_r_v_b_47')
// (8, 11, 'sp4_r_v_b_34')
// (8, 12, 'sp4_r_v_b_23')
// (8, 13, 'local_g2_2')
// (8, 13, 'lutff_7/in_1')
// (8, 13, 'sp4_r_v_b_10')
// (9, 9, 'sp4_h_r_10')
// (9, 9, 'sp4_v_t_47')
// (9, 10, 'sp4_v_b_47')
// (9, 11, 'sp4_v_b_34')
// (9, 12, 'sp4_v_b_23')
// (9, 13, 'sp4_v_b_10')
// (10, 9, 'sp4_h_r_23')
// (11, 9, 'sp4_h_r_34')
// (12, 6, 'neigh_op_tnr_1')
// (12, 6, 'sp4_r_v_b_47')
// (12, 7, 'neigh_op_rgt_1')
// (12, 7, 'sp4_r_v_b_34')
// (12, 8, 'neigh_op_bnr_1')
// (12, 8, 'sp4_r_v_b_23')
// (12, 9, 'sp4_h_r_47')
// (12, 9, 'sp4_r_v_b_10')
// (13, 5, 'sp4_v_t_47')
// (13, 6, 'neigh_op_top_1')
// (13, 6, 'sp4_v_b_47')
// (13, 7, 'lutff_1/out')
// (13, 7, 'sp4_v_b_34')
// (13, 8, 'neigh_op_bot_1')
// (13, 8, 'sp4_v_b_23')
// (13, 9, 'sp4_h_l_47')
// (13, 9, 'sp4_v_b_10')
// (14, 6, 'neigh_op_tnl_1')
// (14, 7, 'neigh_op_lft_1')
// (14, 8, 'neigh_op_bnl_1')

wire n1168;
// (8, 11, 'neigh_op_tnr_3')
// (8, 12, 'neigh_op_rgt_3')
// (8, 13, 'neigh_op_bnr_3')
// (9, 11, 'neigh_op_top_3')
// (9, 12, 'lutff_3/out')
// (9, 13, 'neigh_op_bot_3')
// (10, 11, 'neigh_op_tnl_3')
// (10, 12, 'local_g1_3')
// (10, 12, 'lutff_6/in_0')
// (10, 12, 'neigh_op_lft_3')
// (10, 13, 'neigh_op_bnl_3')

reg n1169 = 0;
// (8, 11, 'neigh_op_tnr_4')
// (8, 12, 'neigh_op_rgt_4')
// (8, 13, 'neigh_op_bnr_4')
// (9, 11, 'local_g1_4')
// (9, 11, 'lutff_4/in_3')
// (9, 11, 'neigh_op_top_4')
// (9, 12, 'lutff_4/out')
// (9, 13, 'neigh_op_bot_4')
// (10, 11, 'neigh_op_tnl_4')
// (10, 12, 'neigh_op_lft_4')
// (10, 13, 'neigh_op_bnl_4')

wire n1170;
// (8, 11, 'neigh_op_tnr_5')
// (8, 12, 'neigh_op_rgt_5')
// (8, 13, 'neigh_op_bnr_5')
// (9, 11, 'local_g1_5')
// (9, 11, 'lutff_3/in_3')
// (9, 11, 'neigh_op_top_5')
// (9, 12, 'lutff_5/out')
// (9, 13, 'neigh_op_bot_5')
// (10, 11, 'neigh_op_tnl_5')
// (10, 12, 'neigh_op_lft_5')
// (10, 13, 'neigh_op_bnl_5')

reg n1171 = 0;
// (8, 11, 'sp4_h_r_2')
// (9, 11, 'sp4_h_r_15')
// (10, 11, 'local_g2_2')
// (10, 11, 'lutff_7/in_3')
// (10, 11, 'sp4_h_r_26')
// (11, 11, 'sp4_h_r_39')
// (11, 12, 'sp4_r_v_b_45')
// (11, 13, 'sp4_r_v_b_32')
// (11, 14, 'local_g3_5')
// (11, 14, 'lutff_7/in_1')
// (11, 14, 'sp4_r_v_b_21')
// (11, 14, 'sp4_r_v_b_45')
// (11, 15, 'sp4_r_v_b_32')
// (11, 15, 'sp4_r_v_b_8')
// (11, 16, 'neigh_op_tnr_4')
// (11, 16, 'sp4_r_v_b_21')
// (11, 16, 'sp4_r_v_b_37')
// (11, 17, 'neigh_op_rgt_4')
// (11, 17, 'sp4_r_v_b_24')
// (11, 17, 'sp4_r_v_b_8')
// (11, 18, 'neigh_op_bnr_4')
// (11, 18, 'sp4_r_v_b_13')
// (11, 19, 'sp4_r_v_b_0')
// (12, 11, 'sp4_h_l_39')
// (12, 11, 'sp4_v_t_45')
// (12, 12, 'sp4_v_b_45')
// (12, 13, 'sp4_v_b_32')
// (12, 13, 'sp4_v_t_45')
// (12, 14, 'sp4_v_b_21')
// (12, 14, 'sp4_v_b_45')
// (12, 15, 'sp4_v_b_32')
// (12, 15, 'sp4_v_b_8')
// (12, 15, 'sp4_v_t_37')
// (12, 16, 'neigh_op_top_4')
// (12, 16, 'sp4_v_b_21')
// (12, 16, 'sp4_v_b_37')
// (12, 17, 'local_g3_4')
// (12, 17, 'lutff_4/in_3')
// (12, 17, 'lutff_4/out')
// (12, 17, 'sp4_v_b_24')
// (12, 17, 'sp4_v_b_8')
// (12, 18, 'neigh_op_bot_4')
// (12, 18, 'sp4_v_b_13')
// (12, 19, 'sp4_v_b_0')
// (13, 16, 'neigh_op_tnl_4')
// (13, 17, 'neigh_op_lft_4')
// (13, 18, 'neigh_op_bnl_4')

reg n1172 = 0;
// (8, 12, 'neigh_op_tnr_0')
// (8, 13, 'local_g2_0')
// (8, 13, 'lutff_7/in_3')
// (8, 13, 'neigh_op_rgt_0')
// (8, 14, 'neigh_op_bnr_0')
// (9, 12, 'neigh_op_top_0')
// (9, 13, 'lutff_0/out')
// (9, 14, 'neigh_op_bot_0')
// (10, 12, 'neigh_op_tnl_0')
// (10, 13, 'neigh_op_lft_0')
// (10, 14, 'neigh_op_bnl_0')

reg n1173 = 0;
// (8, 12, 'neigh_op_tnr_1')
// (8, 13, 'local_g2_1')
// (8, 13, 'lutff_7/in_0')
// (8, 13, 'neigh_op_rgt_1')
// (8, 14, 'neigh_op_bnr_1')
// (9, 12, 'neigh_op_top_1')
// (9, 13, 'lutff_1/out')
// (9, 14, 'neigh_op_bot_1')
// (10, 12, 'neigh_op_tnl_1')
// (10, 13, 'neigh_op_lft_1')
// (10, 14, 'neigh_op_bnl_1')

reg n1174 = 0;
// (8, 12, 'neigh_op_tnr_2')
// (8, 13, 'neigh_op_rgt_2')
// (8, 14, 'neigh_op_bnr_2')
// (9, 12, 'local_g1_2')
// (9, 12, 'lutff_3/in_0')
// (9, 12, 'neigh_op_top_2')
// (9, 13, 'lutff_2/out')
// (9, 14, 'neigh_op_bot_2')
// (10, 12, 'neigh_op_tnl_2')
// (10, 13, 'neigh_op_lft_2')
// (10, 14, 'neigh_op_bnl_2')

wire n1175;
// (8, 12, 'neigh_op_tnr_3')
// (8, 13, 'neigh_op_rgt_3')
// (8, 14, 'neigh_op_bnr_3')
// (9, 12, 'neigh_op_top_3')
// (9, 13, 'local_g1_3')
// (9, 13, 'lutff_3/out')
// (9, 13, 'lutff_5/in_3')
// (9, 14, 'neigh_op_bot_3')
// (10, 12, 'neigh_op_tnl_3')
// (10, 13, 'neigh_op_lft_3')
// (10, 14, 'neigh_op_bnl_3')

reg n1176 = 0;
// (8, 12, 'neigh_op_tnr_4')
// (8, 13, 'neigh_op_rgt_4')
// (8, 14, 'neigh_op_bnr_4')
// (9, 12, 'local_g1_4')
// (9, 12, 'lutff_5/in_0')
// (9, 12, 'neigh_op_top_4')
// (9, 13, 'lutff_4/out')
// (9, 14, 'neigh_op_bot_4')
// (10, 12, 'neigh_op_tnl_4')
// (10, 13, 'neigh_op_lft_4')
// (10, 14, 'neigh_op_bnl_4')

reg n1177 = 0;
// (8, 12, 'neigh_op_tnr_6')
// (8, 13, 'neigh_op_rgt_6')
// (8, 14, 'neigh_op_bnr_6')
// (9, 12, 'local_g1_6')
// (9, 12, 'lutff_5/in_2')
// (9, 12, 'neigh_op_top_6')
// (9, 13, 'lutff_6/out')
// (9, 14, 'neigh_op_bot_6')
// (10, 12, 'neigh_op_tnl_6')
// (10, 13, 'neigh_op_lft_6')
// (10, 14, 'neigh_op_bnl_6')

reg n1178 = 0;
// (8, 12, 'neigh_op_tnr_7')
// (8, 13, 'neigh_op_rgt_7')
// (8, 14, 'neigh_op_bnr_7')
// (9, 12, 'local_g1_7')
// (9, 12, 'lutff_5/in_1')
// (9, 12, 'neigh_op_top_7')
// (9, 13, 'lutff_7/out')
// (9, 14, 'neigh_op_bot_7')
// (10, 12, 'neigh_op_tnl_7')
// (10, 13, 'neigh_op_lft_7')
// (10, 14, 'neigh_op_bnl_7')

wire n1179;
// (8, 12, 'sp4_h_r_0')
// (9, 12, 'local_g1_5')
// (9, 12, 'lutff_6/in_2')
// (9, 12, 'lutff_7/in_3')
// (9, 12, 'sp4_h_r_13')
// (10, 10, 'neigh_op_tnr_6')
// (10, 11, 'neigh_op_rgt_6')
// (10, 12, 'neigh_op_bnr_6')
// (10, 12, 'sp4_h_r_24')
// (11, 5, 'sp4_r_v_b_45')
// (11, 6, 'sp4_r_v_b_32')
// (11, 7, 'sp4_r_v_b_21')
// (11, 8, 'sp4_r_v_b_8')
// (11, 9, 'sp4_r_v_b_37')
// (11, 10, 'neigh_op_top_6')
// (11, 10, 'sp4_r_v_b_24')
// (11, 11, 'lutff_6/out')
// (11, 11, 'sp4_r_v_b_13')
// (11, 12, 'neigh_op_bot_6')
// (11, 12, 'sp4_h_r_37')
// (11, 12, 'sp4_r_v_b_0')
// (12, 4, 'sp4_h_r_8')
// (12, 4, 'sp4_v_t_45')
// (12, 5, 'sp4_v_b_45')
// (12, 6, 'sp4_v_b_32')
// (12, 7, 'sp4_v_b_21')
// (12, 8, 'sp4_v_b_8')
// (12, 8, 'sp4_v_t_37')
// (12, 9, 'sp4_v_b_37')
// (12, 10, 'neigh_op_tnl_6')
// (12, 10, 'sp4_v_b_24')
// (12, 11, 'neigh_op_lft_6')
// (12, 11, 'sp4_v_b_13')
// (12, 12, 'neigh_op_bnl_6')
// (12, 12, 'sp4_h_l_37')
// (12, 12, 'sp4_v_b_0')
// (13, 4, 'sp4_h_r_21')
// (14, 4, 'local_g3_0')
// (14, 4, 'lutff_5/in_2')
// (14, 4, 'sp4_h_r_32')
// (15, 1, 'sp4_r_v_b_45')
// (15, 2, 'sp4_r_v_b_32')
// (15, 3, 'local_g3_5')
// (15, 3, 'lutff_5/in_3')
// (15, 3, 'lutff_6/in_0')
// (15, 3, 'sp4_r_v_b_21')
// (15, 4, 'local_g3_5')
// (15, 4, 'lutff_0/in_2')
// (15, 4, 'sp4_h_r_45')
// (15, 4, 'sp4_r_v_b_8')
// (16, 0, 'span4_vert_45')
// (16, 1, 'sp4_v_b_45')
// (16, 2, 'sp4_v_b_32')
// (16, 3, 'sp4_v_b_21')
// (16, 4, 'sp4_h_l_45')
// (16, 4, 'sp4_v_b_8')

wire n1180;
// (8, 12, 'sp4_h_r_2')
// (9, 12, 'sp4_h_r_15')
// (9, 14, 'sp4_h_r_10')
// (10, 12, 'local_g2_2')
// (10, 12, 'lutff_global/cen')
// (10, 12, 'sp4_h_r_26')
// (10, 14, 'sp4_h_r_23')
// (11, 12, 'sp4_h_r_39')
// (11, 14, 'local_g2_2')
// (11, 14, 'lutff_global/cen')
// (11, 14, 'sp4_h_r_34')
// (11, 15, 'sp4_h_r_7')
// (12, 12, 'sp4_h_l_39')
// (12, 12, 'sp4_h_r_11')
// (12, 14, 'sp4_h_r_47')
// (12, 15, 'local_g0_2')
// (12, 15, 'lutff_global/cen')
// (12, 15, 'sp4_h_r_18')
// (13, 12, 'sp4_h_r_22')
// (13, 14, 'sp4_h_l_47')
// (13, 14, 'sp4_h_r_10')
// (13, 15, 'sp4_h_r_31')
// (14, 12, 'sp4_h_r_35')
// (14, 12, 'sp4_r_v_b_42')
// (14, 13, 'neigh_op_tnr_1')
// (14, 13, 'sp4_r_v_b_31')
// (14, 14, 'neigh_op_rgt_1')
// (14, 14, 'sp4_h_r_23')
// (14, 14, 'sp4_r_v_b_18')
// (14, 15, 'neigh_op_bnr_1')
// (14, 15, 'sp4_h_r_42')
// (14, 15, 'sp4_r_v_b_7')
// (15, 11, 'sp4_v_t_42')
// (15, 12, 'sp4_h_r_46')
// (15, 12, 'sp4_v_b_42')
// (15, 13, 'neigh_op_top_1')
// (15, 13, 'sp4_r_v_b_46')
// (15, 13, 'sp4_v_b_31')
// (15, 14, 'lutff_1/out')
// (15, 14, 'sp4_h_r_34')
// (15, 14, 'sp4_r_v_b_35')
// (15, 14, 'sp4_v_b_18')
// (15, 15, 'local_g0_2')
// (15, 15, 'lutff_global/cen')
// (15, 15, 'neigh_op_bot_1')
// (15, 15, 'sp4_h_l_42')
// (15, 15, 'sp4_h_r_10')
// (15, 15, 'sp4_r_v_b_22')
// (15, 15, 'sp4_v_b_7')
// (15, 16, 'sp4_r_v_b_11')
// (16, 12, 'sp4_h_l_46')
// (16, 12, 'sp4_v_t_46')
// (16, 13, 'neigh_op_tnl_1')
// (16, 13, 'sp4_v_b_46')
// (16, 14, 'neigh_op_lft_1')
// (16, 14, 'sp4_h_r_47')
// (16, 14, 'sp4_v_b_35')
// (16, 15, 'neigh_op_bnl_1')
// (16, 15, 'sp4_h_r_23')
// (16, 15, 'sp4_v_b_22')
// (16, 16, 'sp4_v_b_11')
// (17, 14, 'sp4_h_l_47')
// (17, 15, 'sp4_h_r_34')
// (18, 15, 'sp4_h_r_47')
// (19, 15, 'sp4_h_l_47')

wire n1181;
// (8, 12, 'sp4_h_r_5')
// (9, 12, 'sp4_h_r_16')
// (10, 12, 'local_g3_5')
// (10, 12, 'lutff_1/in_3')
// (10, 12, 'lutff_3/in_1')
// (10, 12, 'lutff_5/in_3')
// (10, 12, 'sp4_h_r_29')
// (11, 12, 'sp4_h_r_40')
// (11, 13, 'sp4_r_v_b_46')
// (11, 14, 'local_g3_3')
// (11, 14, 'lutff_1/in_3')
// (11, 14, 'lutff_4/in_0')
// (11, 14, 'neigh_op_tnr_3')
// (11, 14, 'sp4_r_v_b_35')
// (11, 15, 'neigh_op_rgt_3')
// (11, 15, 'sp4_r_v_b_22')
// (11, 16, 'neigh_op_bnr_3')
// (11, 16, 'sp4_r_v_b_11')
// (12, 12, 'sp4_h_l_40')
// (12, 12, 'sp4_v_t_46')
// (12, 13, 'sp4_v_b_46')
// (12, 14, 'neigh_op_top_3')
// (12, 14, 'sp4_v_b_35')
// (12, 15, 'local_g3_3')
// (12, 15, 'lutff_0/in_0')
// (12, 15, 'lutff_1/in_1')
// (12, 15, 'lutff_3/out')
// (12, 15, 'lutff_6/in_2')
// (12, 15, 'lutff_7/in_3')
// (12, 15, 'sp4_v_b_22')
// (12, 16, 'neigh_op_bot_3')
// (12, 16, 'sp4_v_b_11')
// (13, 14, 'neigh_op_tnl_3')
// (13, 15, 'neigh_op_lft_3')
// (13, 16, 'neigh_op_bnl_3')

reg n1182 = 0;
// (8, 12, 'sp4_h_r_9')
// (9, 12, 'sp4_h_r_20')
// (10, 12, 'local_g2_1')
// (10, 12, 'lutff_3/in_0')
// (10, 12, 'sp4_h_r_33')
// (11, 12, 'neigh_op_tnr_6')
// (11, 12, 'sp4_h_r_44')
// (11, 13, 'neigh_op_rgt_6')
// (11, 13, 'sp4_r_v_b_44')
// (11, 14, 'neigh_op_bnr_6')
// (11, 14, 'sp4_r_v_b_33')
// (11, 15, 'sp4_r_v_b_20')
// (11, 16, 'sp4_r_v_b_9')
// (12, 12, 'neigh_op_top_6')
// (12, 12, 'sp4_h_l_44')
// (12, 12, 'sp4_v_t_44')
// (12, 13, 'lutff_6/out')
// (12, 13, 'sp4_v_b_44')
// (12, 14, 'neigh_op_bot_6')
// (12, 14, 'sp4_v_b_33')
// (12, 15, 'sp4_v_b_20')
// (12, 16, 'sp4_v_b_9')
// (13, 12, 'neigh_op_tnl_6')
// (13, 13, 'neigh_op_lft_6')
// (13, 14, 'neigh_op_bnl_6')

wire n1183;
// (8, 13, 'neigh_op_tnr_1')
// (8, 14, 'neigh_op_rgt_1')
// (8, 15, 'neigh_op_bnr_1')
// (9, 13, 'neigh_op_top_1')
// (9, 14, 'lutff_1/out')
// (9, 15, 'neigh_op_bot_1')
// (10, 13, 'neigh_op_tnl_1')
// (10, 14, 'local_g1_1')
// (10, 14, 'lutff_2/in_0')
// (10, 14, 'neigh_op_lft_1')
// (10, 15, 'neigh_op_bnl_1')

reg n1184 = 0;
// (8, 13, 'neigh_op_tnr_3')
// (8, 14, 'neigh_op_rgt_3')
// (8, 15, 'neigh_op_bnr_3')
// (9, 13, 'neigh_op_top_3')
// (9, 14, 'lutff_3/out')
// (9, 14, 'sp4_r_v_b_39')
// (9, 15, 'local_g1_3')
// (9, 15, 'lutff_3/in_1')
// (9, 15, 'neigh_op_bot_3')
// (9, 15, 'sp4_r_v_b_26')
// (9, 16, 'sp4_r_v_b_15')
// (9, 17, 'sp4_r_v_b_2')
// (10, 13, 'neigh_op_tnl_3')
// (10, 13, 'sp4_v_t_39')
// (10, 14, 'neigh_op_lft_3')
// (10, 14, 'sp4_v_b_39')
// (10, 15, 'neigh_op_bnl_3')
// (10, 15, 'sp4_v_b_26')
// (10, 16, 'local_g0_7')
// (10, 16, 'lutff_6/in_3')
// (10, 16, 'sp4_v_b_15')
// (10, 17, 'sp4_v_b_2')

reg n1185 = 0;
// (8, 13, 'neigh_op_tnr_5')
// (8, 14, 'neigh_op_rgt_5')
// (8, 15, 'neigh_op_bnr_5')
// (9, 11, 'local_g3_6')
// (9, 11, 'lutff_7/in_2')
// (9, 11, 'sp4_r_v_b_46')
// (9, 12, 'sp4_r_v_b_35')
// (9, 13, 'neigh_op_top_5')
// (9, 13, 'sp4_r_v_b_22')
// (9, 14, 'lutff_5/out')
// (9, 14, 'sp4_r_v_b_11')
// (9, 15, 'neigh_op_bot_5')
// (10, 10, 'sp4_v_t_46')
// (10, 11, 'sp4_v_b_46')
// (10, 12, 'sp4_v_b_35')
// (10, 13, 'neigh_op_tnl_5')
// (10, 13, 'sp4_v_b_22')
// (10, 14, 'neigh_op_lft_5')
// (10, 14, 'sp4_v_b_11')
// (10, 15, 'neigh_op_bnl_5')

reg n1186 = 0;
// (8, 13, 'neigh_op_tnr_7')
// (8, 14, 'neigh_op_rgt_7')
// (8, 15, 'neigh_op_bnr_7')
// (9, 13, 'neigh_op_top_7')
// (9, 14, 'lutff_7/out')
// (9, 15, 'neigh_op_bot_7')
// (10, 13, 'local_g3_7')
// (10, 13, 'lutff_7/in_3')
// (10, 13, 'neigh_op_tnl_7')
// (10, 14, 'neigh_op_lft_7')
// (10, 15, 'local_g2_7')
// (10, 15, 'lutff_4/in_1')
// (10, 15, 'neigh_op_bnl_7')

wire n1187;
// (8, 13, 'sp4_h_r_3')
// (9, 13, 'local_g0_6')
// (9, 13, 'lutff_5/in_1')
// (9, 13, 'sp4_h_r_14')
// (10, 6, 'neigh_op_tnr_7')
// (10, 7, 'neigh_op_rgt_7')
// (10, 8, 'neigh_op_bnr_7')
// (10, 13, 'sp4_h_r_27')
// (11, 6, 'neigh_op_top_7')
// (11, 6, 'sp4_r_v_b_42')
// (11, 7, 'lutff_7/out')
// (11, 7, 'sp4_r_v_b_31')
// (11, 8, 'neigh_op_bot_7')
// (11, 8, 'sp4_r_v_b_18')
// (11, 9, 'sp4_r_v_b_7')
// (11, 10, 'sp4_r_v_b_47')
// (11, 11, 'sp4_r_v_b_34')
// (11, 12, 'sp4_r_v_b_23')
// (11, 13, 'sp4_h_r_38')
// (11, 13, 'sp4_r_v_b_10')
// (12, 5, 'sp4_v_t_42')
// (12, 6, 'neigh_op_tnl_7')
// (12, 6, 'sp4_v_b_42')
// (12, 7, 'neigh_op_lft_7')
// (12, 7, 'sp4_v_b_31')
// (12, 8, 'neigh_op_bnl_7')
// (12, 8, 'sp4_v_b_18')
// (12, 9, 'sp4_v_b_7')
// (12, 9, 'sp4_v_t_47')
// (12, 10, 'sp4_v_b_47')
// (12, 11, 'sp4_v_b_34')
// (12, 12, 'sp4_v_b_23')
// (12, 13, 'sp4_h_l_38')
// (12, 13, 'sp4_v_b_10')

reg n1188 = 0;
// (8, 13, 'sp4_h_r_9')
// (9, 13, 'sp4_h_r_20')
// (10, 13, 'local_g3_1')
// (10, 13, 'lutff_3/in_1')
// (10, 13, 'sp4_h_r_33')
// (11, 13, 'sp4_h_r_44')
// (11, 14, 'sp4_r_v_b_44')
// (11, 15, 'sp4_r_v_b_33')
// (11, 16, 'sp4_r_v_b_20')
// (11, 17, 'neigh_op_tnr_2')
// (11, 17, 'sp4_r_v_b_9')
// (11, 18, 'neigh_op_rgt_2')
// (11, 18, 'sp4_r_v_b_36')
// (11, 19, 'neigh_op_bnr_2')
// (11, 19, 'sp4_r_v_b_25')
// (11, 20, 'sp4_r_v_b_12')
// (11, 21, 'sp4_r_v_b_1')
// (12, 13, 'sp4_h_l_44')
// (12, 13, 'sp4_v_t_44')
// (12, 14, 'sp4_v_b_44')
// (12, 15, 'sp4_v_b_33')
// (12, 16, 'sp4_v_b_20')
// (12, 17, 'neigh_op_top_2')
// (12, 17, 'sp4_v_b_9')
// (12, 17, 'sp4_v_t_36')
// (12, 18, 'local_g2_2')
// (12, 18, 'lutff_2/in_2')
// (12, 18, 'lutff_2/out')
// (12, 18, 'sp4_v_b_36')
// (12, 19, 'neigh_op_bot_2')
// (12, 19, 'sp4_v_b_25')
// (12, 20, 'sp4_v_b_12')
// (12, 21, 'sp4_v_b_1')
// (13, 17, 'neigh_op_tnl_2')
// (13, 18, 'neigh_op_lft_2')
// (13, 19, 'neigh_op_bnl_2')

reg n1189 = 0;
// (8, 14, 'local_g2_7')
// (8, 14, 'lutff_5/in_0')
// (8, 14, 'sp4_r_v_b_39')
// (8, 15, 'sp4_r_v_b_26')
// (8, 16, 'sp4_r_v_b_15')
// (8, 17, 'sp4_r_v_b_2')
// (8, 18, 'sp4_r_v_b_39')
// (8, 19, 'sp4_r_v_b_26')
// (8, 20, 'neigh_op_tnr_1')
// (8, 20, 'sp4_r_v_b_15')
// (8, 21, 'neigh_op_rgt_1')
// (8, 21, 'sp4_r_v_b_2')
// (8, 22, 'neigh_op_bnr_1')
// (9, 0, 'span12_vert_18')
// (9, 1, 'sp12_v_b_18')
// (9, 2, 'sp12_v_b_17')
// (9, 3, 'sp12_v_b_14')
// (9, 4, 'sp12_v_b_13')
// (9, 5, 'sp12_v_b_10')
// (9, 6, 'sp12_v_b_9')
// (9, 7, 'sp12_v_b_6')
// (9, 8, 'local_g2_5')
// (9, 8, 'lutff_7/in_2')
// (9, 8, 'sp12_v_b_5')
// (9, 9, 'sp12_v_b_2')
// (9, 10, 'sp12_v_b_1')
// (9, 10, 'sp12_v_t_22')
// (9, 11, 'sp12_v_b_22')
// (9, 12, 'sp12_v_b_21')
// (9, 13, 'sp12_v_b_18')
// (9, 13, 'sp4_v_t_39')
// (9, 14, 'sp12_v_b_17')
// (9, 14, 'sp4_v_b_39')
// (9, 15, 'sp12_v_b_14')
// (9, 15, 'sp4_v_b_26')
// (9, 16, 'sp12_v_b_13')
// (9, 16, 'sp4_v_b_15')
// (9, 17, 'sp12_v_b_10')
// (9, 17, 'sp4_v_b_2')
// (9, 17, 'sp4_v_t_39')
// (9, 18, 'sp12_v_b_9')
// (9, 18, 'sp4_v_b_39')
// (9, 19, 'local_g2_2')
// (9, 19, 'lutff_5/in_3')
// (9, 19, 'lutff_7/in_3')
// (9, 19, 'sp12_v_b_6')
// (9, 19, 'sp4_r_v_b_43')
// (9, 19, 'sp4_v_b_26')
// (9, 20, 'local_g1_1')
// (9, 20, 'lutff_5/in_1')
// (9, 20, 'neigh_op_top_1')
// (9, 20, 'sp12_v_b_5')
// (9, 20, 'sp4_r_v_b_30')
// (9, 20, 'sp4_v_b_15')
// (9, 21, 'lutff_1/out')
// (9, 21, 'sp12_v_b_2')
// (9, 21, 'sp4_r_v_b_19')
// (9, 21, 'sp4_v_b_2')
// (9, 22, 'local_g1_1')
// (9, 22, 'lutff_2/in_2')
// (9, 22, 'neigh_op_bot_1')
// (9, 22, 'sp12_v_b_1')
// (9, 22, 'sp4_r_v_b_6')
// (10, 18, 'sp4_v_t_43')
// (10, 19, 'local_g3_3')
// (10, 19, 'lutff_7/in_3')
// (10, 19, 'sp4_v_b_43')
// (10, 20, 'local_g2_1')
// (10, 20, 'lutff_7/in_2')
// (10, 20, 'neigh_op_tnl_1')
// (10, 20, 'sp4_v_b_30')
// (10, 21, 'neigh_op_lft_1')
// (10, 21, 'sp4_v_b_19')
// (10, 22, 'neigh_op_bnl_1')
// (10, 22, 'sp4_v_b_6')

wire n1190;
// (8, 14, 'neigh_op_tnr_0')
// (8, 15, 'neigh_op_rgt_0')
// (8, 16, 'neigh_op_bnr_0')
// (9, 14, 'neigh_op_top_0')
// (9, 14, 'sp4_r_v_b_44')
// (9, 15, 'lutff_0/out')
// (9, 15, 'sp4_r_v_b_33')
// (9, 16, 'neigh_op_bot_0')
// (9, 16, 'sp4_r_v_b_20')
// (9, 17, 'local_g2_1')
// (9, 17, 'lutff_3/in_2')
// (9, 17, 'sp4_r_v_b_9')
// (10, 13, 'sp4_v_t_44')
// (10, 14, 'neigh_op_tnl_0')
// (10, 14, 'sp4_v_b_44')
// (10, 15, 'neigh_op_lft_0')
// (10, 15, 'sp4_v_b_33')
// (10, 16, 'neigh_op_bnl_0')
// (10, 16, 'sp4_v_b_20')
// (10, 17, 'sp4_v_b_9')

wire n1191;
// (8, 14, 'neigh_op_tnr_2')
// (8, 15, 'neigh_op_rgt_2')
// (8, 16, 'neigh_op_bnr_2')
// (9, 14, 'neigh_op_top_2')
// (9, 15, 'lutff_2/out')
// (9, 16, 'neigh_op_bot_2')
// (10, 14, 'neigh_op_tnl_2')
// (10, 15, 'local_g1_2')
// (10, 15, 'lutff_3/in_0')
// (10, 15, 'neigh_op_lft_2')
// (10, 16, 'neigh_op_bnl_2')

reg n1192 = 0;
// (8, 14, 'neigh_op_tnr_3')
// (8, 15, 'neigh_op_rgt_3')
// (8, 16, 'neigh_op_bnr_3')
// (9, 14, 'local_g0_3')
// (9, 14, 'lutff_1/in_0')
// (9, 14, 'neigh_op_top_3')
// (9, 15, 'lutff_3/out')
// (9, 16, 'neigh_op_bot_3')
// (10, 14, 'neigh_op_tnl_3')
// (10, 15, 'neigh_op_lft_3')
// (10, 16, 'neigh_op_bnl_3')

wire n1193;
// (8, 14, 'neigh_op_tnr_4')
// (8, 15, 'neigh_op_rgt_4')
// (8, 16, 'neigh_op_bnr_4')
// (9, 14, 'neigh_op_top_4')
// (9, 15, 'local_g3_4')
// (9, 15, 'lutff_0/in_3')
// (9, 15, 'lutff_4/out')
// (9, 16, 'neigh_op_bot_4')
// (10, 14, 'neigh_op_tnl_4')
// (10, 15, 'neigh_op_lft_4')
// (10, 16, 'neigh_op_bnl_4')

reg n1194 = 0;
// (8, 14, 'neigh_op_tnr_5')
// (8, 15, 'neigh_op_rgt_5')
// (8, 16, 'neigh_op_bnr_5')
// (9, 14, 'neigh_op_top_5')
// (9, 15, 'local_g2_5')
// (9, 15, 'lutff_2/in_1')
// (9, 15, 'lutff_5/out')
// (9, 16, 'neigh_op_bot_5')
// (10, 14, 'neigh_op_tnl_5')
// (10, 15, 'neigh_op_lft_5')
// (10, 16, 'neigh_op_bnl_5')

wire n1195;
// (8, 14, 'neigh_op_tnr_6')
// (8, 15, 'neigh_op_rgt_6')
// (8, 15, 'sp4_h_r_1')
// (8, 16, 'neigh_op_bnr_6')
// (9, 14, 'neigh_op_top_6')
// (9, 15, 'lutff_6/out')
// (9, 15, 'sp4_h_r_12')
// (9, 16, 'neigh_op_bot_6')
// (10, 14, 'neigh_op_tnl_6')
// (10, 15, 'neigh_op_lft_6')
// (10, 15, 'sp4_h_r_25')
// (10, 16, 'neigh_op_bnl_6')
// (11, 15, 'local_g3_4')
// (11, 15, 'lutff_6/in_3')
// (11, 15, 'sp4_h_r_36')
// (12, 15, 'sp4_h_l_36')

wire n1196;
// (8, 14, 'neigh_op_tnr_7')
// (8, 15, 'neigh_op_rgt_7')
// (8, 16, 'neigh_op_bnr_7')
// (9, 14, 'neigh_op_top_7')
// (9, 15, 'local_g1_7')
// (9, 15, 'lutff_0/in_2')
// (9, 15, 'lutff_7/out')
// (9, 16, 'neigh_op_bot_7')
// (10, 14, 'neigh_op_tnl_7')
// (10, 15, 'neigh_op_lft_7')
// (10, 16, 'neigh_op_bnl_7')

wire n1197;
// (8, 15, 'lutff_7/cout')
// (8, 16, 'carry_in')
// (8, 16, 'carry_in_mux')

wire n1198;
// (8, 16, 'lutff_0/cout')
// (8, 16, 'lutff_1/in_3')

wire n1199;
// (8, 16, 'neigh_op_tnr_1')
// (8, 17, 'neigh_op_rgt_1')
// (8, 18, 'local_g1_1')
// (8, 18, 'lutff_1/in_1')
// (8, 18, 'neigh_op_bnr_1')
// (9, 16, 'neigh_op_top_1')
// (9, 17, 'lutff_1/out')
// (9, 18, 'neigh_op_bot_1')
// (10, 16, 'neigh_op_tnl_1')
// (10, 17, 'neigh_op_lft_1')
// (10, 18, 'neigh_op_bnl_1')

reg n1200 = 0;
// (8, 16, 'neigh_op_tnr_2')
// (8, 17, 'neigh_op_rgt_2')
// (8, 18, 'neigh_op_bnr_2')
// (9, 16, 'neigh_op_top_2')
// (9, 17, 'local_g3_2')
// (9, 17, 'lutff_2/out')
// (9, 17, 'lutff_5/in_0')
// (9, 18, 'neigh_op_bot_2')
// (10, 16, 'neigh_op_tnl_2')
// (10, 17, 'neigh_op_lft_2')
// (10, 18, 'neigh_op_bnl_2')

wire n1201;
// (8, 16, 'neigh_op_tnr_3')
// (8, 17, 'neigh_op_rgt_3')
// (8, 18, 'neigh_op_bnr_3')
// (9, 16, 'neigh_op_top_3')
// (9, 17, 'local_g1_3')
// (9, 17, 'lutff_2/in_2')
// (9, 17, 'lutff_3/out')
// (9, 17, 'lutff_5/in_1')
// (9, 18, 'neigh_op_bot_3')
// (10, 16, 'local_g2_3')
// (10, 16, 'lutff_4/in_3')
// (10, 16, 'neigh_op_tnl_3')
// (10, 17, 'neigh_op_lft_3')
// (10, 18, 'neigh_op_bnl_3')

reg n1202 = 0;
// (8, 16, 'neigh_op_tnr_4')
// (8, 17, 'neigh_op_rgt_4')
// (8, 18, 'neigh_op_bnr_4')
// (9, 16, 'neigh_op_top_4')
// (9, 17, 'local_g3_4')
// (9, 17, 'lutff_4/out')
// (9, 17, 'lutff_5/in_2')
// (9, 18, 'neigh_op_bot_4')
// (10, 16, 'neigh_op_tnl_4')
// (10, 17, 'neigh_op_lft_4')
// (10, 18, 'neigh_op_bnl_4')

wire n1203;
// (8, 16, 'neigh_op_tnr_5')
// (8, 17, 'neigh_op_rgt_5')
// (8, 18, 'neigh_op_bnr_5')
// (9, 16, 'neigh_op_top_5')
// (9, 17, 'lutff_5/out')
// (9, 18, 'neigh_op_bot_5')
// (10, 16, 'local_g3_5')
// (10, 16, 'lutff_6/in_2')
// (10, 16, 'neigh_op_tnl_5')
// (10, 17, 'neigh_op_lft_5')
// (10, 18, 'neigh_op_bnl_5')

wire n1204;
// (8, 16, 'sp12_h_r_1')
// (9, 16, 'sp12_h_r_2')
// (10, 16, 'sp12_h_r_5')
// (11, 16, 'sp12_h_r_6')
// (12, 16, 'local_g0_1')
// (12, 16, 'lutff_1/in_2')
// (12, 16, 'sp12_h_r_9')
// (13, 16, 'sp12_h_r_10')
// (14, 16, 'sp12_h_r_13')
// (15, 16, 'sp12_h_r_14')
// (16, 16, 'sp12_h_r_17')
// (17, 16, 'sp12_h_r_18')
// (18, 15, 'neigh_op_tnr_7')
// (18, 16, 'neigh_op_rgt_7')
// (18, 16, 'sp12_h_r_21')
// (18, 17, 'neigh_op_bnr_7')
// (19, 15, 'neigh_op_top_7')
// (19, 16, 'ram/RDATA_0')
// (19, 16, 'sp12_h_r_22')
// (19, 17, 'neigh_op_bot_7')
// (20, 15, 'neigh_op_tnl_7')
// (20, 16, 'neigh_op_lft_7')
// (20, 16, 'sp12_h_l_22')
// (20, 17, 'neigh_op_bnl_7')

wire n1205;
// (8, 17, 'lutff_7/cout')
// (8, 18, 'carry_in')
// (8, 18, 'carry_in_mux')

wire n1206;
// (8, 17, 'sp4_r_v_b_41')
// (8, 18, 'sp4_r_v_b_28')
// (8, 19, 'neigh_op_tnr_2')
// (8, 19, 'sp4_r_v_b_17')
// (8, 20, 'local_g1_4')
// (8, 20, 'lutff_2/in_1')
// (8, 20, 'neigh_op_rgt_2')
// (8, 20, 'sp4_r_v_b_4')
// (8, 21, 'neigh_op_bnr_2')
// (9, 16, 'sp4_v_t_41')
// (9, 17, 'sp4_v_b_41')
// (9, 18, 'sp4_v_b_28')
// (9, 19, 'neigh_op_top_2')
// (9, 19, 'sp4_v_b_17')
// (9, 20, 'lutff_2/out')
// (9, 20, 'sp4_v_b_4')
// (9, 21, 'neigh_op_bot_2')
// (10, 19, 'neigh_op_tnl_2')
// (10, 20, 'neigh_op_lft_2')
// (10, 21, 'neigh_op_bnl_2')

wire n1207;
// (8, 18, 'local_g3_4')
// (8, 18, 'lutff_5/in_0')
// (8, 18, 'neigh_op_tnr_4')
// (8, 19, 'neigh_op_rgt_4')
// (8, 20, 'neigh_op_bnr_4')
// (9, 18, 'neigh_op_top_4')
// (9, 19, 'lutff_4/out')
// (9, 20, 'neigh_op_bot_4')
// (10, 18, 'neigh_op_tnl_4')
// (10, 19, 'neigh_op_lft_4')
// (10, 20, 'neigh_op_bnl_4')

wire n1208;
// (8, 18, 'lutff_0/cout')
// (8, 18, 'lutff_1/in_3')

wire n1209;
// (8, 18, 'neigh_op_tnr_2')
// (8, 19, 'neigh_op_rgt_2')
// (8, 20, 'neigh_op_bnr_2')
// (9, 18, 'neigh_op_top_2')
// (9, 19, 'local_g0_2')
// (9, 19, 'lutff_2/out')
// (9, 19, 'lutff_5/in_1')
// (9, 20, 'neigh_op_bot_2')
// (10, 18, 'neigh_op_tnl_2')
// (10, 19, 'neigh_op_lft_2')
// (10, 20, 'neigh_op_bnl_2')

wire n1210;
// (8, 18, 'neigh_op_tnr_3')
// (8, 19, 'neigh_op_rgt_3')
// (8, 20, 'neigh_op_bnr_3')
// (9, 18, 'neigh_op_top_3')
// (9, 19, 'local_g0_3')
// (9, 19, 'lutff_3/out')
// (9, 19, 'lutff_4/in_1')
// (9, 19, 'lutff_5/in_2')
// (9, 20, 'neigh_op_bot_3')
// (10, 18, 'neigh_op_tnl_3')
// (10, 19, 'local_g0_3')
// (10, 19, 'lutff_5/in_2')
// (10, 19, 'neigh_op_lft_3')
// (10, 20, 'neigh_op_bnl_3')

wire n1211;
// (8, 18, 'neigh_op_tnr_5')
// (8, 19, 'neigh_op_rgt_5')
// (8, 20, 'local_g0_5')
// (8, 20, 'lutff_1/in_0')
// (8, 20, 'neigh_op_bnr_5')
// (9, 18, 'neigh_op_top_5')
// (9, 19, 'lutff_5/out')
// (9, 20, 'neigh_op_bot_5')
// (10, 18, 'neigh_op_tnl_5')
// (10, 19, 'neigh_op_lft_5')
// (10, 20, 'neigh_op_bnl_5')

wire n1212;
// (8, 18, 'neigh_op_tnr_6')
// (8, 19, 'neigh_op_rgt_6')
// (8, 20, 'neigh_op_bnr_6')
// (9, 18, 'neigh_op_top_6')
// (9, 19, 'local_g0_6')
// (9, 19, 'lutff_1/in_1')
// (9, 19, 'lutff_6/out')
// (9, 20, 'neigh_op_bot_6')
// (10, 18, 'neigh_op_tnl_6')
// (10, 19, 'neigh_op_lft_6')
// (10, 20, 'neigh_op_bnl_6')

wire n1213;
// (8, 18, 'neigh_op_tnr_7')
// (8, 19, 'neigh_op_rgt_7')
// (8, 20, 'neigh_op_bnr_7')
// (9, 18, 'neigh_op_top_7')
// (9, 19, 'local_g1_7')
// (9, 19, 'lutff_4/in_2')
// (9, 19, 'lutff_7/out')
// (9, 20, 'neigh_op_bot_7')
// (10, 18, 'neigh_op_tnl_7')
// (10, 19, 'neigh_op_lft_7')
// (10, 20, 'neigh_op_bnl_7')

wire n1214;
// (8, 19, 'lutff_7/cout')
// (8, 20, 'carry_in')
// (8, 20, 'carry_in_mux')

wire n1215;
// (8, 19, 'neigh_op_tnr_3')
// (8, 20, 'neigh_op_rgt_3')
// (8, 21, 'local_g0_3')
// (8, 21, 'lutff_2/in_3')
// (8, 21, 'neigh_op_bnr_3')
// (9, 19, 'neigh_op_top_3')
// (9, 20, 'lutff_3/out')
// (9, 21, 'neigh_op_bot_3')
// (10, 19, 'neigh_op_tnl_3')
// (10, 20, 'neigh_op_lft_3')
// (10, 21, 'neigh_op_bnl_3')

wire n1216;
// (8, 19, 'neigh_op_tnr_4')
// (8, 20, 'neigh_op_rgt_4')
// (8, 21, 'local_g0_4')
// (8, 21, 'lutff_0/in_2')
// (8, 21, 'neigh_op_bnr_4')
// (9, 19, 'neigh_op_top_4')
// (9, 20, 'lutff_4/out')
// (9, 21, 'neigh_op_bot_4')
// (10, 19, 'neigh_op_tnl_4')
// (10, 20, 'neigh_op_lft_4')
// (10, 21, 'neigh_op_bnl_4')

wire n1217;
// (8, 19, 'neigh_op_tnr_5')
// (8, 20, 'neigh_op_rgt_5')
// (8, 21, 'neigh_op_bnr_5')
// (9, 19, 'neigh_op_top_5')
// (9, 20, 'lutff_5/out')
// (9, 21, 'local_g1_5')
// (9, 21, 'lutff_3/in_1')
// (9, 21, 'neigh_op_bot_5')
// (10, 19, 'neigh_op_tnl_5')
// (10, 20, 'neigh_op_lft_5')
// (10, 21, 'neigh_op_bnl_5')

wire n1218;
// (8, 19, 'neigh_op_tnr_6')
// (8, 20, 'neigh_op_rgt_6')
// (8, 21, 'neigh_op_bnr_6')
// (9, 19, 'neigh_op_top_6')
// (9, 20, 'lutff_6/out')
// (9, 21, 'local_g1_6')
// (9, 21, 'lutff_2/in_3')
// (9, 21, 'neigh_op_bot_6')
// (10, 19, 'neigh_op_tnl_6')
// (10, 20, 'neigh_op_lft_6')
// (10, 21, 'neigh_op_bnl_6')

wire n1219;
// (8, 19, 'neigh_op_tnr_7')
// (8, 20, 'neigh_op_rgt_7')
// (8, 21, 'neigh_op_bnr_7')
// (9, 19, 'neigh_op_top_7')
// (9, 20, 'lutff_7/out')
// (9, 21, 'local_g0_7')
// (9, 21, 'lutff_6/in_1')
// (9, 21, 'neigh_op_bot_7')
// (10, 19, 'neigh_op_tnl_7')
// (10, 20, 'neigh_op_lft_7')
// (10, 21, 'neigh_op_bnl_7')

wire n1220;
// (8, 20, 'lutff_0/cout')
// (8, 20, 'lutff_1/in_3')

wire n1221;
// (8, 20, 'neigh_op_tnr_0')
// (8, 21, 'local_g3_0')
// (8, 21, 'lutff_6/in_3')
// (8, 21, 'neigh_op_rgt_0')
// (8, 22, 'neigh_op_bnr_0')
// (9, 20, 'neigh_op_top_0')
// (9, 21, 'lutff_0/out')
// (9, 22, 'neigh_op_bot_0')
// (10, 20, 'neigh_op_tnl_0')
// (10, 21, 'neigh_op_lft_0')
// (10, 22, 'neigh_op_bnl_0')

wire n1222;
// (8, 20, 'neigh_op_tnr_2')
// (8, 21, 'local_g3_2')
// (8, 21, 'lutff_1/in_0')
// (8, 21, 'neigh_op_rgt_2')
// (8, 22, 'neigh_op_bnr_2')
// (9, 20, 'neigh_op_top_2')
// (9, 21, 'lutff_2/out')
// (9, 22, 'neigh_op_bot_2')
// (10, 20, 'neigh_op_tnl_2')
// (10, 21, 'neigh_op_lft_2')
// (10, 22, 'neigh_op_bnl_2')

wire n1223;
// (8, 20, 'neigh_op_tnr_3')
// (8, 21, 'neigh_op_rgt_3')
// (8, 22, 'neigh_op_bnr_3')
// (9, 20, 'neigh_op_top_3')
// (9, 21, 'local_g0_3')
// (9, 21, 'lutff_1/in_2')
// (9, 21, 'lutff_3/out')
// (9, 22, 'neigh_op_bot_3')
// (10, 20, 'neigh_op_tnl_3')
// (10, 21, 'neigh_op_lft_3')
// (10, 22, 'neigh_op_bnl_3')

wire n1224;
// (8, 20, 'neigh_op_tnr_5')
// (8, 21, 'neigh_op_rgt_5')
// (8, 22, 'neigh_op_bnr_5')
// (9, 20, 'neigh_op_top_5')
// (9, 21, 'local_g0_5')
// (9, 21, 'lutff_4/in_1')
// (9, 21, 'lutff_5/out')
// (9, 22, 'neigh_op_bot_5')
// (10, 20, 'neigh_op_tnl_5')
// (10, 21, 'neigh_op_lft_5')
// (10, 22, 'neigh_op_bnl_5')

wire n1225;
// (8, 20, 'neigh_op_tnr_6')
// (8, 21, 'neigh_op_rgt_6')
// (8, 22, 'neigh_op_bnr_6')
// (9, 20, 'neigh_op_top_6')
// (9, 21, 'local_g2_6')
// (9, 21, 'lutff_4/in_2')
// (9, 21, 'lutff_6/out')
// (9, 22, 'neigh_op_bot_6')
// (10, 20, 'neigh_op_tnl_6')
// (10, 21, 'neigh_op_lft_6')
// (10, 22, 'neigh_op_bnl_6')

wire n1226;
// (8, 20, 'neigh_op_tnr_7')
// (8, 21, 'neigh_op_rgt_7')
// (8, 22, 'neigh_op_bnr_7')
// (9, 20, 'neigh_op_top_7')
// (9, 21, 'local_g3_7')
// (9, 21, 'lutff_1/in_1')
// (9, 21, 'lutff_7/out')
// (9, 22, 'neigh_op_bot_7')
// (10, 20, 'neigh_op_tnl_7')
// (10, 21, 'neigh_op_lft_7')
// (10, 22, 'neigh_op_bnl_7')

wire n1227;
// (8, 21, 'local_g3_5')
// (8, 21, 'lutff_6/in_2')
// (8, 21, 'neigh_op_tnr_5')
// (8, 22, 'neigh_op_rgt_5')
// (8, 23, 'neigh_op_bnr_5')
// (9, 21, 'neigh_op_top_5')
// (9, 22, 'lutff_5/out')
// (9, 23, 'neigh_op_bot_5')
// (10, 21, 'neigh_op_tnl_5')
// (10, 22, 'neigh_op_lft_5')
// (10, 23, 'neigh_op_bnl_5')

wire n1228;
// (8, 21, 'neigh_op_tnr_1')
// (8, 22, 'local_g3_1')
// (8, 22, 'lutff_0/in_0')
// (8, 22, 'neigh_op_rgt_1')
// (8, 23, 'neigh_op_bnr_1')
// (9, 21, 'neigh_op_top_1')
// (9, 22, 'lutff_1/out')
// (9, 23, 'neigh_op_bot_1')
// (10, 21, 'neigh_op_tnl_1')
// (10, 22, 'neigh_op_lft_1')
// (10, 23, 'neigh_op_bnl_1')

wire n1229;
// (8, 21, 'neigh_op_tnr_2')
// (8, 22, 'neigh_op_rgt_2')
// (8, 23, 'neigh_op_bnr_2')
// (9, 21, 'neigh_op_top_2')
// (9, 22, 'local_g1_2')
// (9, 22, 'lutff_2/out')
// (9, 22, 'lutff_7/in_2')
// (9, 23, 'neigh_op_bot_2')
// (10, 21, 'neigh_op_tnl_2')
// (10, 22, 'neigh_op_lft_2')
// (10, 23, 'neigh_op_bnl_2')

wire n1230;
// (8, 21, 'neigh_op_tnr_3')
// (8, 22, 'local_g3_3')
// (8, 22, 'lutff_7/in_1')
// (8, 22, 'neigh_op_rgt_3')
// (8, 23, 'neigh_op_bnr_3')
// (9, 21, 'neigh_op_top_3')
// (9, 22, 'lutff_3/out')
// (9, 23, 'neigh_op_bot_3')
// (10, 21, 'neigh_op_tnl_3')
// (10, 22, 'neigh_op_lft_3')
// (10, 23, 'neigh_op_bnl_3')

wire n1231;
// (8, 21, 'neigh_op_tnr_4')
// (8, 22, 'neigh_op_rgt_4')
// (8, 23, 'neigh_op_bnr_4')
// (9, 21, 'neigh_op_top_4')
// (9, 22, 'local_g2_4')
// (9, 22, 'lutff_4/out')
// (9, 22, 'lutff_6/in_0')
// (9, 23, 'neigh_op_bot_4')
// (10, 21, 'neigh_op_tnl_4')
// (10, 22, 'neigh_op_lft_4')
// (10, 23, 'neigh_op_bnl_4')

wire n1232;
// (8, 21, 'neigh_op_tnr_6')
// (8, 22, 'neigh_op_rgt_6')
// (8, 23, 'neigh_op_bnr_6')
// (9, 21, 'local_g0_6')
// (9, 21, 'lutff_4/in_0')
// (9, 21, 'neigh_op_top_6')
// (9, 22, 'lutff_6/out')
// (9, 23, 'neigh_op_bot_6')
// (10, 21, 'neigh_op_tnl_6')
// (10, 22, 'neigh_op_lft_6')
// (10, 23, 'neigh_op_bnl_6')

wire n1233;
// (8, 21, 'neigh_op_tnr_7')
// (8, 22, 'neigh_op_rgt_7')
// (8, 23, 'neigh_op_bnr_7')
// (9, 21, 'local_g1_7')
// (9, 21, 'lutff_1/in_3')
// (9, 21, 'neigh_op_top_7')
// (9, 22, 'lutff_7/out')
// (9, 23, 'neigh_op_bot_7')
// (10, 21, 'neigh_op_tnl_7')
// (10, 22, 'neigh_op_lft_7')
// (10, 23, 'neigh_op_bnl_7')

wire n1234;
// (9, 0, 'logic_op_tnr_0')
// (9, 1, 'neigh_op_rgt_0')
// (9, 2, 'local_g0_0')
// (9, 2, 'lutff_1/in_1')
// (9, 2, 'neigh_op_bnr_0')
// (10, 0, 'logic_op_top_0')
// (10, 1, 'lutff_0/out')
// (10, 2, 'neigh_op_bot_0')
// (11, 0, 'logic_op_tnl_0')
// (11, 1, 'neigh_op_lft_0')
// (11, 2, 'neigh_op_bnl_0')

reg n1235 = 0;
// (9, 0, 'logic_op_tnr_1')
// (9, 1, 'neigh_op_rgt_1')
// (9, 2, 'neigh_op_bnr_1')
// (9, 2, 'sp4_r_v_b_39')
// (9, 3, 'sp4_r_v_b_26')
// (9, 4, 'sp4_r_v_b_15')
// (9, 5, 'sp4_r_v_b_2')
// (10, 0, 'logic_op_top_1')
// (10, 1, 'local_g2_1')
// (10, 1, 'lutff_1/out')
// (10, 1, 'lutff_6/in_3')
// (10, 1, 'sp4_h_r_2')
// (10, 1, 'sp4_v_t_39')
// (10, 2, 'neigh_op_bot_1')
// (10, 2, 'sp4_v_b_39')
// (10, 3, 'sp4_v_b_26')
// (10, 4, 'local_g1_7')
// (10, 4, 'lutff_0/in_0')
// (10, 4, 'sp4_v_b_15')
// (10, 5, 'sp4_v_b_2')
// (11, 0, 'logic_op_tnl_1')
// (11, 1, 'neigh_op_lft_1')
// (11, 1, 'sp4_h_r_15')
// (11, 2, 'neigh_op_bnl_1')
// (12, 1, 'sp4_h_r_26')
// (13, 1, 'sp4_h_r_39')
// (14, 1, 'sp4_h_l_39')

reg n1236 = 0;
// (9, 0, 'logic_op_tnr_2')
// (9, 1, 'neigh_op_rgt_2')
// (9, 1, 'sp4_r_v_b_36')
// (9, 2, 'neigh_op_bnr_2')
// (9, 2, 'sp4_r_v_b_25')
// (9, 3, 'sp4_r_v_b_12')
// (9, 4, 'sp4_r_v_b_1')
// (10, 0, 'logic_op_top_2')
// (10, 0, 'span4_vert_36')
// (10, 1, 'local_g1_2')
// (10, 1, 'lutff_0/in_3')
// (10, 1, 'lutff_2/out')
// (10, 1, 'sp4_v_b_36')
// (10, 2, 'neigh_op_bot_2')
// (10, 2, 'sp4_v_b_25')
// (10, 3, 'sp4_v_b_12')
// (10, 4, 'local_g1_1')
// (10, 4, 'lutff_2/in_2')
// (10, 4, 'sp4_v_b_1')
// (11, 0, 'logic_op_tnl_2')
// (11, 1, 'neigh_op_lft_2')
// (11, 2, 'neigh_op_bnl_2')

reg n1237 = 0;
// (9, 0, 'logic_op_tnr_3')
// (9, 1, 'neigh_op_rgt_3')
// (9, 2, 'neigh_op_bnr_3')
// (10, 0, 'logic_op_top_3')
// (10, 1, 'local_g2_3')
// (10, 1, 'lutff_3/out')
// (10, 1, 'lutff_4/in_1')
// (10, 2, 'local_g0_3')
// (10, 2, 'lutff_4/in_3')
// (10, 2, 'neigh_op_bot_3')
// (11, 0, 'logic_op_tnl_3')
// (11, 1, 'neigh_op_lft_3')
// (11, 2, 'neigh_op_bnl_3')

wire n1238;
// (9, 0, 'logic_op_tnr_4')
// (9, 1, 'neigh_op_rgt_4')
// (9, 2, 'local_g0_4')
// (9, 2, 'lutff_1/in_3')
// (9, 2, 'neigh_op_bnr_4')
// (10, 0, 'logic_op_top_4')
// (10, 1, 'lutff_4/out')
// (10, 2, 'neigh_op_bot_4')
// (11, 0, 'logic_op_tnl_4')
// (11, 1, 'neigh_op_lft_4')
// (11, 2, 'neigh_op_bnl_4')

reg n1239 = 0;
// (9, 0, 'logic_op_tnr_5')
// (9, 1, 'neigh_op_rgt_5')
// (9, 2, 'local_g1_5')
// (9, 2, 'lutff_4/in_2')
// (9, 2, 'neigh_op_bnr_5')
// (10, 0, 'logic_op_top_5')
// (10, 1, 'local_g1_5')
// (10, 1, 'lutff_4/in_2')
// (10, 1, 'lutff_5/out')
// (10, 2, 'neigh_op_bot_5')
// (11, 0, 'logic_op_tnl_5')
// (11, 1, 'neigh_op_lft_5')
// (11, 2, 'neigh_op_bnl_5')

wire n1240;
// (9, 0, 'logic_op_tnr_6')
// (9, 1, 'local_g3_6')
// (9, 1, 'lutff_6/in_1')
// (9, 1, 'neigh_op_rgt_6')
// (9, 2, 'neigh_op_bnr_6')
// (10, 0, 'logic_op_top_6')
// (10, 1, 'lutff_6/out')
// (10, 2, 'neigh_op_bot_6')
// (11, 0, 'logic_op_tnl_6')
// (11, 1, 'neigh_op_lft_6')
// (11, 2, 'neigh_op_bnl_6')

reg n1241 = 0;
// (9, 0, 'logic_op_tnr_7')
// (9, 1, 'neigh_op_rgt_7')
// (9, 2, 'neigh_op_bnr_7')
// (10, 0, 'logic_op_top_7')
// (10, 1, 'local_g0_7')
// (10, 1, 'lutff_6/in_1')
// (10, 1, 'lutff_7/out')
// (10, 2, 'local_g0_7')
// (10, 2, 'lutff_0/in_3')
// (10, 2, 'neigh_op_bot_7')
// (11, 0, 'logic_op_tnl_7')
// (11, 1, 'neigh_op_lft_7')
// (11, 2, 'neigh_op_bnl_7')

wire n1242;
// (9, 1, 'local_g3_1')
// (9, 1, 'lutff_0/in_0')
// (9, 1, 'neigh_op_tnr_1')
// (9, 2, 'neigh_op_rgt_1')
// (9, 3, 'local_g0_1')
// (9, 3, 'lutff_3/in_0')
// (9, 3, 'neigh_op_bnr_1')
// (10, 1, 'neigh_op_top_1')
// (10, 2, 'lutff_1/out')
// (10, 3, 'neigh_op_bot_1')
// (11, 1, 'neigh_op_tnl_1')
// (11, 2, 'neigh_op_lft_1')
// (11, 3, 'neigh_op_bnl_1')

wire n1243;
// (9, 1, 'local_g3_2')
// (9, 1, 'lutff_6/in_3')
// (9, 1, 'neigh_op_tnr_2')
// (9, 2, 'neigh_op_rgt_2')
// (9, 3, 'neigh_op_bnr_2')
// (10, 1, 'neigh_op_top_2')
// (10, 2, 'lutff_2/out')
// (10, 3, 'neigh_op_bot_2')
// (11, 1, 'neigh_op_tnl_2')
// (11, 2, 'neigh_op_lft_2')
// (11, 3, 'neigh_op_bnl_2')

wire n1244;
// (9, 1, 'neigh_op_tnr_0')
// (9, 2, 'neigh_op_rgt_0')
// (9, 3, 'local_g0_0')
// (9, 3, 'lutff_7/in_1')
// (9, 3, 'neigh_op_bnr_0')
// (10, 1, 'neigh_op_top_0')
// (10, 2, 'lutff_0/out')
// (10, 3, 'neigh_op_bot_0')
// (11, 1, 'neigh_op_tnl_0')
// (11, 2, 'neigh_op_lft_0')
// (11, 3, 'neigh_op_bnl_0')

wire n1245;
// (9, 1, 'neigh_op_tnr_3')
// (9, 2, 'local_g3_3')
// (9, 2, 'lutff_0/in_2')
// (9, 2, 'neigh_op_rgt_3')
// (9, 3, 'neigh_op_bnr_3')
// (10, 1, 'neigh_op_top_3')
// (10, 2, 'lutff_3/out')
// (10, 3, 'neigh_op_bot_3')
// (11, 1, 'neigh_op_tnl_3')
// (11, 2, 'neigh_op_lft_3')
// (11, 3, 'neigh_op_bnl_3')

wire n1246;
// (9, 1, 'neigh_op_tnr_4')
// (9, 2, 'neigh_op_rgt_4')
// (9, 3, 'neigh_op_bnr_4')
// (10, 1, 'neigh_op_top_4')
// (10, 2, 'lutff_4/out')
// (10, 3, 'local_g1_4')
// (10, 3, 'lutff_3/in_0')
// (10, 3, 'neigh_op_bot_4')
// (11, 1, 'neigh_op_tnl_4')
// (11, 2, 'neigh_op_lft_4')
// (11, 3, 'neigh_op_bnl_4')

reg n1247 = 0;
// (9, 1, 'neigh_op_tnr_5')
// (9, 2, 'neigh_op_rgt_5')
// (9, 3, 'neigh_op_bnr_5')
// (10, 1, 'neigh_op_top_5')
// (10, 2, 'local_g1_5')
// (10, 2, 'lutff_5/out')
// (10, 2, 'lutff_6/in_0')
// (10, 3, 'local_g1_5')
// (10, 3, 'lutff_6/in_2')
// (10, 3, 'neigh_op_bot_5')
// (11, 1, 'neigh_op_tnl_5')
// (11, 2, 'neigh_op_lft_5')
// (11, 3, 'neigh_op_bnl_5')

reg n1248 = 0;
// (9, 1, 'neigh_op_tnr_7')
// (9, 2, 'neigh_op_rgt_7')
// (9, 2, 'sp4_r_v_b_46')
// (9, 3, 'neigh_op_bnr_7')
// (9, 3, 'sp4_r_v_b_35')
// (9, 4, 'sp4_r_v_b_22')
// (9, 5, 'sp4_r_v_b_11')
// (10, 1, 'neigh_op_top_7')
// (10, 1, 'sp4_v_t_46')
// (10, 2, 'local_g2_7')
// (10, 2, 'lutff_6/in_1')
// (10, 2, 'lutff_7/out')
// (10, 2, 'sp4_v_b_46')
// (10, 3, 'neigh_op_bot_7')
// (10, 3, 'sp4_v_b_35')
// (10, 4, 'sp4_v_b_22')
// (10, 5, 'local_g1_3')
// (10, 5, 'lutff_5/in_3')
// (10, 5, 'sp4_v_b_11')
// (11, 1, 'neigh_op_tnl_7')
// (11, 2, 'neigh_op_lft_7')
// (11, 3, 'neigh_op_bnl_7')

wire n1249;
// (9, 1, 'sp4_r_v_b_29')
// (9, 2, 'local_g3_0')
// (9, 2, 'lutff_4/in_1')
// (9, 2, 'sp4_r_v_b_16')
// (9, 3, 'sp4_h_r_8')
// (9, 3, 'sp4_r_v_b_5')
// (10, 0, 'span4_vert_29')
// (10, 1, 'sp4_v_b_29')
// (10, 2, 'local_g2_0')
// (10, 2, 'lutff_0/in_2')
// (10, 2, 'lutff_3/in_3')
// (10, 2, 'lutff_4/in_0')
// (10, 2, 'neigh_op_tnr_0')
// (10, 2, 'sp4_v_b_16')
// (10, 3, 'neigh_op_rgt_0')
// (10, 3, 'sp4_h_r_21')
// (10, 3, 'sp4_h_r_5')
// (10, 3, 'sp4_v_b_5')
// (10, 4, 'local_g0_0')
// (10, 4, 'lutff_0/in_2')
// (10, 4, 'lutff_2/in_0')
// (10, 4, 'neigh_op_bnr_0')
// (11, 2, 'local_g0_0')
// (11, 2, 'lutff_2/in_2')
// (11, 2, 'neigh_op_top_0')
// (11, 3, 'local_g3_0')
// (11, 3, 'lutff_0/out')
// (11, 3, 'lutff_6/in_1')
// (11, 3, 'sp4_h_r_0')
// (11, 3, 'sp4_h_r_16')
// (11, 3, 'sp4_h_r_32')
// (11, 4, 'neigh_op_bot_0')
// (12, 2, 'neigh_op_tnl_0')
// (12, 3, 'neigh_op_lft_0')
// (12, 3, 'sp4_h_r_13')
// (12, 3, 'sp4_h_r_29')
// (12, 3, 'sp4_h_r_45')
// (12, 4, 'local_g3_0')
// (12, 4, 'lutff_4/in_3')
// (12, 4, 'neigh_op_bnl_0')
// (12, 4, 'sp4_r_v_b_45')
// (12, 5, 'sp4_r_v_b_32')
// (12, 6, 'sp4_r_v_b_21')
// (12, 7, 'sp4_r_v_b_8')
// (13, 3, 'sp4_h_l_45')
// (13, 3, 'sp4_h_r_24')
// (13, 3, 'sp4_h_r_40')
// (13, 3, 'sp4_v_t_45')
// (13, 4, 'local_g3_7')
// (13, 4, 'lutff_3/in_1')
// (13, 4, 'sp4_r_v_b_47')
// (13, 4, 'sp4_v_b_45')
// (13, 5, 'local_g2_0')
// (13, 5, 'lutff_3/in_1')
// (13, 5, 'lutff_6/in_0')
// (13, 5, 'sp4_r_v_b_34')
// (13, 5, 'sp4_v_b_32')
// (13, 6, 'sp4_r_v_b_23')
// (13, 6, 'sp4_v_b_21')
// (13, 7, 'sp4_r_v_b_10')
// (13, 7, 'sp4_v_b_8')
// (14, 3, 'sp4_h_l_40')
// (14, 3, 'sp4_h_r_37')
// (14, 3, 'sp4_v_t_47')
// (14, 4, 'local_g3_7')
// (14, 4, 'lutff_6/in_2')
// (14, 4, 'sp4_r_v_b_40')
// (14, 4, 'sp4_v_b_47')
// (14, 5, 'local_g2_2')
// (14, 5, 'lutff_4/in_2')
// (14, 5, 'sp4_r_v_b_29')
// (14, 5, 'sp4_v_b_34')
// (14, 6, 'sp4_r_v_b_16')
// (14, 6, 'sp4_v_b_23')
// (14, 7, 'sp4_r_v_b_5')
// (14, 7, 'sp4_v_b_10')
// (15, 3, 'sp4_h_l_37')
// (15, 3, 'sp4_v_t_40')
// (15, 4, 'local_g3_0')
// (15, 4, 'lutff_0/in_3')
// (15, 4, 'lutff_6/in_3')
// (15, 4, 'sp4_v_b_40')
// (15, 5, 'sp4_v_b_29')
// (15, 6, 'sp4_v_b_16')
// (15, 7, 'sp4_v_b_5')

wire n1250;
// (9, 1, 'sp4_r_v_b_37')
// (9, 2, 'sp4_r_v_b_24')
// (9, 3, 'neigh_op_tnr_0')
// (9, 3, 'sp4_r_v_b_13')
// (9, 4, 'local_g1_0')
// (9, 4, 'lutff_3/in_0')
// (9, 4, 'neigh_op_rgt_0')
// (9, 4, 'sp4_r_v_b_0')
// (9, 5, 'neigh_op_bnr_0')
// (10, 0, 'span4_vert_37')
// (10, 1, 'sp4_v_b_37')
// (10, 2, 'sp4_v_b_24')
// (10, 3, 'neigh_op_top_0')
// (10, 3, 'sp4_v_b_13')
// (10, 4, 'lutff_0/out')
// (10, 4, 'sp4_v_b_0')
// (10, 5, 'neigh_op_bot_0')
// (11, 3, 'neigh_op_tnl_0')
// (11, 4, 'neigh_op_lft_0')
// (11, 5, 'neigh_op_bnl_0')

wire n1251;
// (9, 2, 'local_g2_2')
// (9, 2, 'lutff_0/in_0')
// (9, 2, 'neigh_op_tnr_2')
// (9, 3, 'neigh_op_rgt_2')
// (9, 4, 'neigh_op_bnr_2')
// (10, 2, 'neigh_op_top_2')
// (10, 3, 'lutff_2/out')
// (10, 4, 'neigh_op_bot_2')
// (11, 2, 'neigh_op_tnl_2')
// (11, 3, 'neigh_op_lft_2')
// (11, 4, 'neigh_op_bnl_2')

wire n1252;
// (9, 2, 'local_g3_1')
// (9, 2, 'lutff_2/in_0')
// (9, 2, 'neigh_op_tnr_1')
// (9, 3, 'neigh_op_rgt_1')
// (9, 4, 'neigh_op_bnr_1')
// (10, 2, 'neigh_op_top_1')
// (10, 3, 'lutff_1/out')
// (10, 4, 'neigh_op_bot_1')
// (11, 2, 'neigh_op_tnl_1')
// (11, 3, 'neigh_op_lft_1')
// (11, 4, 'neigh_op_bnl_1')

reg n1253 = 0;
// (9, 2, 'neigh_op_tnr_0')
// (9, 3, 'neigh_op_rgt_0')
// (9, 4, 'neigh_op_bnr_0')
// (10, 2, 'neigh_op_top_0')
// (10, 3, 'lutff_0/out')
// (10, 4, 'local_g1_0')
// (10, 4, 'lutff_5/in_2')
// (10, 4, 'neigh_op_bot_0')
// (11, 2, 'local_g2_0')
// (11, 2, 'lutff_3/in_1')
// (11, 2, 'neigh_op_tnl_0')
// (11, 3, 'neigh_op_lft_0')
// (11, 4, 'neigh_op_bnl_0')

wire n1254;
// (9, 2, 'neigh_op_tnr_4')
// (9, 3, 'local_g3_4')
// (9, 3, 'lutff_1/in_0')
// (9, 3, 'neigh_op_rgt_4')
// (9, 4, 'neigh_op_bnr_4')
// (10, 2, 'neigh_op_top_4')
// (10, 3, 'lutff_4/out')
// (10, 4, 'neigh_op_bot_4')
// (11, 2, 'neigh_op_tnl_4')
// (11, 3, 'neigh_op_lft_4')
// (11, 4, 'neigh_op_bnl_4')

reg n1255 = 0;
// (9, 2, 'neigh_op_tnr_5')
// (9, 3, 'local_g3_5')
// (9, 3, 'lutff_5/in_1')
// (9, 3, 'neigh_op_rgt_5')
// (9, 4, 'neigh_op_bnr_5')
// (10, 2, 'neigh_op_top_5')
// (10, 3, 'lutff_5/out')
// (10, 3, 'sp4_r_v_b_43')
// (10, 4, 'neigh_op_bot_5')
// (10, 4, 'sp4_r_v_b_30')
// (10, 5, 'local_g3_3')
// (10, 5, 'lutff_7/in_3')
// (10, 5, 'sp4_r_v_b_19')
// (10, 6, 'sp4_r_v_b_6')
// (11, 2, 'neigh_op_tnl_5')
// (11, 2, 'sp4_v_t_43')
// (11, 3, 'neigh_op_lft_5')
// (11, 3, 'sp4_v_b_43')
// (11, 4, 'neigh_op_bnl_5')
// (11, 4, 'sp4_v_b_30')
// (11, 5, 'sp4_v_b_19')
// (11, 6, 'sp4_v_b_6')

wire n1256;
// (9, 2, 'neigh_op_tnr_6')
// (9, 3, 'neigh_op_rgt_6')
// (9, 4, 'neigh_op_bnr_6')
// (10, 2, 'local_g1_6')
// (10, 2, 'lutff_0/in_1')
// (10, 2, 'neigh_op_top_6')
// (10, 3, 'lutff_6/out')
// (10, 4, 'neigh_op_bot_6')
// (11, 2, 'neigh_op_tnl_6')
// (11, 3, 'neigh_op_lft_6')
// (11, 4, 'neigh_op_bnl_6')

reg n1257 = 0;
// (9, 2, 'sp4_r_v_b_45')
// (9, 3, 'sp4_r_v_b_32')
// (9, 4, 'neigh_op_tnr_4')
// (9, 4, 'sp4_r_v_b_21')
// (9, 5, 'neigh_op_rgt_4')
// (9, 5, 'sp4_r_v_b_8')
// (9, 6, 'neigh_op_bnr_4')
// (10, 1, 'sp4_v_t_45')
// (10, 2, 'sp4_v_b_45')
// (10, 3, 'local_g2_0')
// (10, 3, 'lutff_7/in_3')
// (10, 3, 'sp4_v_b_32')
// (10, 4, 'local_g0_4')
// (10, 4, 'lutff_4/in_0')
// (10, 4, 'neigh_op_top_4')
// (10, 4, 'sp4_v_b_21')
// (10, 5, 'lutff_4/out')
// (10, 5, 'sp4_v_b_8')
// (10, 6, 'neigh_op_bot_4')
// (11, 4, 'neigh_op_tnl_4')
// (11, 5, 'neigh_op_lft_4')
// (11, 6, 'neigh_op_bnl_4')

wire n1258;
// (9, 3, 'local_g2_4')
// (9, 3, 'lutff_1/in_1')
// (9, 3, 'neigh_op_tnr_4')
// (9, 4, 'neigh_op_rgt_4')
// (9, 5, 'neigh_op_bnr_4')
// (10, 3, 'neigh_op_top_4')
// (10, 4, 'lutff_4/out')
// (10, 5, 'neigh_op_bot_4')
// (11, 3, 'neigh_op_tnl_4')
// (11, 4, 'neigh_op_lft_4')
// (11, 5, 'neigh_op_bnl_4')

wire n1259;
// (9, 3, 'neigh_op_tnr_2')
// (9, 4, 'neigh_op_rgt_2')
// (9, 5, 'neigh_op_bnr_2')
// (10, 3, 'neigh_op_top_2')
// (10, 4, 'local_g0_2')
// (10, 4, 'lutff_2/out')
// (10, 4, 'lutff_5/in_1')
// (10, 5, 'neigh_op_bot_2')
// (11, 3, 'neigh_op_tnl_2')
// (11, 4, 'neigh_op_lft_2')
// (11, 5, 'neigh_op_bnl_2')

wire n1260;
// (9, 3, 'neigh_op_tnr_3')
// (9, 4, 'neigh_op_rgt_3')
// (9, 5, 'neigh_op_bnr_3')
// (10, 3, 'neigh_op_top_3')
// (10, 4, 'local_g2_3')
// (10, 4, 'lutff_0/in_3')
// (10, 4, 'lutff_3/out')
// (10, 5, 'neigh_op_bot_3')
// (11, 3, 'neigh_op_tnl_3')
// (11, 4, 'neigh_op_lft_3')
// (11, 5, 'neigh_op_bnl_3')

wire n1261;
// (9, 3, 'neigh_op_tnr_6')
// (9, 4, 'neigh_op_rgt_6')
// (9, 5, 'local_g1_6')
// (9, 5, 'lutff_2/in_1')
// (9, 5, 'neigh_op_bnr_6')
// (10, 3, 'neigh_op_top_6')
// (10, 4, 'lutff_6/out')
// (10, 5, 'neigh_op_bot_6')
// (11, 3, 'neigh_op_tnl_6')
// (11, 4, 'neigh_op_lft_6')
// (11, 5, 'neigh_op_bnl_6')

reg n1262 = 0;
// (9, 3, 'neigh_op_tnr_7')
// (9, 4, 'neigh_op_rgt_7')
// (9, 5, 'neigh_op_bnr_7')
// (10, 3, 'local_g1_7')
// (10, 3, 'lutff_1/in_1')
// (10, 3, 'neigh_op_top_7')
// (10, 4, 'local_g2_7')
// (10, 4, 'lutff_3/in_0')
// (10, 4, 'lutff_7/out')
// (10, 5, 'neigh_op_bot_7')
// (11, 3, 'neigh_op_tnl_7')
// (11, 4, 'neigh_op_lft_7')
// (11, 5, 'neigh_op_bnl_7')

wire n1263;
// (9, 3, 'sp4_h_r_1')
// (10, 3, 'local_g0_4')
// (10, 3, 'lutff_2/in_0')
// (10, 3, 'sp4_h_r_12')
// (11, 3, 'sp4_h_r_25')
// (12, 1, 'neigh_op_tnr_6')
// (12, 1, 'sp4_r_v_b_25')
// (12, 2, 'neigh_op_rgt_6')
// (12, 2, 'sp4_r_v_b_12')
// (12, 3, 'neigh_op_bnr_6')
// (12, 3, 'sp4_h_r_36')
// (12, 3, 'sp4_r_v_b_1')
// (13, 0, 'span4_vert_25')
// (13, 1, 'neigh_op_top_6')
// (13, 1, 'sp4_v_b_25')
// (13, 2, 'lutff_6/out')
// (13, 2, 'sp4_v_b_12')
// (13, 3, 'neigh_op_bot_6')
// (13, 3, 'sp4_h_l_36')
// (13, 3, 'sp4_v_b_1')
// (14, 1, 'neigh_op_tnl_6')
// (14, 2, 'local_g1_6')
// (14, 2, 'lutff_7/in_2')
// (14, 2, 'neigh_op_lft_6')
// (14, 3, 'neigh_op_bnl_6')

wire n1264;
// (9, 4, 'neigh_op_tnr_1')
// (9, 5, 'neigh_op_rgt_1')
// (9, 6, 'neigh_op_bnr_1')
// (10, 4, 'neigh_op_top_1')
// (10, 5, 'lutff_1/out')
// (10, 6, 'neigh_op_bot_1')
// (11, 4, 'neigh_op_tnl_1')
// (11, 5, 'local_g0_1')
// (11, 5, 'lutff_0/in_1')
// (11, 5, 'neigh_op_lft_1')
// (11, 6, 'neigh_op_bnl_1')

wire n1265;
// (9, 4, 'neigh_op_tnr_5')
// (9, 5, 'neigh_op_rgt_5')
// (9, 6, 'neigh_op_bnr_5')
// (10, 4, 'neigh_op_top_5')
// (10, 5, 'local_g2_5')
// (10, 5, 'lutff_5/out')
// (10, 5, 'lutff_7/in_2')
// (10, 6, 'neigh_op_bot_5')
// (11, 4, 'neigh_op_tnl_5')
// (11, 5, 'neigh_op_lft_5')
// (11, 6, 'neigh_op_bnl_5')

wire n1266;
// (9, 4, 'neigh_op_tnr_7')
// (9, 5, 'local_g2_7')
// (9, 5, 'lutff_0/in_1')
// (9, 5, 'neigh_op_rgt_7')
// (9, 6, 'neigh_op_bnr_7')
// (10, 4, 'neigh_op_top_7')
// (10, 5, 'lutff_7/out')
// (10, 6, 'neigh_op_bot_7')
// (11, 4, 'neigh_op_tnl_7')
// (11, 5, 'neigh_op_lft_7')
// (11, 6, 'neigh_op_bnl_7')

wire n1267;
// (9, 5, 'neigh_op_tnr_2')
// (9, 6, 'local_g3_2')
// (9, 6, 'lutff_1/in_0')
// (9, 6, 'neigh_op_rgt_2')
// (9, 6, 'sp4_r_v_b_36')
// (9, 7, 'neigh_op_bnr_2')
// (9, 7, 'sp4_r_v_b_25')
// (9, 8, 'local_g2_4')
// (9, 8, 'lutff_3/in_1')
// (9, 8, 'lutff_4/in_0')
// (9, 8, 'lutff_6/in_0')
// (9, 8, 'sp4_r_v_b_12')
// (9, 9, 'sp4_r_v_b_1')
// (10, 5, 'neigh_op_top_2')
// (10, 5, 'sp4_v_t_36')
// (10, 6, 'local_g2_2')
// (10, 6, 'lutff_2/out')
// (10, 6, 'lutff_4/in_2')
// (10, 6, 'sp4_r_v_b_37')
// (10, 6, 'sp4_v_b_36')
// (10, 7, 'local_g1_2')
// (10, 7, 'lutff_0/in_1')
// (10, 7, 'lutff_1/in_0')
// (10, 7, 'lutff_5/in_2')
// (10, 7, 'neigh_op_bot_2')
// (10, 7, 'sp4_r_v_b_24')
// (10, 7, 'sp4_v_b_25')
// (10, 8, 'local_g1_4')
// (10, 8, 'lutff_2/in_3')
// (10, 8, 'sp4_r_v_b_13')
// (10, 8, 'sp4_v_b_12')
// (10, 9, 'local_g1_0')
// (10, 9, 'lutff_0/in_1')
// (10, 9, 'lutff_4/in_1')
// (10, 9, 'lutff_6/in_3')
// (10, 9, 'sp4_r_v_b_0')
// (10, 9, 'sp4_v_b_1')
// (11, 5, 'neigh_op_tnl_2')
// (11, 5, 'sp4_v_t_37')
// (11, 6, 'neigh_op_lft_2')
// (11, 6, 'sp4_v_b_37')
// (11, 7, 'neigh_op_bnl_2')
// (11, 7, 'sp4_v_b_24')
// (11, 8, 'local_g0_5')
// (11, 8, 'lutff_3/in_2')
// (11, 8, 'lutff_5/in_2')
// (11, 8, 'lutff_6/in_3')
// (11, 8, 'sp4_v_b_13')
// (11, 9, 'local_g0_0')
// (11, 9, 'lutff_5/in_1')
// (11, 9, 'sp4_v_b_0')

wire n1268;
// (9, 5, 'neigh_op_tnr_3')
// (9, 6, 'neigh_op_rgt_3')
// (9, 6, 'sp4_r_v_b_38')
// (9, 7, 'neigh_op_bnr_3')
// (9, 7, 'sp4_r_v_b_27')
// (9, 8, 'sp4_r_v_b_14')
// (9, 9, 'sp4_r_v_b_3')
// (9, 10, 'sp4_r_v_b_38')
// (9, 11, 'sp4_r_v_b_27')
// (9, 12, 'sp4_r_v_b_14')
// (9, 13, 'sp4_r_v_b_3')
// (10, 5, 'neigh_op_top_3')
// (10, 5, 'sp12_v_t_22')
// (10, 5, 'sp4_v_t_38')
// (10, 6, 'lutff_3/out')
// (10, 6, 'sp12_v_b_22')
// (10, 6, 'sp4_r_v_b_39')
// (10, 6, 'sp4_v_b_38')
// (10, 7, 'local_g0_3')
// (10, 7, 'lutff_7/in_2')
// (10, 7, 'neigh_op_bot_3')
// (10, 7, 'sp12_v_b_21')
// (10, 7, 'sp4_r_v_b_26')
// (10, 7, 'sp4_v_b_27')
// (10, 8, 'sp12_v_b_18')
// (10, 8, 'sp4_r_v_b_15')
// (10, 8, 'sp4_v_b_14')
// (10, 9, 'sp12_v_b_17')
// (10, 9, 'sp4_r_v_b_2')
// (10, 9, 'sp4_v_b_3')
// (10, 9, 'sp4_v_t_38')
// (10, 10, 'sp12_v_b_14')
// (10, 10, 'sp4_r_v_b_47')
// (10, 10, 'sp4_v_b_38')
// (10, 11, 'local_g2_3')
// (10, 11, 'lutff_0/in_1')
// (10, 11, 'lutff_5/in_0')
// (10, 11, 'sp12_v_b_13')
// (10, 11, 'sp4_r_v_b_34')
// (10, 11, 'sp4_v_b_27')
// (10, 12, 'local_g3_2')
// (10, 12, 'lutff_0/in_3')
// (10, 12, 'sp12_v_b_10')
// (10, 12, 'sp4_r_v_b_23')
// (10, 12, 'sp4_v_b_14')
// (10, 13, 'local_g0_3')
// (10, 13, 'lutff_3/in_0')
// (10, 13, 'sp12_v_b_9')
// (10, 13, 'sp4_r_v_b_10')
// (10, 13, 'sp4_v_b_3')
// (10, 14, 'local_g3_6')
// (10, 14, 'lutff_1/in_0')
// (10, 14, 'sp12_v_b_6')
// (10, 14, 'sp4_r_v_b_47')
// (10, 15, 'local_g3_5')
// (10, 15, 'lutff_5/in_3')
// (10, 15, 'lutff_6/in_2')
// (10, 15, 'sp12_v_b_5')
// (10, 15, 'sp4_r_v_b_34')
// (10, 16, 'local_g2_2')
// (10, 16, 'lutff_2/in_0')
// (10, 16, 'lutff_4/in_0')
// (10, 16, 'sp12_v_b_2')
// (10, 16, 'sp4_r_v_b_23')
// (10, 17, 'sp12_v_b_1')
// (10, 17, 'sp4_r_v_b_10')
// (11, 5, 'neigh_op_tnl_3')
// (11, 5, 'sp4_v_t_39')
// (11, 6, 'neigh_op_lft_3')
// (11, 6, 'sp4_v_b_39')
// (11, 7, 'neigh_op_bnl_3')
// (11, 7, 'sp4_v_b_26')
// (11, 8, 'sp4_v_b_15')
// (11, 9, 'local_g0_2')
// (11, 9, 'lutff_0/in_0')
// (11, 9, 'sp4_v_b_2')
// (11, 9, 'sp4_v_t_47')
// (11, 10, 'sp4_v_b_47')
// (11, 11, 'local_g3_2')
// (11, 11, 'lutff_5/in_0')
// (11, 11, 'sp4_v_b_34')
// (11, 12, 'sp4_v_b_23')
// (11, 13, 'sp4_v_b_10')
// (11, 13, 'sp4_v_t_47')
// (11, 14, 'sp4_v_b_47')
// (11, 15, 'sp4_v_b_34')
// (11, 16, 'local_g0_7')
// (11, 16, 'lutff_1/in_0')
// (11, 16, 'sp4_v_b_23')
// (11, 17, 'sp4_v_b_10')

reg n1269 = 0;
// (9, 5, 'neigh_op_tnr_4')
// (9, 6, 'local_g3_4')
// (9, 6, 'lutff_3/in_0')
// (9, 6, 'neigh_op_rgt_4')
// (9, 7, 'neigh_op_bnr_4')
// (10, 5, 'neigh_op_top_4')
// (10, 6, 'lutff_4/out')
// (10, 7, 'neigh_op_bot_4')
// (11, 5, 'neigh_op_tnl_4')
// (11, 6, 'neigh_op_lft_4')
// (11, 7, 'neigh_op_bnl_4')

reg n1270 = 0;
// (9, 5, 'sp4_h_r_7')
// (10, 5, 'sp4_h_r_18')
// (11, 4, 'neigh_op_tnr_5')
// (11, 5, 'neigh_op_rgt_5')
// (11, 5, 'sp4_h_r_31')
// (11, 5, 'sp4_r_v_b_42')
// (11, 6, 'neigh_op_bnr_5')
// (11, 6, 'sp4_r_v_b_31')
// (11, 7, 'sp4_r_v_b_18')
// (11, 8, 'local_g1_7')
// (11, 8, 'lutff_5/in_1')
// (11, 8, 'sp4_r_v_b_7')
// (12, 4, 'neigh_op_top_5')
// (12, 4, 'sp4_v_t_42')
// (12, 5, 'lutff_5/out')
// (12, 5, 'sp4_h_r_42')
// (12, 5, 'sp4_v_b_42')
// (12, 6, 'neigh_op_bot_5')
// (12, 6, 'sp4_r_v_b_42')
// (12, 6, 'sp4_v_b_31')
// (12, 7, 'sp4_r_v_b_31')
// (12, 7, 'sp4_v_b_18')
// (12, 8, 'sp4_r_v_b_18')
// (12, 8, 'sp4_v_b_7')
// (12, 9, 'local_g1_7')
// (12, 9, 'lutff_0/in_2')
// (12, 9, 'lutff_7/in_3')
// (12, 9, 'sp4_r_v_b_7')
// (13, 4, 'local_g2_5')
// (13, 4, 'lutff_4/in_1')
// (13, 4, 'neigh_op_tnl_5')
// (13, 5, 'neigh_op_lft_5')
// (13, 5, 'sp4_h_l_42')
// (13, 5, 'sp4_v_t_42')
// (13, 6, 'neigh_op_bnl_5')
// (13, 6, 'sp4_v_b_42')
// (13, 7, 'sp4_v_b_31')
// (13, 8, 'sp4_v_b_18')
// (13, 9, 'sp4_v_b_7')

reg n1271 = 0;
// (9, 5, 'sp4_r_v_b_45')
// (9, 6, 'sp4_r_v_b_32')
// (9, 7, 'sp4_r_v_b_21')
// (9, 8, 'sp4_r_v_b_8')
// (10, 4, 'sp4_v_t_45')
// (10, 5, 'sp4_v_b_45')
// (10, 6, 'sp4_v_b_32')
// (10, 7, 'local_g0_5')
// (10, 7, 'lutff_6/in_3')
// (10, 7, 'sp4_v_b_21')
// (10, 8, 'sp4_h_r_8')
// (10, 8, 'sp4_v_b_8')
// (11, 7, 'local_g3_0')
// (11, 7, 'lutff_2/in_3')
// (11, 7, 'neigh_op_tnr_0')
// (11, 8, 'neigh_op_rgt_0')
// (11, 8, 'sp4_h_r_21')
// (11, 9, 'neigh_op_bnr_0')
// (12, 7, 'neigh_op_top_0')
// (12, 8, 'local_g2_0')
// (12, 8, 'local_g3_0')
// (12, 8, 'lutff_0/out')
// (12, 8, 'lutff_1/in_3')
// (12, 8, 'lutff_5/in_2')
// (12, 8, 'sp4_h_r_32')
// (12, 9, 'neigh_op_bot_0')
// (13, 7, 'neigh_op_tnl_0')
// (13, 8, 'neigh_op_lft_0')
// (13, 8, 'sp4_h_r_45')
// (13, 9, 'neigh_op_bnl_0')
// (14, 8, 'sp4_h_l_45')

reg n1272 = 0;
// (9, 6, 'neigh_op_tnr_0')
// (9, 7, 'neigh_op_rgt_0')
// (9, 8, 'neigh_op_bnr_0')
// (10, 6, 'neigh_op_top_0')
// (10, 7, 'local_g2_0')
// (10, 7, 'lutff_0/out')
// (10, 7, 'lutff_3/in_3')
// (10, 8, 'neigh_op_bot_0')
// (11, 6, 'neigh_op_tnl_0')
// (11, 7, 'neigh_op_lft_0')
// (11, 8, 'neigh_op_bnl_0')

reg n1273 = 0;
// (9, 6, 'neigh_op_tnr_1')
// (9, 7, 'neigh_op_rgt_1')
// (9, 8, 'neigh_op_bnr_1')
// (10, 6, 'neigh_op_top_1')
// (10, 7, 'local_g1_1')
// (10, 7, 'lutff_1/out')
// (10, 7, 'lutff_3/in_1')
// (10, 8, 'neigh_op_bot_1')
// (11, 6, 'neigh_op_tnl_1')
// (11, 7, 'neigh_op_lft_1')
// (11, 8, 'neigh_op_bnl_1')

wire n1274;
// (9, 6, 'neigh_op_tnr_2')
// (9, 7, 'neigh_op_rgt_2')
// (9, 8, 'local_g0_2')
// (9, 8, 'lutff_7/in_1')
// (9, 8, 'neigh_op_bnr_2')
// (10, 6, 'neigh_op_top_2')
// (10, 7, 'lutff_2/out')
// (10, 8, 'neigh_op_bot_2')
// (11, 6, 'neigh_op_tnl_2')
// (11, 7, 'neigh_op_lft_2')
// (11, 8, 'neigh_op_bnl_2')

wire n1275;
// (9, 6, 'neigh_op_tnr_3')
// (9, 7, 'neigh_op_rgt_3')
// (9, 8, 'neigh_op_bnr_3')
// (10, 6, 'neigh_op_top_3')
// (10, 6, 'sp12_v_t_22')
// (10, 7, 'lutff_3/out')
// (10, 7, 'sp12_v_b_22')
// (10, 8, 'neigh_op_bot_3')
// (10, 8, 'sp12_v_b_21')
// (10, 9, 'sp12_v_b_18')
// (10, 10, 'sp12_v_b_17')
// (10, 11, 'sp12_v_b_14')
// (10, 12, 'sp12_v_b_13')
// (10, 13, 'sp12_v_b_10')
// (10, 14, 'sp12_v_b_9')
// (10, 15, 'local_g2_6')
// (10, 15, 'lutff_7/in_3')
// (10, 15, 'sp12_v_b_6')
// (10, 16, 'sp12_v_b_5')
// (10, 17, 'sp12_v_b_2')
// (10, 18, 'sp12_v_b_1')
// (11, 6, 'neigh_op_tnl_3')
// (11, 7, 'neigh_op_lft_3')
// (11, 8, 'neigh_op_bnl_3')

reg n1276 = 0;
// (9, 6, 'neigh_op_tnr_5')
// (9, 7, 'neigh_op_rgt_5')
// (9, 8, 'local_g1_5')
// (9, 8, 'lutff_5/in_3')
// (9, 8, 'neigh_op_bnr_5')
// (10, 6, 'neigh_op_top_5')
// (10, 7, 'lutff_5/out')
// (10, 8, 'neigh_op_bot_5')
// (11, 6, 'neigh_op_tnl_5')
// (11, 7, 'neigh_op_lft_5')
// (11, 8, 'neigh_op_bnl_5')

reg n1277 = 0;
// (9, 6, 'neigh_op_tnr_6')
// (9, 7, 'neigh_op_rgt_6')
// (9, 8, 'neigh_op_bnr_6')
// (10, 6, 'neigh_op_top_6')
// (10, 7, 'local_g1_6')
// (10, 7, 'lutff_3/in_0')
// (10, 7, 'lutff_6/out')
// (10, 8, 'neigh_op_bot_6')
// (11, 6, 'neigh_op_tnl_6')
// (11, 7, 'neigh_op_lft_6')
// (11, 8, 'neigh_op_bnl_6')

reg n1278 = 0;
// (9, 6, 'neigh_op_tnr_7')
// (9, 7, 'neigh_op_rgt_7')
// (9, 8, 'neigh_op_bnr_7')
// (10, 6, 'neigh_op_top_7')
// (10, 7, 'lutff_7/out')
// (10, 8, 'local_g0_7')
// (10, 8, 'lutff_5/in_2')
// (10, 8, 'neigh_op_bot_7')
// (11, 6, 'neigh_op_tnl_7')
// (11, 7, 'neigh_op_lft_7')
// (11, 8, 'neigh_op_bnl_7')

wire n1279;
// (9, 6, 'sp12_h_r_1')
// (10, 6, 'sp12_h_r_2')
// (10, 6, 'sp4_h_r_6')
// (11, 5, 'local_g3_3')
// (11, 5, 'lutff_global/cen')
// (11, 5, 'neigh_op_tnr_7')
// (11, 5, 'sp4_r_v_b_43')
// (11, 6, 'neigh_op_rgt_7')
// (11, 6, 'sp12_h_r_5')
// (11, 6, 'sp4_h_r_19')
// (11, 6, 'sp4_r_v_b_30')
// (11, 6, 'sp4_r_v_b_46')
// (11, 7, 'neigh_op_bnr_7')
// (11, 7, 'sp4_r_v_b_19')
// (11, 7, 'sp4_r_v_b_35')
// (11, 8, 'sp4_r_v_b_22')
// (11, 8, 'sp4_r_v_b_6')
// (11, 9, 'sp4_r_v_b_11')
// (12, 4, 'sp4_r_v_b_39')
// (12, 4, 'sp4_v_t_43')
// (12, 5, 'neigh_op_top_7')
// (12, 5, 'sp4_r_v_b_26')
// (12, 5, 'sp4_v_b_43')
// (12, 5, 'sp4_v_t_46')
// (12, 6, 'lutff_7/out')
// (12, 6, 'sp12_h_r_6')
// (12, 6, 'sp4_h_r_30')
// (12, 6, 'sp4_r_v_b_15')
// (12, 6, 'sp4_v_b_30')
// (12, 6, 'sp4_v_b_46')
// (12, 7, 'local_g3_3')
// (12, 7, 'lutff_global/cen')
// (12, 7, 'neigh_op_bot_7')
// (12, 7, 'sp4_r_v_b_2')
// (12, 7, 'sp4_v_b_19')
// (12, 7, 'sp4_v_b_35')
// (12, 8, 'sp4_v_b_22')
// (12, 8, 'sp4_v_b_6')
// (12, 9, 'sp4_v_b_11')
// (13, 3, 'sp4_v_t_39')
// (13, 4, 'sp4_v_b_39')
// (13, 5, 'local_g2_2')
// (13, 5, 'lutff_global/cen')
// (13, 5, 'neigh_op_tnl_7')
// (13, 5, 'sp4_v_b_26')
// (13, 6, 'neigh_op_lft_7')
// (13, 6, 'sp12_h_r_9')
// (13, 6, 'sp4_h_r_43')
// (13, 6, 'sp4_v_b_15')
// (13, 7, 'neigh_op_bnl_7')
// (13, 7, 'sp4_r_v_b_43')
// (13, 7, 'sp4_v_b_2')
// (13, 8, 'sp4_r_v_b_30')
// (13, 9, 'sp4_r_v_b_19')
// (13, 10, 'sp4_r_v_b_6')
// (14, 6, 'local_g0_2')
// (14, 6, 'lutff_global/cen')
// (14, 6, 'sp12_h_r_10')
// (14, 6, 'sp4_h_l_43')
// (14, 6, 'sp4_v_t_43')
// (14, 7, 'local_g3_3')
// (14, 7, 'lutff_global/cen')
// (14, 7, 'sp4_v_b_43')
// (14, 8, 'sp4_v_b_30')
// (14, 9, 'sp4_v_b_19')
// (14, 10, 'sp4_v_b_6')
// (15, 6, 'sp12_h_r_13')
// (16, 6, 'sp12_h_r_14')
// (17, 6, 'sp12_h_r_17')
// (18, 6, 'sp12_h_r_18')
// (19, 6, 'sp12_h_r_21')
// (20, 6, 'sp12_h_r_22')
// (21, 6, 'sp12_h_l_22')

wire n1280;
// (9, 6, 'sp4_r_v_b_42')
// (9, 7, 'sp4_r_v_b_31')
// (9, 8, 'sp4_r_v_b_18')
// (9, 9, 'sp4_r_v_b_7')
// (10, 5, 'sp4_h_r_1')
// (10, 5, 'sp4_v_t_42')
// (10, 6, 'sp4_v_b_42')
// (10, 7, 'local_g3_7')
// (10, 7, 'lutff_2/in_0')
// (10, 7, 'sp4_v_b_31')
// (10, 8, 'sp4_v_b_18')
// (10, 9, 'sp4_v_b_7')
// (11, 5, 'sp4_h_r_12')
// (12, 4, 'neigh_op_tnr_2')
// (12, 5, 'neigh_op_rgt_2')
// (12, 5, 'sp4_h_r_25')
// (12, 6, 'neigh_op_bnr_2')
// (13, 4, 'neigh_op_top_2')
// (13, 5, 'lutff_2/out')
// (13, 5, 'sp4_h_r_36')
// (13, 6, 'neigh_op_bot_2')
// (14, 4, 'neigh_op_tnl_2')
// (14, 5, 'neigh_op_lft_2')
// (14, 5, 'sp4_h_l_36')
// (14, 6, 'neigh_op_bnl_2')

reg n1281 = 0;
// (9, 6, 'sp4_r_v_b_47')
// (9, 7, 'sp4_r_v_b_34')
// (9, 8, 'sp4_r_v_b_23')
// (9, 9, 'sp4_r_v_b_10')
// (10, 5, 'sp4_h_r_10')
// (10, 5, 'sp4_v_t_47')
// (10, 6, 'local_g2_7')
// (10, 6, 'lutff_4/in_3')
// (10, 6, 'sp4_v_b_47')
// (10, 7, 'sp4_v_b_34')
// (10, 8, 'sp4_v_b_23')
// (10, 9, 'sp4_v_b_10')
// (11, 4, 'neigh_op_tnr_1')
// (11, 5, 'neigh_op_rgt_1')
// (11, 5, 'sp4_h_r_23')
// (11, 6, 'neigh_op_bnr_1')
// (12, 2, 'sp4_r_v_b_38')
// (12, 3, 'sp4_r_v_b_27')
// (12, 4, 'neigh_op_top_1')
// (12, 4, 'sp4_r_v_b_14')
// (12, 5, 'lutff_1/out')
// (12, 5, 'sp4_h_r_34')
// (12, 5, 'sp4_r_v_b_3')
// (12, 6, 'neigh_op_bot_1')
// (12, 6, 'sp4_r_v_b_43')
// (12, 7, 'sp4_r_v_b_30')
// (12, 8, 'sp4_r_v_b_19')
// (12, 9, 'local_g1_6')
// (12, 9, 'lutff_4/in_3')
// (12, 9, 'sp4_r_v_b_6')
// (13, 1, 'sp4_v_t_38')
// (13, 2, 'sp4_v_b_38')
// (13, 3, 'sp4_v_b_27')
// (13, 4, 'local_g2_1')
// (13, 4, 'lutff_7/in_2')
// (13, 4, 'neigh_op_tnl_1')
// (13, 4, 'sp4_v_b_14')
// (13, 5, 'neigh_op_lft_1')
// (13, 5, 'sp4_h_r_47')
// (13, 5, 'sp4_v_b_3')
// (13, 5, 'sp4_v_t_43')
// (13, 6, 'neigh_op_bnl_1')
// (13, 6, 'sp4_v_b_43')
// (13, 7, 'sp4_v_b_30')
// (13, 8, 'sp4_v_b_19')
// (13, 9, 'local_g1_6')
// (13, 9, 'lutff_5/in_0')
// (13, 9, 'sp4_v_b_6')
// (14, 5, 'sp4_h_l_47')

wire n1282;
// (9, 7, 'neigh_op_tnr_0')
// (9, 8, 'neigh_op_rgt_0')
// (9, 9, 'neigh_op_bnr_0')
// (10, 7, 'neigh_op_top_0')
// (10, 8, 'lutff_0/out')
// (10, 9, 'neigh_op_bot_0')
// (11, 7, 'neigh_op_tnl_0')
// (11, 8, 'neigh_op_lft_0')
// (11, 9, 'local_g3_0')
// (11, 9, 'lutff_2/in_1')
// (11, 9, 'neigh_op_bnl_0')

wire n1283;
// (9, 7, 'neigh_op_tnr_1')
// (9, 7, 'sp4_r_v_b_47')
// (9, 8, 'neigh_op_rgt_1')
// (9, 8, 'sp4_r_v_b_34')
// (9, 9, 'neigh_op_bnr_1')
// (9, 9, 'sp4_r_v_b_23')
// (9, 10, 'sp4_r_v_b_10')
// (9, 11, 'sp4_r_v_b_47')
// (9, 12, 'sp4_r_v_b_34')
// (9, 13, 'sp4_r_v_b_23')
// (9, 14, 'sp4_r_v_b_10')
// (10, 6, 'sp4_v_t_47')
// (10, 7, 'neigh_op_top_1')
// (10, 7, 'sp4_v_b_47')
// (10, 8, 'lutff_1/out')
// (10, 8, 'sp4_v_b_34')
// (10, 9, 'neigh_op_bot_1')
// (10, 9, 'sp4_v_b_23')
// (10, 10, 'sp4_v_b_10')
// (10, 10, 'sp4_v_t_47')
// (10, 11, 'sp4_v_b_47')
// (10, 12, 'sp4_v_b_34')
// (10, 13, 'sp4_v_b_23')
// (10, 14, 'local_g1_2')
// (10, 14, 'lutff_5/in_0')
// (10, 14, 'sp4_v_b_10')
// (11, 7, 'neigh_op_tnl_1')
// (11, 8, 'neigh_op_lft_1')
// (11, 9, 'neigh_op_bnl_1')

reg n1284 = 0;
// (9, 7, 'neigh_op_tnr_2')
// (9, 8, 'neigh_op_rgt_2')
// (9, 9, 'neigh_op_bnr_2')
// (10, 7, 'neigh_op_top_2')
// (10, 8, 'local_g1_2')
// (10, 8, 'lutff_2/out')
// (10, 8, 'lutff_7/in_2')
// (10, 9, 'neigh_op_bot_2')
// (11, 7, 'neigh_op_tnl_2')
// (11, 8, 'neigh_op_lft_2')
// (11, 9, 'neigh_op_bnl_2')

reg n1285 = 0;
// (9, 7, 'neigh_op_tnr_3')
// (9, 8, 'neigh_op_rgt_3')
// (9, 9, 'local_g1_3')
// (9, 9, 'lutff_2/in_0')
// (9, 9, 'lutff_5/in_3')
// (9, 9, 'neigh_op_bnr_3')
// (10, 7, 'neigh_op_top_3')
// (10, 8, 'local_g2_3')
// (10, 8, 'lutff_0/in_1')
// (10, 8, 'lutff_3/out')
// (10, 9, 'local_g0_3')
// (10, 9, 'lutff_2/in_1')
// (10, 9, 'lutff_7/in_2')
// (10, 9, 'neigh_op_bot_3')
// (11, 7, 'neigh_op_tnl_3')
// (11, 8, 'neigh_op_lft_3')
// (11, 9, 'neigh_op_bnl_3')

reg n1286 = 0;
// (9, 7, 'neigh_op_tnr_4')
// (9, 8, 'neigh_op_rgt_4')
// (9, 9, 'neigh_op_bnr_4')
// (10, 7, 'neigh_op_top_4')
// (10, 8, 'local_g3_4')
// (10, 8, 'lutff_0/in_3')
// (10, 8, 'lutff_4/out')
// (10, 9, 'neigh_op_bot_4')
// (11, 7, 'neigh_op_tnl_4')
// (11, 8, 'neigh_op_lft_4')
// (11, 9, 'neigh_op_bnl_4')

wire n1287;
// (9, 7, 'neigh_op_tnr_5')
// (9, 8, 'neigh_op_rgt_5')
// (9, 9, 'neigh_op_bnr_5')
// (10, 7, 'neigh_op_top_5')
// (10, 8, 'lutff_5/out')
// (10, 8, 'sp4_r_v_b_43')
// (10, 9, 'neigh_op_bot_5')
// (10, 9, 'sp4_r_v_b_30')
// (10, 10, 'sp4_r_v_b_19')
// (10, 11, 'local_g1_6')
// (10, 11, 'lutff_4/in_1')
// (10, 11, 'sp4_r_v_b_6')
// (11, 7, 'neigh_op_tnl_5')
// (11, 7, 'sp4_v_t_43')
// (11, 8, 'neigh_op_lft_5')
// (11, 8, 'sp4_v_b_43')
// (11, 9, 'neigh_op_bnl_5')
// (11, 9, 'sp4_v_b_30')
// (11, 10, 'sp4_v_b_19')
// (11, 11, 'sp4_v_b_6')

reg n1288 = 0;
// (9, 7, 'neigh_op_tnr_6')
// (9, 8, 'neigh_op_rgt_6')
// (9, 9, 'neigh_op_bnr_6')
// (10, 7, 'neigh_op_top_6')
// (10, 8, 'local_g0_6')
// (10, 8, 'lutff_0/in_2')
// (10, 8, 'lutff_6/out')
// (10, 8, 'sp4_r_v_b_45')
// (10, 9, 'local_g1_6')
// (10, 9, 'lutff_1/in_2')
// (10, 9, 'lutff_3/in_2')
// (10, 9, 'neigh_op_bot_6')
// (10, 9, 'sp4_r_v_b_32')
// (10, 10, 'local_g3_5')
// (10, 10, 'lutff_3/in_3')
// (10, 10, 'sp4_r_v_b_21')
// (10, 11, 'sp4_r_v_b_8')
// (11, 7, 'neigh_op_tnl_6')
// (11, 7, 'sp4_v_t_45')
// (11, 8, 'neigh_op_lft_6')
// (11, 8, 'sp4_v_b_45')
// (11, 9, 'neigh_op_bnl_6')
// (11, 9, 'sp4_v_b_32')
// (11, 10, 'sp4_v_b_21')
// (11, 11, 'sp4_v_b_8')

wire n1289;
// (9, 7, 'neigh_op_tnr_7')
// (9, 8, 'neigh_op_rgt_7')
// (9, 9, 'neigh_op_bnr_7')
// (10, 7, 'neigh_op_top_7')
// (10, 8, 'lutff_7/out')
// (10, 9, 'local_g0_7')
// (10, 9, 'lutff_1/in_0')
// (10, 9, 'neigh_op_bot_7')
// (11, 7, 'neigh_op_tnl_7')
// (11, 8, 'neigh_op_lft_7')
// (11, 9, 'neigh_op_bnl_7')

reg n1290 = 0;
// (9, 7, 'sp4_h_r_1')
// (10, 7, 'local_g0_4')
// (10, 7, 'lutff_1/in_3')
// (10, 7, 'sp4_h_r_12')
// (11, 4, 'neigh_op_tnr_4')
// (11, 5, 'neigh_op_rgt_4')
// (11, 5, 'sp4_r_v_b_40')
// (11, 6, 'neigh_op_bnr_4')
// (11, 6, 'sp4_r_v_b_29')
// (11, 7, 'sp4_h_r_25')
// (11, 7, 'sp4_r_v_b_16')
// (11, 8, 'sp4_r_v_b_5')
// (12, 4, 'neigh_op_top_4')
// (12, 4, 'sp4_r_v_b_36')
// (12, 4, 'sp4_v_t_40')
// (12, 5, 'lutff_4/out')
// (12, 5, 'sp4_r_v_b_25')
// (12, 5, 'sp4_v_b_40')
// (12, 6, 'neigh_op_bot_4')
// (12, 6, 'sp4_r_v_b_12')
// (12, 6, 'sp4_v_b_29')
// (12, 7, 'sp4_h_r_36')
// (12, 7, 'sp4_r_v_b_1')
// (12, 7, 'sp4_v_b_16')
// (12, 8, 'local_g1_5')
// (12, 8, 'lutff_1/in_1')
// (12, 8, 'lutff_5/in_1')
// (12, 8, 'sp4_v_b_5')
// (13, 3, 'sp4_h_r_6')
// (13, 3, 'sp4_v_t_36')
// (13, 4, 'neigh_op_tnl_4')
// (13, 4, 'sp4_v_b_36')
// (13, 5, 'neigh_op_lft_4')
// (13, 5, 'sp4_v_b_25')
// (13, 6, 'neigh_op_bnl_4')
// (13, 6, 'sp4_v_b_12')
// (13, 7, 'sp4_h_l_36')
// (13, 7, 'sp4_v_b_1')
// (14, 3, 'local_g0_3')
// (14, 3, 'lutff_5/in_2')
// (14, 3, 'sp4_h_r_19')
// (15, 3, 'sp4_h_r_30')
// (16, 3, 'sp4_h_r_43')
// (17, 3, 'sp4_h_l_43')

reg n1291 = 0;
// (9, 7, 'sp4_r_v_b_40')
// (9, 8, 'sp4_r_v_b_29')
// (9, 9, 'sp4_r_v_b_16')
// (9, 10, 'sp4_r_v_b_5')
// (10, 6, 'sp4_v_t_40')
// (10, 7, 'sp4_v_b_40')
// (10, 8, 'local_g3_5')
// (10, 8, 'lutff_4/in_0')
// (10, 8, 'sp4_v_b_29')
// (10, 9, 'sp4_v_b_16')
// (10, 10, 'sp4_h_r_0')
// (10, 10, 'sp4_v_b_5')
// (11, 7, 'sp4_r_v_b_45')
// (11, 8, 'sp4_r_v_b_32')
// (11, 9, 'neigh_op_tnr_4')
// (11, 9, 'sp4_r_v_b_21')
// (11, 10, 'neigh_op_rgt_4')
// (11, 10, 'sp4_h_r_13')
// (11, 10, 'sp4_r_v_b_8')
// (11, 11, 'neigh_op_bnr_4')
// (12, 6, 'local_g0_0')
// (12, 6, 'lutff_0/in_0')
// (12, 6, 'sp4_h_r_8')
// (12, 6, 'sp4_v_t_45')
// (12, 7, 'sp4_v_b_45')
// (12, 8, 'sp4_v_b_32')
// (12, 9, 'local_g0_4')
// (12, 9, 'lutff_4/in_2')
// (12, 9, 'neigh_op_top_4')
// (12, 9, 'sp4_v_b_21')
// (12, 10, 'lutff_4/out')
// (12, 10, 'sp4_h_r_24')
// (12, 10, 'sp4_v_b_8')
// (12, 11, 'neigh_op_bot_4')
// (13, 6, 'sp4_h_r_21')
// (13, 9, 'local_g2_4')
// (13, 9, 'lutff_5/in_1')
// (13, 9, 'neigh_op_tnl_4')
// (13, 10, 'neigh_op_lft_4')
// (13, 10, 'sp4_h_r_37')
// (13, 11, 'neigh_op_bnl_4')
// (14, 6, 'sp4_h_r_32')
// (14, 10, 'sp4_h_l_37')
// (15, 6, 'sp4_h_r_45')
// (16, 6, 'sp4_h_l_45')

wire n1292;
// (9, 7, 'sp4_r_v_b_45')
// (9, 8, 'sp4_r_v_b_32')
// (9, 9, 'local_g3_5')
// (9, 9, 'lutff_7/in_3')
// (9, 9, 'sp4_r_v_b_21')
// (9, 10, 'sp4_r_v_b_8')
// (10, 6, 'sp4_h_r_8')
// (10, 6, 'sp4_v_t_45')
// (10, 7, 'sp4_v_b_45')
// (10, 8, 'sp4_v_b_32')
// (10, 9, 'sp4_v_b_21')
// (10, 10, 'sp4_v_b_8')
// (11, 5, 'neigh_op_tnr_0')
// (11, 6, 'neigh_op_rgt_0')
// (11, 6, 'sp4_h_r_21')
// (11, 7, 'neigh_op_bnr_0')
// (12, 5, 'neigh_op_top_0')
// (12, 6, 'lutff_0/out')
// (12, 6, 'sp4_h_r_32')
// (12, 7, 'neigh_op_bot_0')
// (13, 5, 'neigh_op_tnl_0')
// (13, 6, 'neigh_op_lft_0')
// (13, 6, 'sp4_h_r_45')
// (13, 7, 'neigh_op_bnl_0')
// (14, 6, 'sp4_h_l_45')

reg n1293 = 0;
// (9, 8, 'neigh_op_tnr_0')
// (9, 9, 'neigh_op_rgt_0')
// (9, 10, 'neigh_op_bnr_0')
// (10, 8, 'neigh_op_top_0')
// (10, 9, 'local_g0_0')
// (10, 9, 'lutff_0/out')
// (10, 9, 'lutff_7/in_1')
// (10, 10, 'neigh_op_bot_0')
// (11, 8, 'neigh_op_tnl_0')
// (11, 9, 'neigh_op_lft_0')
// (11, 10, 'neigh_op_bnl_0')

wire n1294;
// (9, 8, 'neigh_op_tnr_1')
// (9, 9, 'neigh_op_rgt_1')
// (9, 10, 'neigh_op_bnr_1')
// (9, 10, 'sp4_r_v_b_39')
// (9, 11, 'sp4_r_v_b_26')
// (9, 12, 'sp4_r_v_b_15')
// (9, 13, 'sp4_r_v_b_2')
// (10, 8, 'neigh_op_top_1')
// (10, 9, 'lutff_1/out')
// (10, 9, 'sp4_h_r_2')
// (10, 9, 'sp4_v_t_39')
// (10, 10, 'neigh_op_bot_1')
// (10, 10, 'sp4_v_b_39')
// (10, 11, 'sp4_v_b_26')
// (10, 12, 'sp4_v_b_15')
// (10, 13, 'local_g0_2')
// (10, 13, 'lutff_1/in_3')
// (10, 13, 'sp4_v_b_2')
// (11, 8, 'neigh_op_tnl_1')
// (11, 9, 'neigh_op_lft_1')
// (11, 9, 'sp4_h_r_15')
// (11, 10, 'neigh_op_bnl_1')
// (12, 9, 'sp4_h_r_26')
// (13, 9, 'sp4_h_r_39')
// (14, 9, 'sp4_h_l_39')

wire n1295;
// (9, 8, 'neigh_op_tnr_2')
// (9, 9, 'neigh_op_rgt_2')
// (9, 10, 'neigh_op_bnr_2')
// (10, 7, 'sp4_r_v_b_45')
// (10, 8, 'neigh_op_top_2')
// (10, 8, 'sp4_r_v_b_32')
// (10, 9, 'lutff_2/out')
// (10, 9, 'sp4_r_v_b_21')
// (10, 10, 'neigh_op_bot_2')
// (10, 10, 'sp4_r_v_b_8')
// (11, 6, 'sp4_v_t_45')
// (11, 7, 'sp4_v_b_45')
// (11, 8, 'neigh_op_tnl_2')
// (11, 8, 'sp4_v_b_32')
// (11, 9, 'local_g1_5')
// (11, 9, 'lutff_7/in_1')
// (11, 9, 'neigh_op_lft_2')
// (11, 9, 'sp4_v_b_21')
// (11, 10, 'neigh_op_bnl_2')
// (11, 10, 'sp4_v_b_8')

wire n1296;
// (9, 8, 'neigh_op_tnr_3')
// (9, 9, 'neigh_op_rgt_3')
// (9, 9, 'sp4_r_v_b_38')
// (9, 10, 'neigh_op_bnr_3')
// (9, 10, 'sp4_r_v_b_27')
// (9, 11, 'sp4_r_v_b_14')
// (9, 12, 'sp4_r_v_b_3')
// (10, 8, 'neigh_op_top_3')
// (10, 8, 'sp4_v_t_38')
// (10, 9, 'lutff_3/out')
// (10, 9, 'sp4_v_b_38')
// (10, 10, 'neigh_op_bot_3')
// (10, 10, 'sp4_v_b_27')
// (10, 11, 'sp4_v_b_14')
// (10, 12, 'local_g0_1')
// (10, 12, 'lutff_7/in_2')
// (10, 12, 'sp4_h_r_9')
// (10, 12, 'sp4_v_b_3')
// (11, 8, 'neigh_op_tnl_3')
// (11, 9, 'neigh_op_lft_3')
// (11, 10, 'neigh_op_bnl_3')
// (11, 12, 'sp4_h_r_20')
// (12, 12, 'sp4_h_r_33')
// (13, 12, 'sp4_h_r_44')
// (14, 12, 'sp4_h_l_44')

reg n1297 = 0;
// (9, 8, 'neigh_op_tnr_4')
// (9, 9, 'neigh_op_rgt_4')
// (9, 10, 'neigh_op_bnr_4')
// (10, 8, 'neigh_op_top_4')
// (10, 9, 'lutff_4/out')
// (10, 10, 'neigh_op_bot_4')
// (11, 8, 'neigh_op_tnl_4')
// (11, 9, 'local_g0_4')
// (11, 9, 'lutff_3/in_3')
// (11, 9, 'neigh_op_lft_4')
// (11, 10, 'neigh_op_bnl_4')

reg n1298 = 0;
// (9, 8, 'neigh_op_tnr_5')
// (9, 9, 'neigh_op_rgt_5')
// (9, 10, 'neigh_op_bnr_5')
// (10, 8, 'neigh_op_top_5')
// (10, 9, 'lutff_5/out')
// (10, 10, 'local_g1_5')
// (10, 10, 'lutff_3/in_1')
// (10, 10, 'neigh_op_bot_5')
// (11, 8, 'neigh_op_tnl_5')
// (11, 9, 'neigh_op_lft_5')
// (11, 10, 'neigh_op_bnl_5')

reg n1299 = 0;
// (9, 8, 'neigh_op_tnr_6')
// (9, 9, 'neigh_op_rgt_6')
// (9, 10, 'neigh_op_bnr_6')
// (10, 8, 'neigh_op_top_6')
// (10, 9, 'local_g0_6')
// (10, 9, 'lutff_2/in_2')
// (10, 9, 'lutff_6/out')
// (10, 10, 'neigh_op_bot_6')
// (11, 8, 'neigh_op_tnl_6')
// (11, 9, 'neigh_op_lft_6')
// (11, 10, 'neigh_op_bnl_6')

wire n1300;
// (9, 8, 'neigh_op_tnr_7')
// (9, 9, 'neigh_op_rgt_7')
// (9, 10, 'neigh_op_bnr_7')
// (10, 8, 'neigh_op_top_7')
// (10, 9, 'local_g3_7')
// (10, 9, 'lutff_3/in_1')
// (10, 9, 'lutff_7/out')
// (10, 10, 'neigh_op_bot_7')
// (11, 8, 'neigh_op_tnl_7')
// (11, 9, 'neigh_op_lft_7')
// (11, 10, 'neigh_op_bnl_7')

reg n1301 = 0;
// (9, 8, 'sp4_h_r_7')
// (10, 8, 'sp4_h_r_18')
// (11, 4, 'neigh_op_tnr_3')
// (11, 5, 'neigh_op_rgt_3')
// (11, 6, 'neigh_op_bnr_3')
// (11, 8, 'local_g2_7')
// (11, 8, 'lutff_3/in_0')
// (11, 8, 'sp4_h_r_31')
// (12, 4, 'neigh_op_top_3')
// (12, 5, 'lutff_3/out')
// (12, 5, 'sp4_r_v_b_39')
// (12, 6, 'neigh_op_bot_3')
// (12, 6, 'sp4_r_v_b_26')
// (12, 7, 'sp4_r_v_b_15')
// (12, 8, 'sp4_h_r_42')
// (12, 8, 'sp4_r_v_b_2')
// (13, 4, 'neigh_op_tnl_3')
// (13, 4, 'sp4_h_r_2')
// (13, 4, 'sp4_v_t_39')
// (13, 5, 'neigh_op_lft_3')
// (13, 5, 'sp4_v_b_39')
// (13, 6, 'neigh_op_bnl_3')
// (13, 6, 'sp4_v_b_26')
// (13, 7, 'sp4_v_b_15')
// (13, 8, 'local_g0_2')
// (13, 8, 'lutff_4/in_2')
// (13, 8, 'lutff_7/in_3')
// (13, 8, 'sp4_h_l_42')
// (13, 8, 'sp4_v_b_2')
// (14, 4, 'sp4_h_r_15')
// (15, 4, 'local_g3_2')
// (15, 4, 'lutff_7/in_2')
// (15, 4, 'sp4_h_r_26')
// (16, 4, 'sp4_h_r_39')
// (17, 4, 'sp4_h_l_39')

reg n1302 = 0;
// (9, 9, 'neigh_op_tnr_0')
// (9, 10, 'neigh_op_rgt_0')
// (9, 11, 'neigh_op_bnr_0')
// (10, 9, 'neigh_op_top_0')
// (10, 10, 'local_g2_0')
// (10, 10, 'lutff_0/out')
// (10, 10, 'lutff_5/in_3')
// (10, 11, 'neigh_op_bot_0')
// (11, 9, 'neigh_op_tnl_0')
// (11, 10, 'neigh_op_lft_0')
// (11, 11, 'neigh_op_bnl_0')

reg n1303 = 0;
// (9, 9, 'neigh_op_tnr_1')
// (9, 9, 'sp4_r_v_b_47')
// (9, 10, 'neigh_op_rgt_1')
// (9, 10, 'sp4_r_v_b_34')
// (9, 11, 'neigh_op_bnr_1')
// (9, 11, 'sp4_r_v_b_23')
// (9, 12, 'sp4_r_v_b_10')
// (10, 8, 'sp4_v_t_47')
// (10, 9, 'neigh_op_top_1')
// (10, 9, 'sp4_v_b_47')
// (10, 10, 'lutff_1/out')
// (10, 10, 'sp4_v_b_34')
// (10, 11, 'neigh_op_bot_1')
// (10, 11, 'sp4_v_b_23')
// (10, 12, 'local_g0_4')
// (10, 12, 'lutff_4/in_0')
// (10, 12, 'sp4_h_r_4')
// (10, 12, 'sp4_v_b_10')
// (11, 9, 'neigh_op_tnl_1')
// (11, 10, 'neigh_op_lft_1')
// (11, 11, 'neigh_op_bnl_1')
// (11, 12, 'sp4_h_r_17')
// (12, 12, 'sp4_h_r_28')
// (13, 12, 'sp4_h_r_41')
// (14, 12, 'sp4_h_l_41')

reg n1304 = 0;
// (9, 9, 'neigh_op_tnr_2')
// (9, 10, 'neigh_op_rgt_2')
// (9, 10, 'sp4_r_v_b_36')
// (9, 11, 'neigh_op_bnr_2')
// (9, 11, 'sp4_r_v_b_25')
// (9, 12, 'sp4_r_v_b_12')
// (9, 13, 'sp4_r_v_b_1')
// (10, 9, 'neigh_op_top_2')
// (10, 9, 'sp4_v_t_36')
// (10, 10, 'lutff_2/out')
// (10, 10, 'sp4_v_b_36')
// (10, 11, 'neigh_op_bot_2')
// (10, 11, 'sp4_v_b_25')
// (10, 12, 'sp4_v_b_12')
// (10, 13, 'local_g1_1')
// (10, 13, 'lutff_0/in_2')
// (10, 13, 'sp4_v_b_1')
// (11, 9, 'neigh_op_tnl_2')
// (11, 10, 'neigh_op_lft_2')
// (11, 11, 'neigh_op_bnl_2')

wire n1305;
// (9, 9, 'neigh_op_tnr_3')
// (9, 10, 'neigh_op_rgt_3')
// (9, 11, 'neigh_op_bnr_3')
// (10, 9, 'neigh_op_top_3')
// (10, 10, 'lutff_3/out')
// (10, 11, 'local_g0_3')
// (10, 11, 'lutff_6/in_1')
// (10, 11, 'neigh_op_bot_3')
// (11, 9, 'neigh_op_tnl_3')
// (11, 10, 'neigh_op_lft_3')
// (11, 11, 'neigh_op_bnl_3')

reg n1306 = 0;
// (9, 9, 'neigh_op_tnr_4')
// (9, 10, 'local_g2_4')
// (9, 10, 'lutff_4/in_2')
// (9, 10, 'neigh_op_rgt_4')
// (9, 11, 'neigh_op_bnr_4')
// (10, 9, 'neigh_op_top_4')
// (10, 10, 'lutff_4/out')
// (10, 11, 'neigh_op_bot_4')
// (11, 9, 'neigh_op_tnl_4')
// (11, 10, 'neigh_op_lft_4')
// (11, 11, 'neigh_op_bnl_4')

wire n1307;
// (9, 9, 'neigh_op_tnr_5')
// (9, 10, 'neigh_op_rgt_5')
// (9, 11, 'neigh_op_bnr_5')
// (10, 9, 'neigh_op_top_5')
// (10, 10, 'lutff_5/out')
// (10, 11, 'neigh_op_bot_5')
// (11, 9, 'neigh_op_tnl_5')
// (11, 10, 'local_g1_5')
// (11, 10, 'lutff_5/in_1')
// (11, 10, 'neigh_op_lft_5')
// (11, 11, 'neigh_op_bnl_5')

wire n1308;
// (9, 9, 'neigh_op_tnr_6')
// (9, 10, 'neigh_op_rgt_6')
// (9, 11, 'neigh_op_bnr_6')
// (10, 9, 'neigh_op_top_6')
// (10, 10, 'local_g2_6')
// (10, 10, 'lutff_4/in_2')
// (10, 10, 'lutff_6/out')
// (10, 11, 'neigh_op_bot_6')
// (11, 9, 'neigh_op_tnl_6')
// (11, 10, 'neigh_op_lft_6')
// (11, 11, 'neigh_op_bnl_6')

reg n1309 = 0;
// (9, 9, 'neigh_op_tnr_7')
// (9, 10, 'neigh_op_rgt_7')
// (9, 11, 'neigh_op_bnr_7')
// (10, 9, 'neigh_op_top_7')
// (10, 10, 'lutff_7/out')
// (10, 11, 'local_g0_7')
// (10, 11, 'lutff_3/in_2')
// (10, 11, 'neigh_op_bot_7')
// (11, 9, 'neigh_op_tnl_7')
// (11, 10, 'neigh_op_lft_7')
// (11, 11, 'neigh_op_bnl_7')

reg n1310 = 0;
// (9, 10, 'neigh_op_tnr_0')
// (9, 11, 'neigh_op_rgt_0')
// (9, 12, 'neigh_op_bnr_0')
// (10, 10, 'neigh_op_top_0')
// (10, 11, 'local_g2_0')
// (10, 11, 'lutff_0/out')
// (10, 11, 'lutff_4/in_0')
// (10, 12, 'neigh_op_bot_0')
// (11, 10, 'neigh_op_tnl_0')
// (11, 11, 'neigh_op_lft_0')
// (11, 12, 'neigh_op_bnl_0')

reg n1311 = 0;
// (9, 10, 'neigh_op_tnr_1')
// (9, 11, 'neigh_op_rgt_1')
// (9, 12, 'neigh_op_bnr_1')
// (10, 10, 'local_g0_1')
// (10, 10, 'lutff_5/in_0')
// (10, 10, 'neigh_op_top_1')
// (10, 11, 'local_g3_1')
// (10, 11, 'lutff_1/out')
// (10, 11, 'lutff_6/in_2')
// (10, 12, 'neigh_op_bot_1')
// (11, 10, 'neigh_op_tnl_1')
// (11, 11, 'neigh_op_lft_1')
// (11, 12, 'neigh_op_bnl_1')

reg n1312 = 0;
// (9, 10, 'neigh_op_tnr_2')
// (9, 11, 'neigh_op_rgt_2')
// (9, 12, 'neigh_op_bnr_2')
// (10, 10, 'neigh_op_top_2')
// (10, 11, 'lutff_2/out')
// (10, 12, 'local_g0_2')
// (10, 12, 'lutff_7/in_3')
// (10, 12, 'neigh_op_bot_2')
// (11, 10, 'neigh_op_tnl_2')
// (11, 11, 'neigh_op_lft_2')
// (11, 12, 'neigh_op_bnl_2')

wire n1313;
// (9, 10, 'neigh_op_tnr_3')
// (9, 11, 'neigh_op_rgt_3')
// (9, 12, 'neigh_op_bnr_3')
// (10, 10, 'neigh_op_top_3')
// (10, 11, 'lutff_3/out')
// (10, 12, 'local_g0_3')
// (10, 12, 'lutff_5/in_2')
// (10, 12, 'neigh_op_bot_3')
// (11, 10, 'neigh_op_tnl_3')
// (11, 11, 'neigh_op_lft_3')
// (11, 12, 'neigh_op_bnl_3')

wire n1314;
// (9, 10, 'neigh_op_tnr_4')
// (9, 11, 'neigh_op_rgt_4')
// (9, 12, 'neigh_op_bnr_4')
// (10, 10, 'neigh_op_top_4')
// (10, 11, 'lutff_4/out')
// (10, 12, 'local_g1_4')
// (10, 12, 'lutff_3/in_2')
// (10, 12, 'neigh_op_bot_4')
// (11, 10, 'neigh_op_tnl_4')
// (11, 11, 'neigh_op_lft_4')
// (11, 12, 'neigh_op_bnl_4')

reg n1315 = 0;
// (9, 10, 'neigh_op_tnr_5')
// (9, 11, 'neigh_op_rgt_5')
// (9, 12, 'neigh_op_bnr_5')
// (10, 10, 'neigh_op_top_5')
// (10, 11, 'local_g3_5')
// (10, 11, 'lutff_3/in_1')
// (10, 11, 'lutff_5/out')
// (10, 12, 'neigh_op_bot_5')
// (11, 10, 'neigh_op_tnl_5')
// (11, 11, 'neigh_op_lft_5')
// (11, 12, 'neigh_op_bnl_5')

wire n1316;
// (9, 10, 'neigh_op_tnr_6')
// (9, 11, 'neigh_op_rgt_6')
// (9, 12, 'neigh_op_bnr_6')
// (10, 10, 'neigh_op_top_6')
// (10, 11, 'local_g2_6')
// (10, 11, 'lutff_3/in_3')
// (10, 11, 'lutff_6/out')
// (10, 12, 'neigh_op_bot_6')
// (11, 10, 'neigh_op_tnl_6')
// (11, 11, 'neigh_op_lft_6')
// (11, 12, 'neigh_op_bnl_6')

reg n1317 = 0;
// (9, 10, 'neigh_op_tnr_7')
// (9, 11, 'neigh_op_rgt_7')
// (9, 12, 'neigh_op_bnr_7')
// (10, 10, 'neigh_op_top_7')
// (10, 11, 'local_g1_7')
// (10, 11, 'lutff_6/in_0')
// (10, 11, 'lutff_7/out')
// (10, 12, 'neigh_op_bot_7')
// (11, 10, 'neigh_op_tnl_7')
// (11, 11, 'neigh_op_lft_7')
// (11, 12, 'neigh_op_bnl_7')

wire n1318;
// (9, 10, 'sp4_h_r_11')
// (10, 10, 'local_g1_6')
// (10, 10, 'lutff_4/in_1')
// (10, 10, 'sp4_h_r_22')
// (11, 4, 'neigh_op_tnr_2')
// (11, 5, 'neigh_op_rgt_2')
// (11, 6, 'neigh_op_bnr_2')
// (11, 10, 'sp4_h_r_35')
// (12, 3, 'sp4_r_v_b_45')
// (12, 4, 'neigh_op_top_2')
// (12, 4, 'sp4_r_v_b_32')
// (12, 5, 'lutff_2/out')
// (12, 5, 'sp4_r_v_b_21')
// (12, 6, 'neigh_op_bot_2')
// (12, 6, 'sp4_r_v_b_8')
// (12, 7, 'sp4_r_v_b_46')
// (12, 8, 'sp4_r_v_b_35')
// (12, 9, 'sp4_r_v_b_22')
// (12, 10, 'sp4_h_r_46')
// (12, 10, 'sp4_r_v_b_11')
// (13, 2, 'sp4_v_t_45')
// (13, 3, 'sp4_v_b_45')
// (13, 4, 'neigh_op_tnl_2')
// (13, 4, 'sp4_v_b_32')
// (13, 5, 'neigh_op_lft_2')
// (13, 5, 'sp4_v_b_21')
// (13, 6, 'neigh_op_bnl_2')
// (13, 6, 'sp4_v_b_8')
// (13, 6, 'sp4_v_t_46')
// (13, 7, 'sp4_v_b_46')
// (13, 8, 'sp4_v_b_35')
// (13, 9, 'sp4_v_b_22')
// (13, 10, 'sp4_h_l_46')
// (13, 10, 'sp4_v_b_11')

reg n1319 = 0;
// (9, 10, 'sp4_r_v_b_37')
// (9, 11, 'sp4_r_v_b_24')
// (9, 12, 'sp4_r_v_b_13')
// (9, 13, 'sp4_r_v_b_0')
// (10, 9, 'sp4_v_t_37')
// (10, 10, 'sp4_v_b_37')
// (10, 11, 'sp4_v_b_24')
// (10, 12, 'local_g0_5')
// (10, 12, 'lutff_6/in_3')
// (10, 12, 'sp4_v_b_13')
// (10, 13, 'sp4_h_r_0')
// (10, 13, 'sp4_v_b_0')
// (11, 12, 'neigh_op_tnr_4')
// (11, 13, 'neigh_op_rgt_4')
// (11, 13, 'sp4_h_r_13')
// (11, 14, 'neigh_op_bnr_4')
// (12, 12, 'neigh_op_top_4')
// (12, 13, 'lutff_4/out')
// (12, 13, 'sp4_h_r_24')
// (12, 14, 'neigh_op_bot_4')
// (13, 12, 'neigh_op_tnl_4')
// (13, 13, 'neigh_op_lft_4')
// (13, 13, 'sp4_h_r_37')
// (13, 14, 'neigh_op_bnl_4')
// (14, 13, 'sp4_h_l_37')

wire n1320;
// (9, 11, 'local_g2_0')
// (9, 11, 'lutff_7/in_3')
// (9, 11, 'neigh_op_tnr_0')
// (9, 12, 'neigh_op_rgt_0')
// (9, 13, 'neigh_op_bnr_0')
// (10, 11, 'local_g0_0')
// (10, 11, 'lutff_1/in_1')
// (10, 11, 'neigh_op_top_0')
// (10, 12, 'lutff_0/out')
// (10, 13, 'local_g1_0')
// (10, 13, 'lutff_5/in_0')
// (10, 13, 'neigh_op_bot_0')
// (11, 11, 'neigh_op_tnl_0')
// (11, 12, 'neigh_op_lft_0')
// (11, 13, 'neigh_op_bnl_0')

reg n1321 = 0;
// (9, 11, 'neigh_op_tnr_1')
// (9, 12, 'neigh_op_rgt_1')
// (9, 12, 'sp4_h_r_7')
// (9, 13, 'neigh_op_bnr_1')
// (10, 11, 'neigh_op_top_1')
// (10, 12, 'lutff_1/out')
// (10, 12, 'sp4_h_r_18')
// (10, 13, 'neigh_op_bot_1')
// (11, 11, 'neigh_op_tnl_1')
// (11, 12, 'neigh_op_lft_1')
// (11, 12, 'sp4_h_r_31')
// (11, 13, 'neigh_op_bnl_1')
// (12, 12, 'sp4_h_r_42')
// (13, 12, 'sp4_h_l_42')
// (13, 12, 'sp4_h_r_3')
// (14, 12, 'sp4_h_r_14')
// (15, 12, 'sp4_h_r_27')
// (16, 12, 'sp4_h_r_38')
// (16, 13, 'sp4_r_v_b_45')
// (16, 14, 'sp4_r_v_b_32')
// (16, 15, 'local_g3_5')
// (16, 15, 'lutff_0/in_2')
// (16, 15, 'sp4_r_v_b_21')
// (16, 16, 'sp4_r_v_b_8')
// (17, 12, 'sp4_h_l_38')
// (17, 12, 'sp4_v_t_45')
// (17, 13, 'sp4_v_b_45')
// (17, 14, 'sp4_v_b_32')
// (17, 15, 'sp4_v_b_21')
// (17, 16, 'sp4_v_b_8')

wire n1322;
// (9, 11, 'neigh_op_tnr_2')
// (9, 12, 'local_g3_2')
// (9, 12, 'lutff_1/in_2')
// (9, 12, 'neigh_op_rgt_2')
// (9, 13, 'neigh_op_bnr_2')
// (10, 11, 'neigh_op_top_2')
// (10, 12, 'lutff_2/out')
// (10, 13, 'neigh_op_bot_2')
// (11, 11, 'neigh_op_tnl_2')
// (11, 12, 'neigh_op_lft_2')
// (11, 13, 'neigh_op_bnl_2')

reg n1323 = 0;
// (9, 11, 'neigh_op_tnr_3')
// (9, 12, 'neigh_op_rgt_3')
// (9, 13, 'neigh_op_bnr_3')
// (10, 11, 'neigh_op_top_3')
// (10, 12, 'lutff_3/out')
// (10, 12, 'sp4_r_v_b_39')
// (10, 13, 'neigh_op_bot_3')
// (10, 13, 'sp4_r_v_b_26')
// (10, 14, 'sp4_r_v_b_15')
// (10, 15, 'sp4_r_v_b_2')
// (11, 11, 'neigh_op_tnl_3')
// (11, 11, 'sp4_v_t_39')
// (11, 12, 'neigh_op_lft_3')
// (11, 12, 'sp4_v_b_39')
// (11, 13, 'neigh_op_bnl_3')
// (11, 13, 'sp4_v_b_26')
// (11, 14, 'sp4_v_b_15')
// (11, 15, 'sp4_h_r_2')
// (11, 15, 'sp4_v_b_2')
// (12, 15, 'sp4_h_r_15')
// (13, 15, 'sp4_h_r_26')
// (14, 15, 'sp4_h_r_39')
// (15, 15, 'sp4_h_l_39')
// (15, 15, 'sp4_h_r_2')
// (16, 15, 'local_g1_7')
// (16, 15, 'lutff_4/in_2')
// (16, 15, 'sp4_h_r_15')
// (17, 15, 'sp4_h_r_26')
// (18, 15, 'sp4_h_r_39')
// (19, 15, 'sp4_h_l_39')

wire n1324;
// (9, 11, 'neigh_op_tnr_4')
// (9, 12, 'neigh_op_rgt_4')
// (9, 13, 'neigh_op_bnr_4')
// (10, 11, 'neigh_op_top_4')
// (10, 12, 'lutff_4/out')
// (10, 13, 'local_g0_4')
// (10, 13, 'lutff_1/in_1')
// (10, 13, 'neigh_op_bot_4')
// (11, 11, 'neigh_op_tnl_4')
// (11, 12, 'neigh_op_lft_4')
// (11, 13, 'neigh_op_bnl_4')

reg n1325 = 0;
// (9, 11, 'neigh_op_tnr_5')
// (9, 12, 'neigh_op_rgt_5')
// (9, 13, 'neigh_op_bnr_5')
// (10, 11, 'neigh_op_top_5')
// (10, 12, 'lutff_5/out')
// (10, 12, 'sp4_h_r_10')
// (10, 13, 'neigh_op_bot_5')
// (11, 11, 'neigh_op_tnl_5')
// (11, 12, 'neigh_op_lft_5')
// (11, 12, 'sp4_h_r_23')
// (11, 13, 'neigh_op_bnl_5')
// (12, 12, 'sp4_h_r_34')
// (13, 12, 'sp4_h_r_47')
// (14, 12, 'sp4_h_l_47')
// (14, 12, 'sp4_h_r_1')
// (15, 12, 'sp4_h_r_12')
// (16, 12, 'sp4_h_r_25')
// (17, 12, 'sp4_h_r_36')
// (17, 13, 'sp4_r_v_b_43')
// (17, 14, 'sp4_r_v_b_30')
// (17, 15, 'sp4_r_v_b_19')
// (17, 16, 'local_g1_6')
// (17, 16, 'lutff_3/in_2')
// (17, 16, 'sp4_r_v_b_6')
// (18, 12, 'sp4_h_l_36')
// (18, 12, 'sp4_v_t_43')
// (18, 13, 'sp4_v_b_43')
// (18, 14, 'sp4_v_b_30')
// (18, 15, 'sp4_v_b_19')
// (18, 16, 'sp4_v_b_6')

wire n1326;
// (9, 11, 'neigh_op_tnr_6')
// (9, 12, 'neigh_op_rgt_6')
// (9, 13, 'neigh_op_bnr_6')
// (10, 11, 'neigh_op_top_6')
// (10, 12, 'local_g1_6')
// (10, 12, 'lutff_1/in_0')
// (10, 12, 'lutff_6/out')
// (10, 13, 'neigh_op_bot_6')
// (11, 11, 'neigh_op_tnl_6')
// (11, 12, 'neigh_op_lft_6')
// (11, 13, 'neigh_op_bnl_6')

wire n1327;
// (9, 11, 'neigh_op_tnr_7')
// (9, 12, 'neigh_op_rgt_7')
// (9, 13, 'neigh_op_bnr_7')
// (10, 11, 'neigh_op_top_7')
// (10, 12, 'local_g3_7')
// (10, 12, 'lutff_6/in_2')
// (10, 12, 'lutff_7/out')
// (10, 13, 'neigh_op_bot_7')
// (11, 11, 'neigh_op_tnl_7')
// (11, 12, 'neigh_op_lft_7')
// (11, 13, 'neigh_op_bnl_7')

reg n1328 = 0;
// (9, 11, 'sp4_r_v_b_38')
// (9, 12, 'sp4_r_v_b_27')
// (9, 13, 'sp4_r_v_b_14')
// (9, 14, 'sp4_r_v_b_3')
// (9, 15, 'sp4_r_v_b_38')
// (9, 16, 'neigh_op_tnr_7')
// (9, 16, 'sp4_r_v_b_27')
// (9, 17, 'neigh_op_rgt_7')
// (9, 17, 'sp4_r_v_b_14')
// (9, 18, 'neigh_op_bnr_7')
// (9, 18, 'sp4_r_v_b_3')
// (10, 10, 'sp4_v_t_38')
// (10, 11, 'sp4_v_b_38')
// (10, 12, 'sp4_v_b_27')
// (10, 13, 'local_g1_6')
// (10, 13, 'lutff_6/in_3')
// (10, 13, 'sp4_v_b_14')
// (10, 14, 'sp4_v_b_3')
// (10, 14, 'sp4_v_t_38')
// (10, 15, 'sp4_v_b_38')
// (10, 16, 'neigh_op_top_7')
// (10, 16, 'sp4_v_b_27')
// (10, 17, 'lutff_7/out')
// (10, 17, 'sp4_v_b_14')
// (10, 18, 'neigh_op_bot_7')
// (10, 18, 'sp4_v_b_3')
// (11, 16, 'neigh_op_tnl_7')
// (11, 17, 'local_g0_7')
// (11, 17, 'lutff_7/in_0')
// (11, 17, 'neigh_op_lft_7')
// (11, 18, 'neigh_op_bnl_7')

reg n1329 = 0;
// (9, 12, 'local_g0_0')
// (9, 12, 'lutff_2/in_0')
// (9, 12, 'sp4_h_r_8')
// (10, 11, 'neigh_op_tnr_0')
// (10, 12, 'neigh_op_rgt_0')
// (10, 12, 'sp4_h_r_21')
// (10, 13, 'neigh_op_bnr_0')
// (11, 11, 'local_g0_0')
// (11, 11, 'lutff_3/in_1')
// (11, 11, 'neigh_op_top_0')
// (11, 12, 'local_g3_0')
// (11, 12, 'lutff_0/out')
// (11, 12, 'lutff_1/in_0')
// (11, 12, 'lutff_7/in_0')
// (11, 12, 'sp4_h_r_0')
// (11, 12, 'sp4_h_r_32')
// (11, 13, 'neigh_op_bot_0')
// (12, 11, 'local_g2_0')
// (12, 11, 'lutff_7/in_3')
// (12, 11, 'neigh_op_tnl_0')
// (12, 12, 'neigh_op_lft_0')
// (12, 12, 'sp4_h_r_13')
// (12, 12, 'sp4_h_r_45')
// (12, 13, 'neigh_op_bnl_0')
// (13, 12, 'sp4_h_l_45')
// (13, 12, 'sp4_h_r_24')
// (14, 9, 'sp4_r_v_b_37')
// (14, 10, 'sp4_r_v_b_24')
// (14, 11, 'sp4_r_v_b_13')
// (14, 12, 'sp4_h_r_37')
// (14, 12, 'sp4_r_v_b_0')
// (14, 13, 'sp4_r_v_b_40')
// (14, 14, 'sp4_r_v_b_29')
// (14, 15, 'sp4_r_v_b_16')
// (14, 16, 'sp4_r_v_b_5')
// (15, 8, 'sp4_v_t_37')
// (15, 9, 'sp4_v_b_37')
// (15, 10, 'sp4_v_b_24')
// (15, 11, 'local_g1_5')
// (15, 11, 'lutff_4/in_0')
// (15, 11, 'sp4_v_b_13')
// (15, 12, 'sp4_h_l_37')
// (15, 12, 'sp4_h_r_3')
// (15, 12, 'sp4_v_b_0')
// (15, 12, 'sp4_v_t_40')
// (15, 13, 'sp4_v_b_40')
// (15, 14, 'local_g3_5')
// (15, 14, 'lutff_0/in_0')
// (15, 14, 'sp4_v_b_29')
// (15, 15, 'sp4_v_b_16')
// (15, 16, 'sp4_v_b_5')
// (16, 12, 'sp4_h_r_14')
// (17, 12, 'local_g2_3')
// (17, 12, 'lutff_5/in_0')
// (17, 12, 'sp4_h_r_27')
// (18, 12, 'sp4_h_r_38')
// (19, 12, 'sp4_h_l_38')

reg n1330 = 0;
// (9, 12, 'local_g0_6')
// (9, 12, 'lutff_2/in_2')
// (9, 12, 'sp4_h_r_6')
// (10, 11, 'neigh_op_tnr_7')
// (10, 12, 'local_g2_7')
// (10, 12, 'lutff_2/in_1')
// (10, 12, 'neigh_op_rgt_7')
// (10, 12, 'sp4_h_r_19')
// (10, 12, 'sp4_r_v_b_46')
// (10, 13, 'neigh_op_bnr_7')
// (10, 13, 'sp4_r_v_b_35')
// (10, 14, 'sp4_r_v_b_22')
// (10, 15, 'sp4_r_v_b_11')
// (11, 11, 'local_g0_7')
// (11, 11, 'lutff_4/in_1')
// (11, 11, 'neigh_op_top_7')
// (11, 11, 'sp4_h_r_11')
// (11, 11, 'sp4_r_v_b_42')
// (11, 11, 'sp4_v_t_46')
// (11, 12, 'lutff_7/out')
// (11, 12, 'sp4_h_r_30')
// (11, 12, 'sp4_r_v_b_31')
// (11, 12, 'sp4_v_b_46')
// (11, 13, 'neigh_op_bot_7')
// (11, 13, 'sp4_r_v_b_18')
// (11, 13, 'sp4_v_b_35')
// (11, 14, 'sp4_r_v_b_7')
// (11, 14, 'sp4_v_b_22')
// (11, 15, 'sp4_v_b_11')
// (12, 10, 'sp4_v_t_42')
// (12, 11, 'local_g3_7')
// (12, 11, 'lutff_7/in_1')
// (12, 11, 'neigh_op_tnl_7')
// (12, 11, 'sp4_h_r_22')
// (12, 11, 'sp4_v_b_42')
// (12, 12, 'local_g0_7')
// (12, 12, 'lutff_4/in_3')
// (12, 12, 'lutff_7/in_2')
// (12, 12, 'neigh_op_lft_7')
// (12, 12, 'sp4_h_r_43')
// (12, 12, 'sp4_v_b_31')
// (12, 13, 'neigh_op_bnl_7')
// (12, 13, 'sp4_v_b_18')
// (12, 14, 'sp4_h_r_1')
// (12, 14, 'sp4_h_r_7')
// (12, 14, 'sp4_v_b_7')
// (13, 11, 'sp4_h_r_35')
// (13, 12, 'sp4_h_l_43')
// (13, 14, 'local_g1_4')
// (13, 14, 'lutff_0/in_3')
// (13, 14, 'sp4_h_r_12')
// (13, 14, 'sp4_h_r_18')
// (14, 11, 'sp4_h_r_46')
// (14, 14, 'sp4_h_r_25')
// (14, 14, 'sp4_h_r_31')
// (15, 11, 'local_g1_2')
// (15, 11, 'lutff_2/in_1')
// (15, 11, 'lutff_4/in_3')
// (15, 11, 'sp4_h_l_46')
// (15, 11, 'sp4_h_r_2')
// (15, 14, 'local_g2_2')
// (15, 14, 'lutff_6/in_2')
// (15, 14, 'sp4_h_r_36')
// (15, 14, 'sp4_h_r_42')
// (16, 11, 'sp4_h_r_15')
// (16, 14, 'sp4_h_l_36')
// (16, 14, 'sp4_h_l_42')
// (17, 11, 'sp4_h_r_26')
// (18, 11, 'sp4_h_r_39')
// (19, 11, 'sp4_h_l_39')

reg n1331 = 0;
// (9, 12, 'local_g3_5')
// (9, 12, 'lutff_3/in_1')
// (9, 12, 'neigh_op_tnr_5')
// (9, 13, 'neigh_op_rgt_5')
// (9, 14, 'neigh_op_bnr_5')
// (10, 12, 'neigh_op_top_5')
// (10, 13, 'lutff_5/out')
// (10, 14, 'neigh_op_bot_5')
// (11, 12, 'neigh_op_tnl_5')
// (11, 13, 'neigh_op_lft_5')
// (11, 14, 'neigh_op_bnl_5')

wire n1332;
// (9, 12, 'lutff_1/cout')
// (9, 12, 'lutff_2/in_3')

wire n1333;
// (9, 12, 'neigh_op_tnr_0')
// (9, 13, 'neigh_op_rgt_0')
// (9, 14, 'neigh_op_bnr_0')
// (10, 12, 'neigh_op_top_0')
// (10, 12, 'sp4_r_v_b_44')
// (10, 13, 'lutff_0/out')
// (10, 13, 'sp4_r_v_b_33')
// (10, 14, 'neigh_op_bot_0')
// (10, 14, 'sp4_r_v_b_20')
// (10, 15, 'sp4_r_v_b_9')
// (11, 11, 'sp4_v_t_44')
// (11, 12, 'neigh_op_tnl_0')
// (11, 12, 'sp4_v_b_44')
// (11, 13, 'neigh_op_lft_0')
// (11, 13, 'sp4_v_b_33')
// (11, 14, 'neigh_op_bnl_0')
// (11, 14, 'sp4_v_b_20')
// (11, 15, 'local_g1_1')
// (11, 15, 'lutff_2/in_0')
// (11, 15, 'sp4_v_b_9')

wire n1334;
// (9, 12, 'neigh_op_tnr_1')
// (9, 13, 'neigh_op_rgt_1')
// (9, 14, 'neigh_op_bnr_1')
// (10, 12, 'neigh_op_top_1')
// (10, 13, 'lutff_1/out')
// (10, 14, 'neigh_op_bot_1')
// (11, 12, 'neigh_op_tnl_1')
// (11, 13, 'local_g1_1')
// (11, 13, 'lutff_5/in_3')
// (11, 13, 'neigh_op_lft_1')
// (11, 14, 'neigh_op_bnl_1')

reg n1335 = 0;
// (9, 12, 'neigh_op_tnr_2')
// (9, 13, 'neigh_op_rgt_2')
// (9, 14, 'neigh_op_bnr_2')
// (10, 12, 'local_g1_2')
// (10, 12, 'lutff_4/in_1')
// (10, 12, 'neigh_op_top_2')
// (10, 13, 'lutff_2/out')
// (10, 14, 'neigh_op_bot_2')
// (11, 12, 'neigh_op_tnl_2')
// (11, 13, 'neigh_op_lft_2')
// (11, 14, 'neigh_op_bnl_2')

reg n1336 = 0;
// (9, 12, 'neigh_op_tnr_3')
// (9, 13, 'neigh_op_rgt_3')
// (9, 14, 'neigh_op_bnr_3')
// (10, 12, 'neigh_op_top_3')
// (10, 13, 'local_g2_3')
// (10, 13, 'lutff_1/in_0')
// (10, 13, 'lutff_3/out')
// (10, 14, 'neigh_op_bot_3')
// (11, 12, 'neigh_op_tnl_3')
// (11, 13, 'neigh_op_lft_3')
// (11, 14, 'neigh_op_bnl_3')

reg n1337 = 0;
// (9, 12, 'neigh_op_tnr_4')
// (9, 13, 'neigh_op_rgt_4')
// (9, 14, 'neigh_op_bnr_4')
// (10, 12, 'neigh_op_top_4')
// (10, 13, 'lutff_4/out')
// (10, 14, 'neigh_op_bot_4')
// (11, 12, 'neigh_op_tnl_4')
// (11, 13, 'local_g0_4')
// (11, 13, 'lutff_5/in_1')
// (11, 13, 'neigh_op_lft_4')
// (11, 14, 'neigh_op_bnl_4')

reg n1338 = 0;
// (9, 12, 'neigh_op_tnr_6')
// (9, 13, 'neigh_op_rgt_6')
// (9, 14, 'neigh_op_bnr_6')
// (10, 12, 'local_g0_6')
// (10, 12, 'lutff_3/in_3')
// (10, 12, 'neigh_op_top_6')
// (10, 13, 'lutff_6/out')
// (10, 14, 'neigh_op_bot_6')
// (11, 12, 'neigh_op_tnl_6')
// (11, 13, 'neigh_op_lft_6')
// (11, 14, 'neigh_op_bnl_6')

reg n1339 = 0;
// (9, 12, 'neigh_op_tnr_7')
// (9, 13, 'neigh_op_rgt_7')
// (9, 14, 'neigh_op_bnr_7')
// (10, 12, 'neigh_op_top_7')
// (10, 13, 'local_g2_7')
// (10, 13, 'lutff_0/in_3')
// (10, 13, 'lutff_7/out')
// (10, 14, 'neigh_op_bot_7')
// (11, 12, 'neigh_op_tnl_7')
// (11, 13, 'neigh_op_lft_7')
// (11, 14, 'neigh_op_bnl_7')

reg n1340 = 0;
// (9, 12, 'sp4_r_v_b_47')
// (9, 13, 'sp4_r_v_b_34')
// (9, 14, 'neigh_op_tnr_5')
// (9, 14, 'sp4_r_v_b_23')
// (9, 15, 'neigh_op_rgt_5')
// (9, 15, 'sp4_r_v_b_10')
// (9, 16, 'neigh_op_bnr_5')
// (10, 11, 'sp4_v_t_47')
// (10, 12, 'sp4_v_b_47')
// (10, 13, 'local_g3_2')
// (10, 13, 'lutff_1/in_2')
// (10, 13, 'sp4_v_b_34')
// (10, 14, 'neigh_op_top_5')
// (10, 14, 'sp4_v_b_23')
// (10, 15, 'lutff_5/out')
// (10, 15, 'sp4_v_b_10')
// (10, 16, 'neigh_op_bot_5')
// (11, 14, 'neigh_op_tnl_5')
// (11, 15, 'neigh_op_lft_5')
// (11, 16, 'neigh_op_bnl_5')

reg n1341 = 0;
// (9, 13, 'neigh_op_tnr_0')
// (9, 14, 'neigh_op_rgt_0')
// (9, 15, 'neigh_op_bnr_0')
// (10, 13, 'neigh_op_top_0')
// (10, 14, 'local_g0_0')
// (10, 14, 'lutff_0/out')
// (10, 14, 'lutff_2/in_2')
// (10, 15, 'neigh_op_bot_0')
// (11, 13, 'neigh_op_tnl_0')
// (11, 14, 'neigh_op_lft_0')
// (11, 15, 'neigh_op_bnl_0')

wire n1342;
// (9, 13, 'neigh_op_tnr_1')
// (9, 14, 'neigh_op_rgt_1')
// (9, 15, 'neigh_op_bnr_1')
// (10, 13, 'neigh_op_top_1')
// (10, 14, 'local_g0_1')
// (10, 14, 'lutff_1/out')
// (10, 14, 'lutff_3/in_2')
// (10, 14, 'lutff_4/in_1')
// (10, 15, 'neigh_op_bot_1')
// (11, 13, 'neigh_op_tnl_1')
// (11, 14, 'neigh_op_lft_1')
// (11, 15, 'neigh_op_bnl_1')

wire n1343;
// (9, 13, 'neigh_op_tnr_2')
// (9, 14, 'neigh_op_rgt_2')
// (9, 15, 'neigh_op_bnr_2')
// (10, 13, 'neigh_op_top_2')
// (10, 14, 'lutff_2/out')
// (10, 15, 'neigh_op_bot_2')
// (11, 13, 'neigh_op_tnl_2')
// (11, 14, 'local_g1_2')
// (11, 14, 'lutff_4/in_1')
// (11, 14, 'neigh_op_lft_2')
// (11, 15, 'neigh_op_bnl_2')

reg n1344 = 0;
// (9, 13, 'neigh_op_tnr_3')
// (9, 14, 'neigh_op_rgt_3')
// (9, 15, 'neigh_op_bnr_3')
// (10, 13, 'neigh_op_top_3')
// (10, 14, 'local_g2_3')
// (10, 14, 'lutff_2/in_1')
// (10, 14, 'lutff_3/out')
// (10, 15, 'neigh_op_bot_3')
// (11, 13, 'neigh_op_tnl_3')
// (11, 14, 'neigh_op_lft_3')
// (11, 15, 'neigh_op_bnl_3')

reg n1345 = 0;
// (9, 13, 'neigh_op_tnr_4')
// (9, 14, 'neigh_op_rgt_4')
// (9, 15, 'neigh_op_bnr_4')
// (10, 13, 'neigh_op_top_4')
// (10, 14, 'local_g0_4')
// (10, 14, 'lutff_4/out')
// (10, 14, 'lutff_5/in_1')
// (10, 15, 'neigh_op_bot_4')
// (11, 13, 'neigh_op_tnl_4')
// (11, 14, 'neigh_op_lft_4')
// (11, 15, 'neigh_op_bnl_4')

wire n1346;
// (9, 13, 'neigh_op_tnr_5')
// (9, 14, 'neigh_op_rgt_5')
// (9, 15, 'neigh_op_bnr_5')
// (10, 13, 'neigh_op_top_5')
// (10, 14, 'lutff_5/out')
// (10, 15, 'neigh_op_bot_5')
// (11, 13, 'neigh_op_tnl_5')
// (11, 14, 'local_g0_5')
// (11, 14, 'lutff_6/in_3')
// (11, 14, 'neigh_op_lft_5')
// (11, 15, 'neigh_op_bnl_5')

reg n1347 = 0;
// (9, 13, 'neigh_op_tnr_6')
// (9, 14, 'neigh_op_rgt_6')
// (9, 14, 'sp4_h_r_1')
// (9, 15, 'neigh_op_bnr_6')
// (10, 13, 'neigh_op_top_6')
// (10, 14, 'lutff_6/out')
// (10, 14, 'sp4_h_r_12')
// (10, 15, 'neigh_op_bot_6')
// (11, 13, 'neigh_op_tnl_6')
// (11, 14, 'local_g3_1')
// (11, 14, 'lutff_6/in_0')
// (11, 14, 'neigh_op_lft_6')
// (11, 14, 'sp4_h_r_25')
// (11, 15, 'neigh_op_bnl_6')
// (12, 14, 'sp4_h_r_36')
// (13, 14, 'sp4_h_l_36')

reg n1348 = 0;
// (9, 13, 'neigh_op_tnr_7')
// (9, 14, 'neigh_op_rgt_7')
// (9, 15, 'neigh_op_bnr_7')
// (10, 13, 'local_g1_7')
// (10, 13, 'lutff_0/in_0')
// (10, 13, 'neigh_op_top_7')
// (10, 14, 'lutff_7/out')
// (10, 15, 'neigh_op_bot_7')
// (11, 13, 'neigh_op_tnl_7')
// (11, 14, 'local_g0_7')
// (11, 14, 'lutff_3/in_0')
// (11, 14, 'neigh_op_lft_7')
// (11, 15, 'neigh_op_bnl_7')

wire n1349;
// (9, 13, 'sp4_h_r_8')
// (10, 13, 'local_g0_5')
// (10, 13, 'lutff_6/in_1')
// (10, 13, 'sp4_h_r_21')
// (11, 3, 'neigh_op_tnr_6')
// (11, 4, 'neigh_op_rgt_6')
// (11, 4, 'sp4_r_v_b_44')
// (11, 5, 'neigh_op_bnr_6')
// (11, 5, 'sp4_r_v_b_33')
// (11, 6, 'sp4_r_v_b_20')
// (11, 7, 'sp4_r_v_b_9')
// (11, 8, 'sp4_r_v_b_37')
// (11, 9, 'sp4_r_v_b_24')
// (11, 10, 'local_g2_5')
// (11, 10, 'lutff_7/in_0')
// (11, 10, 'sp4_r_v_b_13')
// (11, 11, 'sp4_r_v_b_0')
// (11, 13, 'sp4_h_r_32')
// (12, 2, 'sp4_r_v_b_37')
// (12, 3, 'neigh_op_top_6')
// (12, 3, 'sp4_r_v_b_24')
// (12, 3, 'sp4_v_t_44')
// (12, 4, 'lutff_6/out')
// (12, 4, 'sp4_r_v_b_13')
// (12, 4, 'sp4_v_b_44')
// (12, 5, 'neigh_op_bot_6')
// (12, 5, 'sp4_r_v_b_0')
// (12, 5, 'sp4_v_b_33')
// (12, 6, 'sp4_r_v_b_45')
// (12, 6, 'sp4_v_b_20')
// (12, 7, 'sp4_r_v_b_32')
// (12, 7, 'sp4_v_b_9')
// (12, 7, 'sp4_v_t_37')
// (12, 8, 'sp4_r_v_b_21')
// (12, 8, 'sp4_v_b_37')
// (12, 9, 'sp4_r_v_b_8')
// (12, 9, 'sp4_v_b_24')
// (12, 10, 'sp4_r_v_b_41')
// (12, 10, 'sp4_r_v_b_45')
// (12, 10, 'sp4_v_b_13')
// (12, 11, 'sp4_r_v_b_28')
// (12, 11, 'sp4_r_v_b_32')
// (12, 11, 'sp4_v_b_0')
// (12, 12, 'local_g3_5')
// (12, 12, 'lutff_5/in_1')
// (12, 12, 'sp4_r_v_b_17')
// (12, 12, 'sp4_r_v_b_21')
// (12, 13, 'local_g1_4')
// (12, 13, 'local_g2_0')
// (12, 13, 'lutff_1/in_1')
// (12, 13, 'lutff_3/in_1')
// (12, 13, 'lutff_4/in_0')
// (12, 13, 'lutff_5/in_0')
// (12, 13, 'lutff_6/in_2')
// (12, 13, 'lutff_7/in_2')
// (12, 13, 'sp4_h_r_45')
// (12, 13, 'sp4_r_v_b_4')
// (12, 13, 'sp4_r_v_b_8')
// (12, 14, 'sp4_r_v_b_45')
// (12, 15, 'sp4_r_v_b_32')
// (12, 16, 'local_g3_5')
// (12, 16, 'lutff_0/in_2')
// (12, 16, 'lutff_1/in_1')
// (12, 16, 'sp4_r_v_b_21')
// (12, 17, 'sp4_r_v_b_8')
// (13, 1, 'sp4_v_t_37')
// (13, 2, 'sp4_v_b_37')
// (13, 3, 'neigh_op_tnl_6')
// (13, 3, 'sp4_v_b_24')
// (13, 4, 'neigh_op_lft_6')
// (13, 4, 'sp4_v_b_13')
// (13, 5, 'neigh_op_bnl_6')
// (13, 5, 'sp4_v_b_0')
// (13, 5, 'sp4_v_t_45')
// (13, 6, 'sp4_v_b_45')
// (13, 7, 'sp4_v_b_32')
// (13, 8, 'sp4_v_b_21')
// (13, 9, 'sp4_v_b_8')
// (13, 9, 'sp4_v_t_41')
// (13, 9, 'sp4_v_t_45')
// (13, 10, 'sp4_v_b_41')
// (13, 10, 'sp4_v_b_45')
// (13, 11, 'sp4_v_b_28')
// (13, 11, 'sp4_v_b_32')
// (13, 12, 'sp4_v_b_17')
// (13, 12, 'sp4_v_b_21')
// (13, 13, 'sp4_h_l_45')
// (13, 13, 'sp4_v_b_4')
// (13, 13, 'sp4_v_b_8')
// (13, 13, 'sp4_v_t_45')
// (13, 14, 'sp4_v_b_45')
// (13, 15, 'sp4_v_b_32')
// (13, 16, 'sp4_v_b_21')
// (13, 17, 'sp4_v_b_8')

reg n1350 = 0;
// (9, 13, 'sp4_r_v_b_45')
// (9, 14, 'sp4_r_v_b_32')
// (9, 15, 'neigh_op_tnr_4')
// (9, 15, 'sp4_r_v_b_21')
// (9, 16, 'neigh_op_rgt_4')
// (9, 16, 'sp4_r_v_b_8')
// (9, 17, 'neigh_op_bnr_4')
// (10, 12, 'local_g1_1')
// (10, 12, 'lutff_7/in_1')
// (10, 12, 'sp4_h_r_1')
// (10, 12, 'sp4_v_t_45')
// (10, 13, 'sp4_v_b_45')
// (10, 14, 'sp4_v_b_32')
// (10, 15, 'neigh_op_top_4')
// (10, 15, 'sp4_v_b_21')
// (10, 16, 'lutff_4/out')
// (10, 16, 'sp4_v_b_8')
// (10, 17, 'neigh_op_bot_4')
// (11, 12, 'sp4_h_r_12')
// (11, 15, 'neigh_op_tnl_4')
// (11, 16, 'neigh_op_lft_4')
// (11, 17, 'neigh_op_bnl_4')
// (12, 12, 'sp4_h_r_25')
// (13, 12, 'sp4_h_r_36')
// (14, 12, 'sp4_h_l_36')

reg n1351 = 0;
// (9, 14, 'local_g3_2')
// (9, 14, 'lutff_1/in_2')
// (9, 14, 'neigh_op_tnr_2')
// (9, 15, 'neigh_op_rgt_2')
// (9, 16, 'neigh_op_bnr_2')
// (10, 14, 'local_g0_2')
// (10, 14, 'lutff_5/in_3')
// (10, 14, 'neigh_op_top_2')
// (10, 15, 'lutff_2/out')
// (10, 16, 'neigh_op_bot_2')
// (11, 14, 'neigh_op_tnl_2')
// (11, 15, 'neigh_op_lft_2')
// (11, 16, 'neigh_op_bnl_2')

reg n1352 = 0;
// (9, 14, 'neigh_op_tnr_0')
// (9, 15, 'neigh_op_rgt_0')
// (9, 16, 'neigh_op_bnr_0')
// (10, 14, 'neigh_op_top_0')
// (10, 15, 'local_g3_0')
// (10, 15, 'lutff_0/out')
// (10, 15, 'lutff_3/in_2')
// (10, 16, 'neigh_op_bot_0')
// (11, 14, 'neigh_op_tnl_0')
// (11, 15, 'neigh_op_lft_0')
// (11, 16, 'neigh_op_bnl_0')

reg n1353 = 0;
// (9, 14, 'neigh_op_tnr_1')
// (9, 15, 'local_g3_1')
// (9, 15, 'lutff_2/in_2')
// (9, 15, 'neigh_op_rgt_1')
// (9, 16, 'neigh_op_bnr_1')
// (10, 14, 'neigh_op_top_1')
// (10, 15, 'local_g0_1')
// (10, 15, 'lutff_1/out')
// (10, 15, 'lutff_7/in_0')
// (10, 16, 'neigh_op_bot_1')
// (11, 14, 'neigh_op_tnl_1')
// (11, 15, 'neigh_op_lft_1')
// (11, 16, 'neigh_op_bnl_1')

wire n1354;
// (9, 14, 'neigh_op_tnr_3')
// (9, 15, 'neigh_op_rgt_3')
// (9, 16, 'neigh_op_bnr_3')
// (10, 14, 'neigh_op_top_3')
// (10, 15, 'lutff_3/out')
// (10, 15, 'sp4_h_r_6')
// (10, 16, 'neigh_op_bot_3')
// (11, 14, 'neigh_op_tnl_3')
// (11, 15, 'neigh_op_lft_3')
// (11, 15, 'sp4_h_r_19')
// (11, 16, 'neigh_op_bnl_3')
// (12, 15, 'local_g2_6')
// (12, 15, 'lutff_7/in_1')
// (12, 15, 'sp4_h_r_30')
// (13, 15, 'sp4_h_r_43')
// (14, 15, 'sp4_h_l_43')

wire n1355;
// (9, 14, 'neigh_op_tnr_4')
// (9, 15, 'neigh_op_rgt_4')
// (9, 16, 'neigh_op_bnr_4')
// (10, 14, 'neigh_op_top_4')
// (10, 15, 'lutff_4/out')
// (10, 16, 'neigh_op_bot_4')
// (11, 14, 'neigh_op_tnl_4')
// (11, 15, 'local_g0_4')
// (11, 15, 'lutff_0/in_0')
// (11, 15, 'neigh_op_lft_4')
// (11, 16, 'neigh_op_bnl_4')

reg n1356 = 0;
// (9, 14, 'neigh_op_tnr_6')
// (9, 15, 'neigh_op_rgt_6')
// (9, 16, 'neigh_op_bnr_6')
// (10, 14, 'local_g1_6')
// (10, 14, 'lutff_2/in_3')
// (10, 14, 'lutff_5/in_2')
// (10, 14, 'neigh_op_top_6')
// (10, 15, 'local_g0_6')
// (10, 15, 'local_g1_6')
// (10, 15, 'lutff_3/in_3')
// (10, 15, 'lutff_6/out')
// (10, 15, 'lutff_7/in_2')
// (10, 16, 'neigh_op_bot_6')
// (11, 14, 'local_g3_6')
// (11, 14, 'lutff_3/in_2')
// (11, 14, 'neigh_op_tnl_6')
// (11, 15, 'local_g1_6')
// (11, 15, 'lutff_2/in_3')
// (11, 15, 'neigh_op_lft_6')
// (11, 16, 'neigh_op_bnl_6')

wire n1357;
// (9, 14, 'neigh_op_tnr_7')
// (9, 15, 'neigh_op_rgt_7')
// (9, 16, 'neigh_op_bnr_7')
// (10, 14, 'neigh_op_top_7')
// (10, 15, 'lutff_7/out')
// (10, 16, 'neigh_op_bot_7')
// (11, 14, 'neigh_op_tnl_7')
// (11, 15, 'local_g0_7')
// (11, 15, 'lutff_5/in_2')
// (11, 15, 'neigh_op_lft_7')
// (11, 16, 'neigh_op_bnl_7')

reg n1358 = 0;
// (9, 14, 'sp4_r_v_b_38')
// (9, 15, 'sp4_r_v_b_27')
// (9, 16, 'sp4_r_v_b_14')
// (9, 17, 'sp4_r_v_b_3')
// (10, 13, 'sp4_v_t_38')
// (10, 14, 'sp4_v_b_38')
// (10, 15, 'local_g2_3')
// (10, 15, 'lutff_5/in_2')
// (10, 15, 'sp4_v_b_27')
// (10, 16, 'sp4_v_b_14')
// (10, 17, 'sp4_h_r_10')
// (10, 17, 'sp4_v_b_3')
// (11, 16, 'neigh_op_tnr_1')
// (11, 17, 'neigh_op_rgt_1')
// (11, 17, 'sp4_h_r_23')
// (11, 18, 'neigh_op_bnr_1')
// (12, 16, 'neigh_op_top_1')
// (12, 17, 'local_g1_1')
// (12, 17, 'lutff_1/in_3')
// (12, 17, 'lutff_1/out')
// (12, 17, 'lutff_7/in_1')
// (12, 17, 'sp4_h_r_34')
// (12, 18, 'neigh_op_bot_1')
// (13, 16, 'neigh_op_tnl_1')
// (13, 17, 'neigh_op_lft_1')
// (13, 17, 'sp4_h_r_47')
// (13, 18, 'neigh_op_bnl_1')
// (14, 17, 'sp4_h_l_47')

reg n1359 = 0;
// (9, 14, 'sp4_r_v_b_46')
// (9, 15, 'local_g0_0')
// (9, 15, 'lutff_5/in_1')
// (9, 15, 'sp4_r_v_b_35')
// (9, 16, 'sp4_r_v_b_22')
// (9, 17, 'sp4_r_v_b_11')
// (10, 13, 'sp4_v_t_46')
// (10, 14, 'sp4_v_b_46')
// (10, 15, 'sp4_v_b_35')
// (10, 16, 'neigh_op_tnr_3')
// (10, 16, 'sp4_v_b_22')
// (10, 17, 'neigh_op_rgt_3')
// (10, 17, 'sp4_h_r_11')
// (10, 17, 'sp4_v_b_11')
// (10, 18, 'neigh_op_bnr_3')
// (11, 16, 'neigh_op_top_3')
// (11, 17, 'local_g2_3')
// (11, 17, 'lutff_3/out')
// (11, 17, 'lutff_7/in_2')
// (11, 17, 'sp4_h_r_22')
// (11, 18, 'neigh_op_bot_3')
// (12, 16, 'neigh_op_tnl_3')
// (12, 17, 'neigh_op_lft_3')
// (12, 17, 'sp4_h_r_35')
// (12, 18, 'neigh_op_bnl_3')
// (13, 17, 'sp4_h_r_46')
// (14, 17, 'sp4_h_l_46')

reg n1360 = 0;
// (9, 14, 'sp4_r_v_b_47')
// (9, 15, 'sp4_r_v_b_34')
// (9, 16, 'neigh_op_tnr_5')
// (9, 16, 'sp4_r_v_b_23')
// (9, 17, 'neigh_op_rgt_5')
// (9, 17, 'sp4_r_v_b_10')
// (9, 18, 'neigh_op_bnr_5')
// (10, 13, 'sp4_v_t_47')
// (10, 14, 'local_g2_7')
// (10, 14, 'lutff_6/in_1')
// (10, 14, 'sp4_v_b_47')
// (10, 15, 'local_g3_2')
// (10, 15, 'lutff_4/in_3')
// (10, 15, 'sp4_v_b_34')
// (10, 16, 'neigh_op_top_5')
// (10, 16, 'sp4_v_b_23')
// (10, 17, 'lutff_5/out')
// (10, 17, 'sp4_v_b_10')
// (10, 18, 'neigh_op_bot_5')
// (11, 16, 'neigh_op_tnl_5')
// (11, 17, 'neigh_op_lft_5')
// (11, 18, 'neigh_op_bnl_5')

reg n1361 = 0;
// (9, 15, 'neigh_op_tnr_0')
// (9, 16, 'neigh_op_rgt_0')
// (9, 17, 'neigh_op_bnr_0')
// (10, 15, 'local_g0_0')
// (10, 15, 'lutff_3/in_1')
// (10, 15, 'neigh_op_top_0')
// (10, 16, 'lutff_0/out')
// (10, 17, 'neigh_op_bot_0')
// (11, 15, 'neigh_op_tnl_0')
// (11, 16, 'neigh_op_lft_0')
// (11, 17, 'neigh_op_bnl_0')

wire n1362;
// (9, 15, 'neigh_op_tnr_2')
// (9, 16, 'neigh_op_rgt_2')
// (9, 17, 'neigh_op_bnr_2')
// (10, 15, 'neigh_op_top_2')
// (10, 16, 'local_g3_2')
// (10, 16, 'lutff_0/in_3')
// (10, 16, 'lutff_2/out')
// (10, 16, 'lutff_7/in_2')
// (10, 17, 'neigh_op_bot_2')
// (11, 15, 'neigh_op_tnl_2')
// (11, 16, 'neigh_op_lft_2')
// (11, 17, 'neigh_op_bnl_2')

reg n1363 = 0;
// (9, 15, 'neigh_op_tnr_3')
// (9, 16, 'neigh_op_rgt_3')
// (9, 17, 'neigh_op_bnr_3')
// (10, 15, 'neigh_op_top_3')
// (10, 16, 'lutff_3/out')
// (10, 17, 'neigh_op_bot_3')
// (11, 15, 'local_g2_3')
// (11, 15, 'lutff_5/in_0')
// (11, 15, 'neigh_op_tnl_3')
// (11, 16, 'neigh_op_lft_3')
// (11, 17, 'neigh_op_bnl_3')

wire n1364;
// (9, 15, 'neigh_op_tnr_6')
// (9, 16, 'neigh_op_rgt_6')
// (9, 17, 'neigh_op_bnr_6')
// (10, 15, 'neigh_op_top_6')
// (10, 16, 'lutff_6/out')
// (10, 17, 'neigh_op_bot_6')
// (11, 15, 'local_g2_6')
// (11, 15, 'lutff_1/in_1')
// (11, 15, 'neigh_op_tnl_6')
// (11, 16, 'neigh_op_lft_6')
// (11, 17, 'neigh_op_bnl_6')

reg n1365 = 0;
// (9, 15, 'neigh_op_tnr_7')
// (9, 16, 'neigh_op_rgt_7')
// (9, 17, 'neigh_op_bnr_7')
// (10, 15, 'local_g1_7')
// (10, 15, 'lutff_7/in_1')
// (10, 15, 'neigh_op_top_7')
// (10, 16, 'lutff_7/out')
// (10, 17, 'neigh_op_bot_7')
// (11, 15, 'neigh_op_tnl_7')
// (11, 16, 'neigh_op_lft_7')
// (11, 17, 'neigh_op_bnl_7')

reg n1366 = 0;
// (9, 15, 'sp4_h_r_11')
// (10, 15, 'sp4_h_r_22')
// (11, 14, 'neigh_op_tnr_7')
// (11, 15, 'neigh_op_rgt_7')
// (11, 15, 'sp4_h_r_35')
// (11, 16, 'neigh_op_bnr_7')
// (12, 14, 'neigh_op_top_7')
// (12, 15, 'lutff_7/out')
// (12, 15, 'sp4_h_r_46')
// (12, 16, 'neigh_op_bot_7')
// (13, 14, 'neigh_op_tnl_7')
// (13, 15, 'neigh_op_lft_7')
// (13, 15, 'sp4_h_l_46')
// (13, 15, 'sp4_h_r_7')
// (13, 16, 'neigh_op_bnl_7')
// (14, 15, 'sp4_h_r_18')
// (15, 15, 'sp4_h_r_31')
// (16, 15, 'local_g2_2')
// (16, 15, 'lutff_3/in_3')
// (16, 15, 'sp4_h_r_42')
// (17, 15, 'sp4_h_l_42')

reg n1367 = 0;
// (9, 15, 'sp4_r_v_b_43')
// (9, 16, 'sp4_r_v_b_30')
// (9, 17, 'sp4_r_v_b_19')
// (9, 18, 'sp4_r_v_b_6')
// (9, 19, 'sp4_r_v_b_38')
// (9, 20, 'neigh_op_tnr_7')
// (9, 20, 'sp4_r_v_b_27')
// (9, 21, 'neigh_op_rgt_7')
// (9, 21, 'sp4_r_v_b_14')
// (9, 22, 'neigh_op_bnr_7')
// (9, 22, 'sp4_r_v_b_3')
// (10, 14, 'sp4_v_t_43')
// (10, 15, 'sp4_v_b_43')
// (10, 16, 'local_g3_6')
// (10, 16, 'lutff_2/in_1')
// (10, 16, 'sp4_v_b_30')
// (10, 17, 'sp4_v_b_19')
// (10, 18, 'sp4_v_b_6')
// (10, 18, 'sp4_v_t_38')
// (10, 19, 'sp4_v_b_38')
// (10, 20, 'neigh_op_top_7')
// (10, 20, 'sp4_v_b_27')
// (10, 21, 'local_g1_7')
// (10, 21, 'lutff_4/in_2')
// (10, 21, 'lutff_7/out')
// (10, 21, 'sp4_v_b_14')
// (10, 22, 'neigh_op_bot_7')
// (10, 22, 'sp4_v_b_3')
// (11, 20, 'neigh_op_tnl_7')
// (11, 21, 'neigh_op_lft_7')
// (11, 22, 'neigh_op_bnl_7')

wire n1368;
// (9, 16, 'lutff_7/cout')
// (9, 17, 'carry_in')
// (9, 17, 'carry_in_mux')

reg n1369 = 0;
// (9, 16, 'neigh_op_tnr_1')
// (9, 17, 'neigh_op_rgt_1')
// (9, 18, 'neigh_op_bnr_1')
// (10, 16, 'neigh_op_top_1')
// (10, 17, 'lutff_1/out')
// (10, 18, 'neigh_op_bot_1')
// (11, 16, 'local_g3_1')
// (11, 16, 'lutff_0/in_2')
// (11, 16, 'neigh_op_tnl_1')
// (11, 17, 'local_g0_1')
// (11, 17, 'lutff_6/in_1')
// (11, 17, 'neigh_op_lft_1')
// (11, 18, 'neigh_op_bnl_1')

reg n1370 = 0;
// (9, 16, 'neigh_op_tnr_4')
// (9, 17, 'neigh_op_rgt_4')
// (9, 18, 'neigh_op_bnr_4')
// (10, 16, 'local_g1_4')
// (10, 16, 'lutff_3/in_2')
// (10, 16, 'lutff_6/in_1')
// (10, 16, 'neigh_op_top_4')
// (10, 17, 'lutff_4/out')
// (10, 18, 'neigh_op_bot_4')
// (11, 16, 'neigh_op_tnl_4')
// (11, 17, 'neigh_op_lft_4')
// (11, 18, 'neigh_op_bnl_4')

wire n1371;
// (9, 17, 'lutff_0/cout')
// (9, 17, 'lutff_1/in_3')

wire n1372;
// (9, 18, 'lutff_7/cout')
// (9, 19, 'carry_in')
// (9, 19, 'carry_in_mux')

wire n1373;
// (9, 18, 'neigh_op_tnr_0')
// (9, 19, 'neigh_op_rgt_0')
// (9, 20, 'neigh_op_bnr_0')
// (10, 18, 'neigh_op_top_0')
// (10, 19, 'local_g2_0')
// (10, 19, 'lutff_0/out')
// (10, 19, 'lutff_1/in_1')
// (10, 20, 'neigh_op_bot_0')
// (11, 18, 'neigh_op_tnl_0')
// (11, 19, 'neigh_op_lft_0')
// (11, 20, 'neigh_op_bnl_0')

wire n1374;
// (9, 18, 'neigh_op_tnr_3')
// (9, 19, 'neigh_op_rgt_3')
// (9, 20, 'neigh_op_bnr_3')
// (10, 18, 'neigh_op_top_3')
// (10, 19, 'local_g2_3')
// (10, 19, 'lutff_1/in_2')
// (10, 19, 'lutff_3/out')
// (10, 20, 'neigh_op_bot_3')
// (11, 18, 'neigh_op_tnl_3')
// (11, 19, 'neigh_op_lft_3')
// (11, 20, 'neigh_op_bnl_3')

wire n1375;
// (9, 18, 'neigh_op_tnr_4')
// (9, 19, 'neigh_op_rgt_4')
// (9, 20, 'neigh_op_bnr_4')
// (10, 18, 'neigh_op_top_4')
// (10, 19, 'local_g0_4')
// (10, 19, 'lutff_4/out')
// (10, 19, 'lutff_7/in_1')
// (10, 20, 'neigh_op_bot_4')
// (11, 18, 'neigh_op_tnl_4')
// (11, 19, 'neigh_op_lft_4')
// (11, 20, 'neigh_op_bnl_4')

wire n1376;
// (9, 18, 'neigh_op_tnr_5')
// (9, 19, 'neigh_op_rgt_5')
// (9, 20, 'neigh_op_bnr_5')
// (10, 18, 'neigh_op_top_5')
// (10, 19, 'local_g2_5')
// (10, 19, 'lutff_3/in_2')
// (10, 19, 'lutff_5/out')
// (10, 20, 'neigh_op_bot_5')
// (11, 18, 'neigh_op_tnl_5')
// (11, 19, 'neigh_op_lft_5')
// (11, 20, 'neigh_op_bnl_5')

wire n1377;
// (9, 18, 'neigh_op_tnr_7')
// (9, 19, 'neigh_op_rgt_7')
// (9, 20, 'neigh_op_bnr_7')
// (10, 18, 'neigh_op_top_7')
// (10, 19, 'local_g3_7')
// (10, 19, 'lutff_5/in_3')
// (10, 19, 'lutff_7/out')
// (10, 20, 'neigh_op_bot_7')
// (11, 18, 'neigh_op_tnl_7')
// (11, 19, 'neigh_op_lft_7')
// (11, 20, 'neigh_op_bnl_7')

wire n1378;
// (9, 19, 'lutff_0/cout')
// (9, 19, 'lutff_1/in_3')

wire n1379;
// (9, 19, 'neigh_op_tnr_1')
// (9, 20, 'neigh_op_rgt_1')
// (9, 21, 'neigh_op_bnr_1')
// (10, 19, 'neigh_op_top_1')
// (10, 20, 'local_g1_1')
// (10, 20, 'lutff_1/out')
// (10, 20, 'lutff_6/in_2')
// (10, 21, 'neigh_op_bot_1')
// (11, 19, 'neigh_op_tnl_1')
// (11, 20, 'neigh_op_lft_1')
// (11, 21, 'neigh_op_bnl_1')

reg n1380 = 0;
// (9, 19, 'neigh_op_tnr_5')
// (9, 20, 'neigh_op_rgt_5')
// (9, 21, 'neigh_op_bnr_5')
// (10, 19, 'neigh_op_top_5')
// (10, 20, 'local_g3_5')
// (10, 20, 'lutff_5/in_3')
// (10, 20, 'lutff_5/out')
// (10, 21, 'neigh_op_bot_5')
// (11, 19, 'local_g3_5')
// (11, 19, 'lutff_7/in_1')
// (11, 19, 'neigh_op_tnl_5')
// (11, 20, 'local_g0_5')
// (11, 20, 'local_g1_5')
// (11, 20, 'lutff_1/in_1')
// (11, 20, 'lutff_6/in_3')
// (11, 20, 'neigh_op_lft_5')
// (11, 21, 'neigh_op_bnl_5')

wire n1381;
// (9, 19, 'neigh_op_tnr_6')
// (9, 20, 'neigh_op_rgt_6')
// (9, 21, 'neigh_op_bnr_6')
// (10, 19, 'local_g0_6')
// (10, 19, 'lutff_3/in_3')
// (10, 19, 'neigh_op_top_6')
// (10, 20, 'lutff_6/out')
// (10, 21, 'neigh_op_bot_6')
// (11, 19, 'neigh_op_tnl_6')
// (11, 20, 'neigh_op_lft_6')
// (11, 21, 'neigh_op_bnl_6')

wire n1382;
// (9, 20, 'lutff_1/cout')
// (9, 20, 'lutff_2/in_3')

wire n1383;
// (9, 20, 'lutff_2/cout')
// (9, 20, 'lutff_3/in_3')

wire n1384;
// (9, 20, 'lutff_3/cout')
// (9, 20, 'lutff_4/in_3')

wire n1385;
// (9, 20, 'lutff_4/cout')
// (9, 20, 'lutff_5/in_3')

wire n1386;
// (9, 20, 'lutff_5/cout')
// (9, 20, 'lutff_6/in_3')

wire n1387;
// (9, 20, 'lutff_6/cout')
// (9, 20, 'lutff_7/in_3')

wire n1388;
// (9, 20, 'lutff_7/cout')
// (9, 21, 'carry_in')
// (9, 21, 'carry_in_mux')
// (9, 21, 'lutff_0/in_3')

wire n1389;
// (9, 20, 'neigh_op_tnr_4')
// (9, 21, 'neigh_op_rgt_4')
// (9, 22, 'neigh_op_bnr_4')
// (10, 20, 'neigh_op_top_4')
// (10, 21, 'local_g3_4')
// (10, 21, 'lutff_4/out')
// (10, 21, 'lutff_7/in_2')
// (10, 22, 'neigh_op_bot_4')
// (11, 20, 'neigh_op_tnl_4')
// (11, 21, 'neigh_op_lft_4')
// (11, 22, 'neigh_op_bnl_4')

wire n1390;
// (9, 20, 'sp12_h_r_0')
// (10, 19, 'neigh_op_tnr_6')
// (10, 20, 'local_g1_3')
// (10, 20, 'lutff_global/cen')
// (10, 20, 'neigh_op_rgt_6')
// (10, 20, 'sp12_h_r_3')
// (10, 21, 'neigh_op_bnr_6')
// (11, 19, 'neigh_op_top_6')
// (11, 20, 'lutff_6/out')
// (11, 20, 'sp12_h_r_4')
// (11, 21, 'neigh_op_bot_6')
// (12, 19, 'neigh_op_tnl_6')
// (12, 20, 'neigh_op_lft_6')
// (12, 20, 'sp12_h_r_7')
// (12, 21, 'neigh_op_bnl_6')
// (13, 20, 'sp12_h_r_8')
// (14, 20, 'sp12_h_r_11')
// (15, 20, 'sp12_h_r_12')
// (16, 20, 'sp12_h_r_15')
// (17, 20, 'sp12_h_r_16')
// (18, 20, 'sp12_h_r_19')
// (19, 20, 'sp12_h_r_20')
// (20, 20, 'sp12_h_r_23')
// (21, 20, 'sp12_h_l_23')

reg n1391 = 0;
// (9, 21, 'sp4_h_r_7')
// (10, 21, 'local_g1_2')
// (10, 21, 'lutff_4/in_3')
// (10, 21, 'sp4_h_r_18')
// (11, 20, 'neigh_op_tnr_5')
// (11, 21, 'local_g3_5')
// (11, 21, 'lutff_1/in_3')
// (11, 21, 'lutff_6/in_0')
// (11, 21, 'neigh_op_rgt_5')
// (11, 21, 'sp4_h_r_31')
// (11, 22, 'neigh_op_bnr_5')
// (12, 20, 'neigh_op_top_5')
// (12, 21, 'lutff_5/out')
// (12, 21, 'sp4_h_r_42')
// (12, 22, 'neigh_op_bot_5')
// (13, 20, 'neigh_op_tnl_5')
// (13, 21, 'neigh_op_lft_5')
// (13, 21, 'sp4_h_l_42')
// (13, 22, 'neigh_op_bnl_5')

wire n1392;
// (9, 22, 'lutff_1/cout')
// (9, 22, 'lutff_2/in_3')

wire n1393;
// (9, 22, 'lutff_2/cout')
// (9, 22, 'lutff_3/in_3')

wire n1394;
// (9, 22, 'lutff_3/cout')
// (9, 22, 'lutff_4/in_3')

wire n1395;
// (9, 22, 'lutff_4/cout')
// (9, 22, 'lutff_5/in_3')

reg n1396 = 0;
// (10, 1, 'local_g2_4')
// (10, 1, 'lutff_0/in_2')
// (10, 1, 'neigh_op_tnr_4')
// (10, 2, 'local_g3_4')
// (10, 2, 'lutff_3/in_2')
// (10, 2, 'neigh_op_rgt_4')
// (10, 3, 'neigh_op_bnr_4')
// (11, 1, 'neigh_op_top_4')
// (11, 2, 'lutff_4/out')
// (11, 3, 'neigh_op_bot_4')
// (12, 1, 'neigh_op_tnl_4')
// (12, 2, 'neigh_op_lft_4')
// (12, 3, 'neigh_op_bnl_4')

wire n1397;
// (10, 1, 'neigh_op_tnr_0')
// (10, 2, 'neigh_op_rgt_0')
// (10, 3, 'neigh_op_bnr_0')
// (11, 1, 'neigh_op_top_0')
// (11, 1, 'sp4_r_v_b_44')
// (11, 2, 'lutff_0/out')
// (11, 2, 'sp4_r_v_b_33')
// (11, 3, 'neigh_op_bot_0')
// (11, 3, 'sp4_r_v_b_20')
// (11, 4, 'sp4_r_v_b_9')
// (12, 0, 'span4_vert_44')
// (12, 1, 'neigh_op_tnl_0')
// (12, 1, 'sp4_v_b_44')
// (12, 2, 'neigh_op_lft_0')
// (12, 2, 'sp4_v_b_33')
// (12, 3, 'neigh_op_bnl_0')
// (12, 3, 'sp4_v_b_20')
// (12, 4, 'local_g0_1')
// (12, 4, 'lutff_6/in_1')
// (12, 4, 'sp4_v_b_9')

reg n1398 = 0;
// (10, 1, 'neigh_op_tnr_1')
// (10, 2, 'local_g3_1')
// (10, 2, 'lutff_2/in_2')
// (10, 2, 'neigh_op_rgt_1')
// (10, 3, 'neigh_op_bnr_1')
// (11, 1, 'neigh_op_top_1')
// (11, 2, 'local_g0_1')
// (11, 2, 'lutff_1/out')
// (11, 2, 'lutff_2/in_1')
// (11, 3, 'neigh_op_bot_1')
// (12, 1, 'neigh_op_tnl_1')
// (12, 2, 'neigh_op_lft_1')
// (12, 3, 'neigh_op_bnl_1')

wire n1399;
// (10, 1, 'neigh_op_tnr_2')
// (10, 2, 'neigh_op_rgt_2')
// (10, 3, 'neigh_op_bnr_2')
// (11, 1, 'neigh_op_top_2')
// (11, 2, 'lutff_2/out')
// (11, 3, 'local_g1_2')
// (11, 3, 'lutff_5/in_0')
// (11, 3, 'neigh_op_bot_2')
// (12, 1, 'neigh_op_tnl_2')
// (12, 2, 'neigh_op_lft_2')
// (12, 3, 'neigh_op_bnl_2')

wire n1400;
// (10, 1, 'neigh_op_tnr_3')
// (10, 2, 'local_g3_3')
// (10, 2, 'lutff_1/in_3')
// (10, 2, 'neigh_op_rgt_3')
// (10, 3, 'neigh_op_bnr_3')
// (11, 1, 'neigh_op_top_3')
// (11, 2, 'lutff_3/out')
// (11, 3, 'neigh_op_bot_3')
// (12, 1, 'neigh_op_tnl_3')
// (12, 2, 'neigh_op_lft_3')
// (12, 3, 'neigh_op_bnl_3')

reg n1401 = 0;
// (10, 1, 'neigh_op_tnr_5')
// (10, 2, 'local_g2_5')
// (10, 2, 'lutff_2/in_3')
// (10, 2, 'neigh_op_rgt_5')
// (10, 3, 'neigh_op_bnr_5')
// (11, 1, 'neigh_op_top_5')
// (11, 2, 'lutff_5/out')
// (11, 3, 'local_g1_5')
// (11, 3, 'lutff_6/in_2')
// (11, 3, 'neigh_op_bot_5')
// (12, 1, 'neigh_op_tnl_5')
// (12, 2, 'neigh_op_lft_5')
// (12, 3, 'neigh_op_bnl_5')

wire n1402;
// (10, 1, 'sp4_r_v_b_32')
// (10, 2, 'neigh_op_tnr_4')
// (10, 2, 'sp4_r_v_b_21')
// (10, 3, 'neigh_op_rgt_4')
// (10, 3, 'sp4_r_v_b_8')
// (10, 4, 'neigh_op_bnr_4')
// (11, 0, 'span4_vert_32')
// (11, 1, 'local_g3_0')
// (11, 1, 'lutff_1/in_2')
// (11, 1, 'sp4_r_v_b_33')
// (11, 1, 'sp4_v_b_32')
// (11, 2, 'neigh_op_top_4')
// (11, 2, 'sp4_r_v_b_20')
// (11, 2, 'sp4_r_v_b_36')
// (11, 2, 'sp4_v_b_21')
// (11, 3, 'lutff_4/out')
// (11, 3, 'sp4_r_v_b_25')
// (11, 3, 'sp4_r_v_b_9')
// (11, 3, 'sp4_v_b_8')
// (11, 4, 'neigh_op_bot_4')
// (11, 4, 'sp4_r_v_b_12')
// (11, 5, 'sp4_r_v_b_1')
// (12, 0, 'span4_vert_33')
// (12, 1, 'local_g2_1')
// (12, 1, 'lutff_1/in_2')
// (12, 1, 'sp4_h_r_6')
// (12, 1, 'sp4_v_b_33')
// (12, 1, 'sp4_v_t_36')
// (12, 2, 'neigh_op_tnl_4')
// (12, 2, 'sp4_v_b_20')
// (12, 2, 'sp4_v_b_36')
// (12, 3, 'local_g1_4')
// (12, 3, 'lutff_0/in_1')
// (12, 3, 'neigh_op_lft_4')
// (12, 3, 'sp4_v_b_25')
// (12, 3, 'sp4_v_b_9')
// (12, 4, 'neigh_op_bnl_4')
// (12, 4, 'sp4_v_b_12')
// (12, 5, 'sp4_v_b_1')
// (13, 1, 'local_g1_3')
// (13, 1, 'lutff_1/in_1')
// (13, 1, 'sp4_h_r_19')
// (14, 1, 'sp4_h_r_30')
// (15, 1, 'sp4_h_r_43')
// (16, 1, 'sp4_h_l_43')

reg n1403 = 0;
// (10, 2, 'neigh_op_tnr_1')
// (10, 3, 'local_g2_1')
// (10, 3, 'local_g3_1')
// (10, 3, 'lutff_2/in_2')
// (10, 3, 'lutff_4/in_3')
// (10, 3, 'neigh_op_rgt_1')
// (10, 4, 'neigh_op_bnr_1')
// (11, 2, 'neigh_op_top_1')
// (11, 3, 'lutff_1/out')
// (11, 4, 'neigh_op_bot_1')
// (12, 2, 'neigh_op_tnl_1')
// (12, 3, 'neigh_op_lft_1')
// (12, 4, 'neigh_op_bnl_1')

wire n1404;
// (10, 2, 'neigh_op_tnr_2')
// (10, 3, 'local_g2_2')
// (10, 3, 'lutff_3/in_3')
// (10, 3, 'neigh_op_rgt_2')
// (10, 4, 'neigh_op_bnr_2')
// (11, 2, 'neigh_op_top_2')
// (11, 3, 'lutff_2/out')
// (11, 4, 'neigh_op_bot_2')
// (12, 2, 'neigh_op_tnl_2')
// (12, 3, 'neigh_op_lft_2')
// (12, 4, 'neigh_op_bnl_2')

wire n1405;
// (10, 2, 'neigh_op_tnr_5')
// (10, 3, 'neigh_op_rgt_5')
// (10, 4, 'local_g1_5')
// (10, 4, 'lutff_6/in_2')
// (10, 4, 'neigh_op_bnr_5')
// (11, 2, 'neigh_op_top_5')
// (11, 3, 'lutff_5/out')
// (11, 4, 'neigh_op_bot_5')
// (12, 2, 'neigh_op_tnl_5')
// (12, 3, 'neigh_op_lft_5')
// (12, 4, 'neigh_op_bnl_5')

wire n1406;
// (10, 2, 'neigh_op_tnr_6')
// (10, 3, 'neigh_op_rgt_6')
// (10, 4, 'neigh_op_bnr_6')
// (11, 2, 'neigh_op_top_6')
// (11, 3, 'lutff_6/out')
// (11, 4, 'local_g0_6')
// (11, 4, 'lutff_1/in_3')
// (11, 4, 'neigh_op_bot_6')
// (12, 2, 'neigh_op_tnl_6')
// (12, 3, 'neigh_op_lft_6')
// (12, 4, 'neigh_op_bnl_6')

reg n1407 = 0;
// (10, 2, 'neigh_op_tnr_7')
// (10, 3, 'local_g2_7')
// (10, 3, 'lutff_1/in_2')
// (10, 3, 'neigh_op_rgt_7')
// (10, 4, 'neigh_op_bnr_7')
// (11, 2, 'neigh_op_top_7')
// (11, 3, 'local_g1_7')
// (11, 3, 'lutff_5/in_3')
// (11, 3, 'lutff_7/out')
// (11, 4, 'neigh_op_bot_7')
// (12, 2, 'neigh_op_tnl_7')
// (12, 3, 'neigh_op_lft_7')
// (12, 4, 'neigh_op_bnl_7')

wire n1408;
// (10, 3, 'local_g0_6')
// (10, 3, 'lutff_7/in_1')
// (10, 3, 'sp4_h_r_6')
// (11, 3, 'sp4_h_r_19')
// (12, 3, 'sp4_h_r_30')
// (13, 1, 'neigh_op_tnr_6')
// (13, 1, 'sp4_r_v_b_25')
// (13, 2, 'neigh_op_rgt_6')
// (13, 2, 'sp4_r_v_b_12')
// (13, 3, 'neigh_op_bnr_6')
// (13, 3, 'sp4_h_r_43')
// (13, 3, 'sp4_r_v_b_1')
// (14, 0, 'span4_vert_25')
// (14, 1, 'neigh_op_top_6')
// (14, 1, 'sp4_v_b_25')
// (14, 2, 'lutff_6/out')
// (14, 2, 'sp4_v_b_12')
// (14, 3, 'neigh_op_bot_6')
// (14, 3, 'sp4_h_l_43')
// (14, 3, 'sp4_v_b_1')
// (15, 1, 'neigh_op_tnl_6')
// (15, 2, 'local_g0_6')
// (15, 2, 'lutff_7/in_1')
// (15, 2, 'neigh_op_lft_6')
// (15, 3, 'neigh_op_bnl_6')

reg n1409 = 0;
// (10, 3, 'local_g2_4')
// (10, 3, 'lutff_4/in_2')
// (10, 3, 'neigh_op_tnr_4')
// (10, 4, 'neigh_op_rgt_4')
// (10, 5, 'neigh_op_bnr_4')
// (11, 3, 'local_g0_4')
// (11, 3, 'lutff_2/in_0')
// (11, 3, 'neigh_op_top_4')
// (11, 4, 'lutff_4/out')
// (11, 5, 'neigh_op_bot_4')
// (12, 3, 'neigh_op_tnl_4')
// (12, 4, 'neigh_op_lft_4')
// (12, 5, 'neigh_op_bnl_4')

wire n1410;
// (10, 3, 'local_g3_2')
// (10, 3, 'lutff_2/in_1')
// (10, 3, 'lutff_6/in_1')
// (10, 3, 'lutff_7/in_2')
// (10, 3, 'neigh_op_tnr_2')
// (10, 4, 'local_g2_2')
// (10, 4, 'lutff_3/in_1')
// (10, 4, 'neigh_op_rgt_2')
// (10, 5, 'local_g1_2')
// (10, 5, 'lutff_5/in_0')
// (10, 5, 'neigh_op_bnr_2')
// (11, 2, 'sp4_r_v_b_45')
// (11, 3, 'local_g0_2')
// (11, 3, 'lutff_2/in_2')
// (11, 3, 'lutff_5/in_1')
// (11, 3, 'neigh_op_top_2')
// (11, 3, 'sp4_r_v_b_32')
// (11, 4, 'local_g1_2')
// (11, 4, 'lutff_2/out')
// (11, 4, 'lutff_5/in_0')
// (11, 4, 'sp4_h_r_4')
// (11, 4, 'sp4_r_v_b_21')
// (11, 4, 'sp4_r_v_b_37')
// (11, 5, 'neigh_op_bot_2')
// (11, 5, 'sp4_r_v_b_24')
// (11, 5, 'sp4_r_v_b_8')
// (11, 6, 'sp4_r_v_b_13')
// (11, 7, 'sp4_r_v_b_0')
// (12, 1, 'sp4_v_t_45')
// (12, 2, 'sp4_v_b_45')
// (12, 3, 'neigh_op_tnl_2')
// (12, 3, 'sp4_v_b_32')
// (12, 3, 'sp4_v_t_37')
// (12, 4, 'local_g0_2')
// (12, 4, 'lutff_5/in_1')
// (12, 4, 'neigh_op_lft_2')
// (12, 4, 'sp4_h_r_17')
// (12, 4, 'sp4_v_b_21')
// (12, 4, 'sp4_v_b_37')
// (12, 5, 'neigh_op_bnl_2')
// (12, 5, 'sp4_h_r_8')
// (12, 5, 'sp4_v_b_24')
// (12, 5, 'sp4_v_b_8')
// (12, 6, 'local_g1_5')
// (12, 6, 'lutff_3/in_3')
// (12, 6, 'sp4_v_b_13')
// (12, 7, 'local_g1_0')
// (12, 7, 'lutff_7/in_0')
// (12, 7, 'sp4_h_r_6')
// (12, 7, 'sp4_v_b_0')
// (13, 4, 'sp4_h_r_28')
// (13, 5, 'local_g0_5')
// (13, 5, 'local_g1_5')
// (13, 5, 'lutff_2/in_1')
// (13, 5, 'lutff_4/in_0')
// (13, 5, 'sp4_h_r_21')
// (13, 7, 'sp4_h_r_19')
// (14, 4, 'local_g2_1')
// (14, 4, 'lutff_2/in_1')
// (14, 4, 'lutff_5/in_0')
// (14, 4, 'sp4_h_r_41')
// (14, 5, 'local_g2_0')
// (14, 5, 'lutff_1/in_3')
// (14, 5, 'sp4_h_r_32')
// (14, 7, 'local_g3_6')
// (14, 7, 'lutff_5/in_2')
// (14, 7, 'sp4_h_r_30')
// (15, 4, 'sp4_h_l_41')
// (15, 5, 'sp4_h_r_45')
// (15, 7, 'sp4_h_r_43')
// (16, 5, 'sp4_h_l_45')
// (16, 7, 'sp4_h_l_43')

wire n1411;
// (10, 3, 'neigh_op_tnr_1')
// (10, 4, 'neigh_op_rgt_1')
// (10, 5, 'local_g0_1')
// (10, 5, 'lutff_5/in_2')
// (10, 5, 'neigh_op_bnr_1')
// (11, 3, 'neigh_op_top_1')
// (11, 4, 'lutff_1/out')
// (11, 5, 'neigh_op_bot_1')
// (12, 3, 'neigh_op_tnl_1')
// (12, 4, 'neigh_op_lft_1')
// (12, 5, 'neigh_op_bnl_1')

wire n1412;
// (10, 3, 'neigh_op_tnr_3')
// (10, 4, 'neigh_op_rgt_3')
// (10, 4, 'sp4_r_v_b_38')
// (10, 5, 'neigh_op_bnr_3')
// (10, 5, 'sp4_r_v_b_27')
// (10, 6, 'sp4_r_v_b_14')
// (10, 7, 'sp4_r_v_b_3')
// (10, 8, 'sp4_r_v_b_38')
// (10, 9, 'sp4_r_v_b_27')
// (10, 10, 'sp4_r_v_b_14')
// (10, 11, 'sp4_r_v_b_3')
// (11, 3, 'local_g0_3')
// (11, 3, 'lutff_3/in_0')
// (11, 3, 'neigh_op_top_3')
// (11, 3, 'sp4_v_t_38')
// (11, 4, 'local_g0_3')
// (11, 4, 'lutff_3/out')
// (11, 4, 'lutff_7/in_0')
// (11, 4, 'sp4_v_b_38')
// (11, 5, 'neigh_op_bot_3')
// (11, 5, 'sp4_v_b_27')
// (11, 6, 'sp4_v_b_14')
// (11, 7, 'sp4_v_b_3')
// (11, 7, 'sp4_v_t_38')
// (11, 8, 'sp4_v_b_38')
// (11, 9, 'sp4_v_b_27')
// (11, 10, 'local_g1_6')
// (11, 10, 'lutff_2/in_3')
// (11, 10, 'sp4_v_b_14')
// (11, 11, 'sp4_v_b_3')
// (12, 3, 'neigh_op_tnl_3')
// (12, 4, 'neigh_op_lft_3')
// (12, 5, 'neigh_op_bnl_3')

wire n1413;
// (10, 3, 'neigh_op_tnr_5')
// (10, 4, 'local_g3_5')
// (10, 4, 'lutff_5/in_3')
// (10, 4, 'neigh_op_rgt_5')
// (10, 5, 'neigh_op_bnr_5')
// (11, 3, 'neigh_op_top_5')
// (11, 4, 'lutff_5/out')
// (11, 5, 'neigh_op_bot_5')
// (12, 3, 'neigh_op_tnl_5')
// (12, 4, 'neigh_op_lft_5')
// (12, 5, 'neigh_op_bnl_5')

reg n1414 = 0;
// (10, 3, 'neigh_op_tnr_6')
// (10, 4, 'local_g3_6')
// (10, 4, 'lutff_4/in_1')
// (10, 4, 'neigh_op_rgt_6')
// (10, 5, 'neigh_op_bnr_6')
// (11, 3, 'neigh_op_top_6')
// (11, 4, 'local_g2_6')
// (11, 4, 'lutff_5/in_3')
// (11, 4, 'lutff_6/out')
// (11, 5, 'neigh_op_bot_6')
// (12, 3, 'neigh_op_tnl_6')
// (12, 4, 'neigh_op_lft_6')
// (12, 5, 'neigh_op_bnl_6')

wire n1415;
// (10, 3, 'neigh_op_tnr_7')
// (10, 4, 'neigh_op_rgt_7')
// (10, 5, 'neigh_op_bnr_7')
// (11, 3, 'neigh_op_top_7')
// (11, 4, 'local_g3_7')
// (11, 4, 'lutff_0/in_2')
// (11, 4, 'lutff_7/out')
// (11, 5, 'neigh_op_bot_7')
// (12, 3, 'neigh_op_tnl_7')
// (12, 4, 'neigh_op_lft_7')
// (12, 5, 'neigh_op_bnl_7')

reg n1416 = 0;
// (10, 3, 'sp4_r_v_b_40')
// (10, 4, 'sp4_r_v_b_29')
// (10, 5, 'sp4_r_v_b_16')
// (10, 6, 'sp4_r_v_b_5')
// (11, 2, 'sp4_v_t_40')
// (11, 3, 'local_g2_0')
// (11, 3, 'lutff_4/in_0')
// (11, 3, 'sp4_v_b_40')
// (11, 4, 'local_g2_5')
// (11, 4, 'lutff_3/in_0')
// (11, 4, 'sp4_v_b_29')
// (11, 5, 'local_g1_0')
// (11, 5, 'lutff_1/in_2')
// (11, 5, 'lutff_7/in_0')
// (11, 5, 'sp4_v_b_16')
// (11, 6, 'local_g0_3')
// (11, 6, 'lutff_2/in_3')
// (11, 6, 'sp4_h_r_0')
// (11, 6, 'sp4_h_r_3')
// (11, 6, 'sp4_v_b_5')
// (12, 3, 'sp4_r_v_b_36')
// (12, 4, 'local_g1_1')
// (12, 4, 'lutff_7/in_1')
// (12, 4, 'sp4_r_v_b_25')
// (12, 5, 'sp4_r_v_b_12')
// (12, 6, 'sp4_h_r_13')
// (12, 6, 'sp4_h_r_14')
// (12, 6, 'sp4_r_v_b_1')
// (12, 11, 'sp4_r_v_b_42')
// (12, 12, 'sp4_r_v_b_31')
// (12, 13, 'sp4_r_v_b_18')
// (12, 14, 'sp4_r_v_b_7')
// (13, 2, 'sp4_v_t_36')
// (13, 3, 'sp4_v_b_36')
// (13, 4, 'sp4_v_b_25')
// (13, 5, 'sp4_v_b_12')
// (13, 6, 'sp4_h_r_24')
// (13, 6, 'sp4_h_r_27')
// (13, 6, 'sp4_h_r_8')
// (13, 6, 'sp4_v_b_1')
// (13, 10, 'sp4_h_r_1')
// (13, 10, 'sp4_v_t_42')
// (13, 11, 'sp4_v_b_42')
// (13, 12, 'sp4_v_b_31')
// (13, 13, 'sp4_v_b_18')
// (13, 14, 'local_g0_7')
// (13, 14, 'lutff_5/in_2')
// (13, 14, 'lutff_7/in_2')
// (13, 14, 'sp4_v_b_7')
// (14, 3, 'sp4_r_v_b_37')
// (14, 4, 'sp4_r_v_b_24')
// (14, 5, 'local_g3_0')
// (14, 5, 'lutff_2/in_1')
// (14, 5, 'lutff_5/in_2')
// (14, 5, 'neigh_op_tnr_0')
// (14, 5, 'sp4_r_v_b_13')
// (14, 6, 'neigh_op_rgt_0')
// (14, 6, 'sp4_h_r_21')
// (14, 6, 'sp4_h_r_37')
// (14, 6, 'sp4_h_r_38')
// (14, 6, 'sp4_r_v_b_0')
// (14, 7, 'neigh_op_bnr_0')
// (14, 10, 'sp4_h_r_12')
// (15, 2, 'sp4_v_t_37')
// (15, 3, 'local_g2_5')
// (15, 3, 'lutff_3/in_0')
// (15, 3, 'sp4_v_b_37')
// (15, 4, 'sp4_v_b_24')
// (15, 5, 'local_g0_0')
// (15, 5, 'lutff_5/in_1')
// (15, 5, 'lutff_7/in_1')
// (15, 5, 'neigh_op_top_0')
// (15, 5, 'sp4_v_b_13')
// (15, 6, 'local_g3_0')
// (15, 6, 'lutff_0/in_3')
// (15, 6, 'lutff_0/out')
// (15, 6, 'sp4_h_l_37')
// (15, 6, 'sp4_h_l_38')
// (15, 6, 'sp4_h_r_0')
// (15, 6, 'sp4_h_r_32')
// (15, 6, 'sp4_v_b_0')
// (15, 7, 'neigh_op_bot_0')
// (15, 10, 'sp4_h_r_25')
// (16, 5, 'neigh_op_tnl_0')
// (16, 6, 'neigh_op_lft_0')
// (16, 6, 'sp4_h_r_13')
// (16, 6, 'sp4_h_r_45')
// (16, 7, 'neigh_op_bnl_0')
// (16, 7, 'sp4_r_v_b_45')
// (16, 8, 'sp4_r_v_b_32')
// (16, 9, 'sp4_r_v_b_21')
// (16, 10, 'sp4_h_r_36')
// (16, 10, 'sp4_r_v_b_8')
// (17, 6, 'local_g3_0')
// (17, 6, 'lutff_2/in_1')
// (17, 6, 'sp4_h_l_45')
// (17, 6, 'sp4_h_r_24')
// (17, 6, 'sp4_v_t_45')
// (17, 7, 'sp4_v_b_45')
// (17, 8, 'sp4_v_b_32')
// (17, 9, 'sp4_v_b_21')
// (17, 10, 'sp4_h_l_36')
// (17, 10, 'sp4_v_b_8')
// (18, 6, 'sp4_h_r_37')
// (19, 6, 'sp4_h_l_37')

wire n1417;
// (10, 3, 'sp4_r_v_b_45')
// (10, 4, 'sp4_r_v_b_32')
// (10, 5, 'sp4_r_v_b_21')
// (10, 6, 'sp4_r_v_b_8')
// (11, 2, 'sp4_h_r_2')
// (11, 2, 'sp4_v_t_45')
// (11, 3, 'local_g2_5')
// (11, 3, 'lutff_2/in_3')
// (11, 3, 'sp4_v_b_45')
// (11, 4, 'sp4_v_b_32')
// (11, 5, 'sp4_v_b_21')
// (11, 6, 'sp4_v_b_8')
// (12, 1, 'neigh_op_tnr_5')
// (12, 2, 'neigh_op_rgt_5')
// (12, 2, 'sp4_h_r_15')
// (12, 3, 'neigh_op_bnr_5')
// (13, 1, 'neigh_op_top_5')
// (13, 2, 'lutff_5/out')
// (13, 2, 'sp4_h_r_26')
// (13, 3, 'local_g0_5')
// (13, 3, 'lutff_1/in_2')
// (13, 3, 'neigh_op_bot_5')
// (14, 1, 'neigh_op_tnl_5')
// (14, 2, 'neigh_op_lft_5')
// (14, 2, 'sp4_h_r_39')
// (14, 3, 'neigh_op_bnl_5')
// (15, 2, 'sp4_h_l_39')

reg n1418 = 0;
// (10, 3, 'sp4_r_v_b_46')
// (10, 4, 'neigh_op_tnr_3')
// (10, 4, 'sp4_r_v_b_35')
// (10, 5, 'neigh_op_rgt_3')
// (10, 5, 'sp4_r_v_b_22')
// (10, 6, 'neigh_op_bnr_3')
// (10, 6, 'sp4_r_v_b_11')
// (11, 2, 'sp4_v_t_46')
// (11, 3, 'sp4_v_b_46')
// (11, 4, 'neigh_op_top_3')
// (11, 4, 'sp4_v_b_35')
// (11, 5, 'lutff_3/out')
// (11, 5, 'sp4_v_b_22')
// (11, 6, 'neigh_op_bot_3')
// (11, 6, 'sp4_h_r_11')
// (11, 6, 'sp4_v_b_11')
// (12, 4, 'neigh_op_tnl_3')
// (12, 5, 'neigh_op_lft_3')
// (12, 6, 'local_g3_3')
// (12, 6, 'lutff_3/in_1')
// (12, 6, 'lutff_6/in_0')
// (12, 6, 'neigh_op_bnl_3')
// (12, 6, 'sp4_h_r_22')
// (13, 6, 'local_g2_3')
// (13, 6, 'lutff_0/in_1')
// (13, 6, 'sp4_h_r_35')
// (14, 6, 'sp4_h_r_46')
// (15, 6, 'sp4_h_l_46')

wire n1419;
// (10, 4, 'neigh_op_tnr_2')
// (10, 5, 'neigh_op_rgt_2')
// (10, 5, 'sp4_r_v_b_36')
// (10, 6, 'neigh_op_bnr_2')
// (10, 6, 'sp4_r_v_b_25')
// (10, 7, 'sp4_r_v_b_12')
// (10, 8, 'sp4_r_v_b_1')
// (11, 4, 'neigh_op_top_2')
// (11, 4, 'sp4_v_t_36')
// (11, 5, 'lutff_2/out')
// (11, 5, 'sp4_v_b_36')
// (11, 6, 'neigh_op_bot_2')
// (11, 6, 'sp4_v_b_25')
// (11, 7, 'local_g1_4')
// (11, 7, 'lutff_5/in_0')
// (11, 7, 'lutff_6/in_1')
// (11, 7, 'sp4_v_b_12')
// (11, 8, 'sp4_v_b_1')
// (12, 4, 'local_g2_2')
// (12, 4, 'lutff_0/in_0')
// (12, 4, 'lutff_3/in_1')
// (12, 4, 'neigh_op_tnl_2')
// (12, 5, 'neigh_op_lft_2')
// (12, 6, 'neigh_op_bnl_2')

wire n1420;
// (10, 4, 'neigh_op_tnr_5')
// (10, 4, 'sp4_r_v_b_39')
// (10, 5, 'neigh_op_rgt_5')
// (10, 5, 'sp4_r_v_b_26')
// (10, 6, 'neigh_op_bnr_5')
// (10, 6, 'sp4_r_v_b_15')
// (10, 7, 'sp4_r_v_b_2')
// (11, 3, 'sp4_h_r_2')
// (11, 3, 'sp4_v_t_39')
// (11, 4, 'neigh_op_top_5')
// (11, 4, 'sp4_v_b_39')
// (11, 5, 'lutff_5/out')
// (11, 5, 'sp4_v_b_26')
// (11, 6, 'neigh_op_bot_5')
// (11, 6, 'sp4_v_b_15')
// (11, 7, 'sp4_v_b_2')
// (12, 3, 'sp4_h_r_15')
// (12, 4, 'neigh_op_tnl_5')
// (12, 5, 'neigh_op_lft_5')
// (12, 6, 'neigh_op_bnl_5')
// (13, 3, 'local_g2_2')
// (13, 3, 'lutff_5/in_3')
// (13, 3, 'sp4_h_r_26')
// (14, 3, 'sp4_h_r_39')
// (15, 3, 'sp4_h_l_39')

wire n1421;
// (10, 4, 'neigh_op_tnr_7')
// (10, 5, 'neigh_op_rgt_7')
// (10, 6, 'neigh_op_bnr_7')
// (11, 4, 'neigh_op_top_7')
// (11, 5, 'local_g0_7')
// (11, 5, 'lutff_4/in_1')
// (11, 5, 'lutff_7/out')
// (11, 6, 'neigh_op_bot_7')
// (12, 4, 'neigh_op_tnl_7')
// (12, 5, 'neigh_op_lft_7')
// (12, 6, 'neigh_op_bnl_7')

wire n1422;
// (10, 4, 'sp4_h_r_8')
// (11, 3, 'neigh_op_tnr_0')
// (11, 4, 'neigh_op_rgt_0')
// (11, 4, 'sp4_h_r_21')
// (11, 5, 'local_g0_0')
// (11, 5, 'lutff_6/in_2')
// (11, 5, 'neigh_op_bnr_0')
// (12, 3, 'neigh_op_top_0')
// (12, 4, 'lutff_0/out')
// (12, 4, 'sp4_h_r_0')
// (12, 4, 'sp4_h_r_32')
// (12, 5, 'neigh_op_bot_0')
// (13, 1, 'sp4_r_v_b_45')
// (13, 2, 'sp4_r_v_b_32')
// (13, 3, 'local_g2_0')
// (13, 3, 'lutff_3/in_1')
// (13, 3, 'neigh_op_tnl_0')
// (13, 3, 'sp4_r_v_b_21')
// (13, 4, 'local_g0_0')
// (13, 4, 'lutff_4/in_0')
// (13, 4, 'lutff_5/in_1')
// (13, 4, 'lutff_6/in_2')
// (13, 4, 'lutff_7/in_1')
// (13, 4, 'neigh_op_lft_0')
// (13, 4, 'sp4_h_r_13')
// (13, 4, 'sp4_h_r_45')
// (13, 4, 'sp4_r_v_b_8')
// (13, 5, 'neigh_op_bnl_0')
// (14, 0, 'span4_vert_45')
// (14, 1, 'sp4_v_b_45')
// (14, 2, 'sp4_v_b_32')
// (14, 3, 'local_g1_5')
// (14, 3, 'lutff_5/in_3')
// (14, 3, 'sp4_v_b_21')
// (14, 4, 'local_g2_0')
// (14, 4, 'lutff_3/in_3')
// (14, 4, 'sp4_h_l_45')
// (14, 4, 'sp4_h_r_24')
// (14, 4, 'sp4_v_b_8')
// (15, 4, 'local_g2_5')
// (15, 4, 'lutff_7/in_0')
// (15, 4, 'sp4_h_r_37')
// (16, 4, 'sp4_h_l_37')

wire n1423;
// (10, 4, 'sp4_h_r_9')
// (11, 4, 'sp4_h_r_20')
// (12, 1, 'neigh_op_tnr_0')
// (12, 2, 'neigh_op_rgt_0')
// (12, 3, 'neigh_op_bnr_0')
// (12, 4, 'local_g2_1')
// (12, 4, 'lutff_3/in_2')
// (12, 4, 'sp4_h_r_33')
// (13, 1, 'neigh_op_top_0')
// (13, 1, 'sp4_r_v_b_44')
// (13, 2, 'lutff_0/out')
// (13, 2, 'sp4_r_v_b_33')
// (13, 3, 'neigh_op_bot_0')
// (13, 3, 'sp4_r_v_b_20')
// (13, 4, 'sp4_h_r_44')
// (13, 4, 'sp4_r_v_b_9')
// (14, 0, 'span4_vert_44')
// (14, 1, 'neigh_op_tnl_0')
// (14, 1, 'sp4_v_b_44')
// (14, 2, 'neigh_op_lft_0')
// (14, 2, 'sp4_v_b_33')
// (14, 3, 'neigh_op_bnl_0')
// (14, 3, 'sp4_v_b_20')
// (14, 4, 'sp4_h_l_44')
// (14, 4, 'sp4_v_b_9')

wire n1424;
// (10, 5, 'local_g3_2')
// (10, 5, 'lutff_1/in_2')
// (10, 5, 'neigh_op_tnr_2')
// (10, 6, 'local_g3_2')
// (10, 6, 'lutff_1/in_0')
// (10, 6, 'neigh_op_rgt_2')
// (10, 7, 'neigh_op_bnr_2')
// (11, 5, 'local_g1_2')
// (11, 5, 'lutff_2/in_3')
// (11, 5, 'neigh_op_top_2')
// (11, 6, 'local_g3_2')
// (11, 6, 'lutff_2/out')
// (11, 6, 'lutff_5/in_2')
// (11, 7, 'neigh_op_bot_2')
// (12, 5, 'neigh_op_tnl_2')
// (12, 6, 'neigh_op_lft_2')
// (12, 7, 'neigh_op_bnl_2')

wire n1425;
// (10, 5, 'local_g3_5')
// (10, 5, 'lutff_0/in_0')
// (10, 5, 'neigh_op_tnr_5')
// (10, 6, 'neigh_op_rgt_5')
// (10, 7, 'neigh_op_bnr_5')
// (11, 0, 'span12_vert_21')
// (11, 1, 'sp12_v_b_21')
// (11, 2, 'sp12_v_b_18')
// (11, 3, 'sp12_v_b_17')
// (11, 3, 'sp4_r_v_b_46')
// (11, 4, 'sp12_v_b_14')
// (11, 4, 'sp4_r_v_b_35')
// (11, 5, 'local_g1_5')
// (11, 5, 'lutff_5/in_1')
// (11, 5, 'neigh_op_top_5')
// (11, 5, 'sp12_v_b_13')
// (11, 5, 'sp4_r_v_b_22')
// (11, 6, 'lutff_5/out')
// (11, 6, 'sp12_v_b_10')
// (11, 6, 'sp4_r_v_b_11')
// (11, 7, 'neigh_op_bot_5')
// (11, 7, 'sp12_v_b_9')
// (11, 8, 'sp12_v_b_6')
// (11, 9, 'sp12_v_b_5')
// (11, 10, 'local_g3_2')
// (11, 10, 'lutff_4/in_3')
// (11, 10, 'lutff_6/in_3')
// (11, 10, 'sp12_v_b_2')
// (11, 11, 'sp12_v_b_1')
// (12, 2, 'local_g1_3')
// (12, 2, 'lutff_3/in_1')
// (12, 2, 'sp4_h_r_11')
// (12, 2, 'sp4_v_t_46')
// (12, 3, 'sp4_v_b_46')
// (12, 4, 'sp4_v_b_35')
// (12, 5, 'neigh_op_tnl_5')
// (12, 5, 'sp4_v_b_22')
// (12, 6, 'neigh_op_lft_5')
// (12, 6, 'sp4_v_b_11')
// (12, 7, 'neigh_op_bnl_5')
// (13, 2, 'sp4_h_r_22')
// (14, 2, 'sp4_h_r_35')
// (15, 2, 'sp4_h_r_46')
// (16, 2, 'sp4_h_l_46')

wire n1426;
// (10, 5, 'neigh_op_tnr_0')
// (10, 6, 'neigh_op_rgt_0')
// (10, 7, 'neigh_op_bnr_0')
// (11, 3, 'sp4_r_v_b_36')
// (11, 3, 'sp4_r_v_b_43')
// (11, 4, 'sp4_r_v_b_25')
// (11, 4, 'sp4_r_v_b_30')
// (11, 5, 'neigh_op_top_0')
// (11, 5, 'sp4_r_v_b_12')
// (11, 5, 'sp4_r_v_b_19')
// (11, 5, 'sp4_r_v_b_44')
// (11, 6, 'local_g0_2')
// (11, 6, 'lutff_0/out')
// (11, 6, 'lutff_global/cen')
// (11, 6, 'sp4_r_v_b_1')
// (11, 6, 'sp4_r_v_b_33')
// (11, 6, 'sp4_r_v_b_6')
// (11, 7, 'neigh_op_bot_0')
// (11, 7, 'sp4_r_v_b_20')
// (11, 8, 'sp4_r_v_b_9')
// (12, 2, 'sp4_h_r_6')
// (12, 2, 'sp4_v_t_36')
// (12, 2, 'sp4_v_t_43')
// (12, 3, 'sp4_v_b_36')
// (12, 3, 'sp4_v_b_43')
// (12, 4, 'sp4_v_b_25')
// (12, 4, 'sp4_v_b_30')
// (12, 4, 'sp4_v_t_44')
// (12, 5, 'local_g1_3')
// (12, 5, 'lutff_global/cen')
// (12, 5, 'neigh_op_tnl_0')
// (12, 5, 'sp4_v_b_12')
// (12, 5, 'sp4_v_b_19')
// (12, 5, 'sp4_v_b_44')
// (12, 6, 'neigh_op_lft_0')
// (12, 6, 'sp4_v_b_1')
// (12, 6, 'sp4_v_b_33')
// (12, 6, 'sp4_v_b_6')
// (12, 7, 'neigh_op_bnl_0')
// (12, 7, 'sp4_v_b_20')
// (12, 8, 'sp4_v_b_9')
// (13, 2, 'sp4_h_r_19')
// (14, 2, 'sp4_h_r_30')
// (15, 2, 'sp4_h_r_43')
// (16, 2, 'sp4_h_l_43')

reg n1427 = 0;
// (10, 5, 'neigh_op_tnr_3')
// (10, 6, 'neigh_op_rgt_3')
// (10, 6, 'sp4_h_r_11')
// (10, 7, 'local_g1_3')
// (10, 7, 'lutff_5/in_1')
// (10, 7, 'neigh_op_bnr_3')
// (11, 5, 'neigh_op_top_3')
// (11, 6, 'lutff_3/out')
// (11, 6, 'sp4_h_r_22')
// (11, 7, 'neigh_op_bot_3')
// (12, 5, 'neigh_op_tnl_3')
// (12, 6, 'neigh_op_lft_3')
// (12, 6, 'sp4_h_r_35')
// (12, 7, 'local_g2_3')
// (12, 7, 'lutff_2/in_3')
// (12, 7, 'lutff_5/in_2')
// (12, 7, 'neigh_op_bnl_3')
// (13, 3, 'sp4_r_v_b_46')
// (13, 4, 'local_g2_3')
// (13, 4, 'lutff_5/in_2')
// (13, 4, 'sp4_r_v_b_35')
// (13, 5, 'sp4_r_v_b_22')
// (13, 6, 'sp4_h_r_46')
// (13, 6, 'sp4_r_v_b_11')
// (14, 2, 'sp4_v_t_46')
// (14, 3, 'sp4_v_b_46')
// (14, 4, 'sp4_v_b_35')
// (14, 5, 'sp4_v_b_22')
// (14, 6, 'sp4_h_l_46')
// (14, 6, 'sp4_v_b_11')

reg n1428 = 0;
// (10, 5, 'neigh_op_tnr_6')
// (10, 5, 'sp4_r_v_b_41')
// (10, 6, 'neigh_op_rgt_6')
// (10, 6, 'sp4_r_v_b_28')
// (10, 7, 'neigh_op_bnr_6')
// (10, 7, 'sp4_r_v_b_17')
// (10, 8, 'sp4_r_v_b_4')
// (11, 4, 'sp4_h_r_9')
// (11, 4, 'sp4_v_t_41')
// (11, 5, 'neigh_op_top_6')
// (11, 5, 'sp4_v_b_41')
// (11, 6, 'lutff_6/out')
// (11, 6, 'sp4_r_v_b_45')
// (11, 6, 'sp4_v_b_28')
// (11, 7, 'neigh_op_bot_6')
// (11, 7, 'sp4_r_v_b_32')
// (11, 7, 'sp4_v_b_17')
// (11, 8, 'local_g3_5')
// (11, 8, 'lutff_6/in_2')
// (11, 8, 'sp4_r_v_b_21')
// (11, 8, 'sp4_v_b_4')
// (11, 9, 'sp4_r_v_b_8')
// (12, 4, 'sp4_h_r_20')
// (12, 5, 'neigh_op_tnl_6')
// (12, 5, 'sp4_v_t_45')
// (12, 6, 'neigh_op_lft_6')
// (12, 6, 'sp4_v_b_45')
// (12, 7, 'neigh_op_bnl_6')
// (12, 7, 'sp4_v_b_32')
// (12, 8, 'local_g0_5')
// (12, 8, 'lutff_3/in_2')
// (12, 8, 'lutff_7/in_0')
// (12, 8, 'sp4_v_b_21')
// (12, 9, 'sp4_v_b_8')
// (13, 4, 'sp4_h_r_33')
// (14, 4, 'local_g3_4')
// (14, 4, 'lutff_3/in_2')
// (14, 4, 'sp4_h_r_44')
// (15, 4, 'sp4_h_l_44')

reg n1429 = 0;
// (10, 5, 'neigh_op_tnr_7')
// (10, 6, 'neigh_op_rgt_7')
// (10, 7, 'neigh_op_bnr_7')
// (11, 4, 'sp4_r_v_b_39')
// (11, 5, 'neigh_op_top_7')
// (11, 5, 'sp4_r_v_b_26')
// (11, 6, 'lutff_7/out')
// (11, 6, 'sp4_r_v_b_15')
// (11, 6, 'sp4_r_v_b_47')
// (11, 7, 'neigh_op_bot_7')
// (11, 7, 'sp4_r_v_b_2')
// (11, 7, 'sp4_r_v_b_34')
// (11, 8, 'sp4_r_v_b_23')
// (11, 9, 'local_g2_2')
// (11, 9, 'lutff_5/in_3')
// (11, 9, 'sp4_r_v_b_10')
// (12, 3, 'sp4_h_r_2')
// (12, 3, 'sp4_v_t_39')
// (12, 4, 'sp4_v_b_39')
// (12, 5, 'neigh_op_tnl_7')
// (12, 5, 'sp4_v_b_26')
// (12, 5, 'sp4_v_t_47')
// (12, 6, 'neigh_op_lft_7')
// (12, 6, 'sp4_v_b_15')
// (12, 6, 'sp4_v_b_47')
// (12, 7, 'local_g0_2')
// (12, 7, 'lutff_1/in_1')
// (12, 7, 'neigh_op_bnl_7')
// (12, 7, 'sp4_v_b_2')
// (12, 7, 'sp4_v_b_34')
// (12, 8, 'sp4_v_b_23')
// (12, 9, 'local_g1_2')
// (12, 9, 'lutff_5/in_0')
// (12, 9, 'sp4_v_b_10')
// (13, 3, 'local_g0_7')
// (13, 3, 'lutff_3/in_0')
// (13, 3, 'sp4_h_r_15')
// (14, 3, 'sp4_h_r_26')
// (15, 3, 'sp4_h_r_39')
// (16, 3, 'sp4_h_l_39')

wire n1430;
// (10, 5, 'sp4_r_v_b_42')
// (10, 6, 'neigh_op_tnr_1')
// (10, 6, 'sp4_r_v_b_31')
// (10, 7, 'neigh_op_rgt_1')
// (10, 7, 'sp4_r_v_b_18')
// (10, 8, 'neigh_op_bnr_1')
// (10, 8, 'sp4_r_v_b_7')
// (11, 4, 'sp4_r_v_b_38')
// (11, 4, 'sp4_v_t_42')
// (11, 5, 'sp4_r_v_b_27')
// (11, 5, 'sp4_v_b_42')
// (11, 6, 'neigh_op_top_1')
// (11, 6, 'sp4_r_v_b_14')
// (11, 6, 'sp4_v_b_31')
// (11, 7, 'lutff_1/out')
// (11, 7, 'sp4_r_v_b_3')
// (11, 7, 'sp4_v_b_18')
// (11, 8, 'neigh_op_bot_1')
// (11, 8, 'sp4_h_r_7')
// (11, 8, 'sp4_r_v_b_43')
// (11, 8, 'sp4_v_b_7')
// (11, 9, 'sp4_r_v_b_30')
// (11, 10, 'sp4_r_v_b_19')
// (11, 11, 'sp4_r_v_b_6')
// (12, 3, 'sp4_v_t_38')
// (12, 4, 'sp4_v_b_38')
// (12, 5, 'sp4_v_b_27')
// (12, 6, 'neigh_op_tnl_1')
// (12, 6, 'sp4_v_b_14')
// (12, 7, 'neigh_op_lft_1')
// (12, 7, 'sp4_v_b_3')
// (12, 7, 'sp4_v_t_43')
// (12, 8, 'local_g0_2')
// (12, 8, 'lutff_global/cen')
// (12, 8, 'neigh_op_bnl_1')
// (12, 8, 'sp4_h_r_18')
// (12, 8, 'sp4_v_b_43')
// (12, 9, 'sp4_v_b_30')
// (12, 10, 'local_g1_3')
// (12, 10, 'lutff_global/cen')
// (12, 10, 'sp4_v_b_19')
// (12, 11, 'sp4_v_b_6')
// (13, 8, 'sp4_h_r_31')
// (14, 8, 'sp4_h_r_42')
// (15, 8, 'sp4_h_l_42')

wire n1431;
// (10, 6, 'neigh_op_tnr_4')
// (10, 7, 'local_g2_4')
// (10, 7, 'lutff_7/in_3')
// (10, 7, 'neigh_op_rgt_4')
// (10, 8, 'neigh_op_bnr_4')
// (11, 6, 'neigh_op_top_4')
// (11, 7, 'lutff_4/out')
// (11, 8, 'neigh_op_bot_4')
// (12, 6, 'neigh_op_tnl_4')
// (12, 7, 'neigh_op_lft_4')
// (12, 8, 'neigh_op_bnl_4')

wire n1432;
// (10, 6, 'neigh_op_tnr_5')
// (10, 7, 'neigh_op_rgt_5')
// (10, 8, 'neigh_op_bnr_5')
// (11, 6, 'neigh_op_top_5')
// (11, 7, 'local_g1_5')
// (11, 7, 'lutff_1/in_3')
// (11, 7, 'lutff_5/out')
// (11, 8, 'neigh_op_bot_5')
// (12, 6, 'neigh_op_tnl_5')
// (12, 7, 'neigh_op_lft_5')
// (12, 8, 'neigh_op_bnl_5')

wire n1433;
// (10, 6, 'sp4_h_r_7')
// (11, 6, 'sp4_h_r_18')
// (12, 6, 'sp4_h_r_31')
// (13, 3, 'neigh_op_tnr_5')
// (13, 3, 'sp4_r_v_b_39')
// (13, 3, 'sp4_r_v_b_42')
// (13, 4, 'local_g0_2')
// (13, 4, 'lutff_global/cen')
// (13, 4, 'neigh_op_rgt_5')
// (13, 4, 'sp4_r_v_b_26')
// (13, 4, 'sp4_r_v_b_31')
// (13, 5, 'neigh_op_bnr_5')
// (13, 5, 'sp4_r_v_b_15')
// (13, 5, 'sp4_r_v_b_18')
// (13, 6, 'local_g2_2')
// (13, 6, 'lutff_global/cen')
// (13, 6, 'sp4_h_r_42')
// (13, 6, 'sp4_r_v_b_2')
// (13, 6, 'sp4_r_v_b_7')
// (14, 2, 'sp4_h_r_7')
// (14, 2, 'sp4_v_t_39')
// (14, 2, 'sp4_v_t_42')
// (14, 3, 'neigh_op_top_5')
// (14, 3, 'sp4_v_b_39')
// (14, 3, 'sp4_v_b_42')
// (14, 4, 'lutff_5/out')
// (14, 4, 'sp4_v_b_26')
// (14, 4, 'sp4_v_b_31')
// (14, 5, 'local_g0_2')
// (14, 5, 'lutff_global/cen')
// (14, 5, 'neigh_op_bot_5')
// (14, 5, 'sp4_v_b_15')
// (14, 5, 'sp4_v_b_18')
// (14, 6, 'sp4_h_l_42')
// (14, 6, 'sp4_h_r_10')
// (14, 6, 'sp4_v_b_2')
// (14, 6, 'sp4_v_b_7')
// (15, 2, 'sp4_h_r_18')
// (15, 3, 'neigh_op_tnl_5')
// (15, 4, 'neigh_op_lft_5')
// (15, 5, 'neigh_op_bnl_5')
// (15, 6, 'sp4_h_r_23')
// (16, 2, 'sp4_h_r_31')
// (16, 6, 'local_g2_2')
// (16, 6, 'lutff_global/cen')
// (16, 6, 'sp4_h_r_34')
// (17, 2, 'sp4_h_r_42')
// (17, 6, 'sp4_h_r_47')
// (18, 2, 'sp4_h_l_42')
// (18, 6, 'sp4_h_l_47')

reg n1434 = 0;
// (10, 6, 'sp4_h_r_9')
// (11, 6, 'sp4_h_r_20')
// (12, 6, 'local_g2_1')
// (12, 6, 'lutff_6/in_1')
// (12, 6, 'sp4_h_r_33')
// (12, 9, 'neigh_op_tnr_4')
// (12, 10, 'neigh_op_rgt_4')
// (12, 11, 'local_g0_4')
// (12, 11, 'lutff_6/in_2')
// (12, 11, 'neigh_op_bnr_4')
// (13, 6, 'sp4_h_r_44')
// (13, 7, 'sp4_r_v_b_44')
// (13, 8, 'sp4_r_v_b_33')
// (13, 9, 'neigh_op_top_4')
// (13, 9, 'sp4_r_v_b_20')
// (13, 10, 'lutff_4/out')
// (13, 10, 'sp4_r_v_b_9')
// (13, 11, 'neigh_op_bot_4')
// (13, 11, 'sp4_r_v_b_40')
// (13, 12, 'sp4_r_v_b_29')
// (13, 13, 'sp4_r_v_b_16')
// (13, 14, 'sp4_r_v_b_5')
// (14, 6, 'local_g0_1')
// (14, 6, 'lutff_0/in_1')
// (14, 6, 'sp4_h_l_44')
// (14, 6, 'sp4_h_r_9')
// (14, 6, 'sp4_v_t_44')
// (14, 7, 'sp4_v_b_44')
// (14, 8, 'sp4_v_b_33')
// (14, 9, 'neigh_op_tnl_4')
// (14, 9, 'sp4_v_b_20')
// (14, 10, 'neigh_op_lft_4')
// (14, 10, 'sp4_v_b_9')
// (14, 10, 'sp4_v_t_40')
// (14, 11, 'neigh_op_bnl_4')
// (14, 11, 'sp4_v_b_40')
// (14, 12, 'sp4_v_b_29')
// (14, 13, 'local_g0_0')
// (14, 13, 'lutff_4/in_0')
// (14, 13, 'sp4_v_b_16')
// (14, 14, 'sp4_v_b_5')
// (15, 6, 'sp4_h_r_20')
// (16, 6, 'sp4_h_r_33')
// (17, 6, 'sp4_h_r_44')
// (18, 6, 'sp4_h_l_44')

reg n1435 = 0;
// (10, 6, 'sp4_r_v_b_40')
// (10, 7, 'sp4_r_v_b_29')
// (10, 8, 'sp4_r_v_b_16')
// (10, 9, 'local_g1_5')
// (10, 9, 'lutff_0/in_0')
// (10, 9, 'sp4_r_v_b_5')
// (11, 4, 'neigh_op_tnr_0')
// (11, 5, 'neigh_op_rgt_0')
// (11, 5, 'sp4_h_r_5')
// (11, 5, 'sp4_v_t_40')
// (11, 6, 'neigh_op_bnr_0')
// (11, 6, 'sp4_r_v_b_43')
// (11, 6, 'sp4_v_b_40')
// (11, 7, 'sp4_r_v_b_30')
// (11, 7, 'sp4_v_b_29')
// (11, 8, 'sp4_r_v_b_19')
// (11, 8, 'sp4_v_b_16')
// (11, 9, 'sp4_r_v_b_6')
// (11, 9, 'sp4_v_b_5')
// (12, 4, 'neigh_op_top_0')
// (12, 5, 'lutff_0/out')
// (12, 5, 'sp4_h_r_0')
// (12, 5, 'sp4_h_r_16')
// (12, 5, 'sp4_v_t_43')
// (12, 6, 'local_g1_0')
// (12, 6, 'lutff_2/in_3')
// (12, 6, 'neigh_op_bot_0')
// (12, 6, 'sp4_v_b_43')
// (12, 7, 'sp4_v_b_30')
// (12, 8, 'sp4_v_b_19')
// (12, 9, 'local_g0_6')
// (12, 9, 'lutff_3/in_3')
// (12, 9, 'sp4_v_b_6')
// (13, 4, 'local_g2_0')
// (13, 4, 'lutff_6/in_0')
// (13, 4, 'neigh_op_tnl_0')
// (13, 5, 'neigh_op_lft_0')
// (13, 5, 'sp4_h_r_13')
// (13, 5, 'sp4_h_r_29')
// (13, 6, 'neigh_op_bnl_0')
// (14, 5, 'sp4_h_r_24')
// (14, 5, 'sp4_h_r_40')
// (15, 5, 'sp4_h_l_40')
// (15, 5, 'sp4_h_r_37')
// (16, 5, 'sp4_h_l_37')

reg n1436 = 0;
// (10, 7, 'neigh_op_tnr_0')
// (10, 8, 'local_g2_0')
// (10, 8, 'lutff_5/in_1')
// (10, 8, 'neigh_op_rgt_0')
// (10, 9, 'neigh_op_bnr_0')
// (11, 4, 'sp12_v_t_23')
// (11, 5, 'sp12_v_b_23')
// (11, 6, 'sp12_v_b_20')
// (11, 7, 'neigh_op_top_0')
// (11, 7, 'sp12_v_b_19')
// (11, 8, 'lutff_0/out')
// (11, 8, 'sp12_v_b_16')
// (11, 9, 'neigh_op_bot_0')
// (11, 9, 'sp12_v_b_15')
// (11, 10, 'sp12_v_b_12')
// (11, 11, 'sp12_v_b_11')
// (11, 12, 'sp12_v_b_8')
// (11, 13, 'sp12_v_b_7')
// (11, 14, 'local_g2_4')
// (11, 14, 'lutff_6/in_2')
// (11, 14, 'sp12_v_b_4')
// (11, 15, 'local_g3_3')
// (11, 15, 'lutff_5/in_1')
// (11, 15, 'lutff_7/in_1')
// (11, 15, 'sp12_v_b_3')
// (11, 16, 'sp12_v_b_0')
// (12, 7, 'neigh_op_tnl_0')
// (12, 8, 'neigh_op_lft_0')
// (12, 9, 'neigh_op_bnl_0')

reg n1437 = 0;
// (10, 7, 'neigh_op_tnr_2')
// (10, 8, 'neigh_op_rgt_2')
// (10, 9, 'neigh_op_bnr_2')
// (11, 7, 'neigh_op_top_2')
// (11, 8, 'lutff_2/out')
// (11, 9, 'local_g1_2')
// (11, 9, 'lutff_3/in_0')
// (11, 9, 'neigh_op_bot_2')
// (12, 7, 'neigh_op_tnl_2')
// (12, 8, 'neigh_op_lft_2')
// (12, 9, 'neigh_op_bnl_2')

reg n1438 = 0;
// (10, 7, 'neigh_op_tnr_3')
// (10, 8, 'neigh_op_rgt_3')
// (10, 9, 'neigh_op_bnr_3')
// (11, 7, 'neigh_op_top_3')
// (11, 8, 'lutff_3/out')
// (11, 9, 'local_g0_3')
// (11, 9, 'lutff_3/in_2')
// (11, 9, 'neigh_op_bot_3')
// (12, 7, 'neigh_op_tnl_3')
// (12, 8, 'neigh_op_lft_3')
// (12, 9, 'neigh_op_bnl_3')

reg n1439 = 0;
// (10, 7, 'neigh_op_tnr_4')
// (10, 8, 'local_g2_4')
// (10, 8, 'lutff_7/in_3')
// (10, 8, 'neigh_op_rgt_4')
// (10, 9, 'neigh_op_bnr_4')
// (11, 7, 'neigh_op_top_4')
// (11, 8, 'lutff_4/out')
// (11, 9, 'neigh_op_bot_4')
// (12, 7, 'neigh_op_tnl_4')
// (12, 8, 'neigh_op_lft_4')
// (12, 9, 'neigh_op_bnl_4')

reg n1440 = 0;
// (10, 7, 'neigh_op_tnr_5')
// (10, 8, 'local_g2_5')
// (10, 8, 'lutff_1/in_0')
// (10, 8, 'neigh_op_rgt_5')
// (10, 9, 'neigh_op_bnr_5')
// (11, 7, 'neigh_op_top_5')
// (11, 8, 'lutff_5/out')
// (11, 9, 'neigh_op_bot_5')
// (12, 7, 'neigh_op_tnl_5')
// (12, 8, 'neigh_op_lft_5')
// (12, 9, 'neigh_op_bnl_5')

reg n1441 = 0;
// (10, 7, 'neigh_op_tnr_6')
// (10, 8, 'local_g3_6')
// (10, 8, 'lutff_7/in_0')
// (10, 8, 'neigh_op_rgt_6')
// (10, 9, 'neigh_op_bnr_6')
// (11, 7, 'neigh_op_top_6')
// (11, 8, 'lutff_6/out')
// (11, 9, 'neigh_op_bot_6')
// (12, 7, 'neigh_op_tnl_6')
// (12, 8, 'neigh_op_lft_6')
// (12, 9, 'neigh_op_bnl_6')

reg n1442 = 0;
// (10, 7, 'neigh_op_tnr_7')
// (10, 8, 'local_g2_7')
// (10, 8, 'lutff_1/in_2')
// (10, 8, 'neigh_op_rgt_7')
// (10, 9, 'neigh_op_bnr_7')
// (11, 7, 'neigh_op_top_7')
// (11, 8, 'lutff_7/out')
// (11, 9, 'neigh_op_bot_7')
// (12, 7, 'neigh_op_tnl_7')
// (12, 8, 'neigh_op_lft_7')
// (12, 9, 'neigh_op_bnl_7')

wire n1443;
// (10, 7, 'sp4_h_r_5')
// (11, 7, 'local_g1_0')
// (11, 7, 'lutff_3/in_0')
// (11, 7, 'sp4_h_r_16')
// (12, 7, 'sp4_h_r_29')
// (13, 4, 'neigh_op_tnr_4')
// (13, 4, 'sp4_r_v_b_37')
// (13, 5, 'neigh_op_rgt_4')
// (13, 5, 'sp4_r_v_b_24')
// (13, 6, 'neigh_op_bnr_4')
// (13, 6, 'sp4_r_v_b_13')
// (13, 7, 'sp4_h_r_40')
// (13, 7, 'sp4_r_v_b_0')
// (14, 3, 'sp4_v_t_37')
// (14, 4, 'neigh_op_top_4')
// (14, 4, 'sp4_v_b_37')
// (14, 5, 'lutff_4/out')
// (14, 5, 'sp4_v_b_24')
// (14, 6, 'neigh_op_bot_4')
// (14, 6, 'sp4_v_b_13')
// (14, 7, 'sp4_h_l_40')
// (14, 7, 'sp4_v_b_0')
// (15, 4, 'neigh_op_tnl_4')
// (15, 5, 'neigh_op_lft_4')
// (15, 6, 'neigh_op_bnl_4')

wire n1444;
// (10, 7, 'sp4_h_r_6')
// (11, 6, 'neigh_op_tnr_7')
// (11, 7, 'local_g0_3')
// (11, 7, 'lutff_3/in_2')
// (11, 7, 'neigh_op_rgt_7')
// (11, 7, 'sp4_h_r_19')
// (11, 8, 'neigh_op_bnr_7')
// (12, 6, 'neigh_op_top_7')
// (12, 7, 'lutff_7/out')
// (12, 7, 'sp4_h_r_30')
// (12, 8, 'neigh_op_bot_7')
// (13, 6, 'neigh_op_tnl_7')
// (13, 7, 'neigh_op_lft_7')
// (13, 7, 'sp4_h_r_43')
// (13, 8, 'neigh_op_bnl_7')
// (14, 7, 'sp4_h_l_43')

wire n1445;
// (10, 7, 'sp4_r_v_b_46')
// (10, 8, 'neigh_op_tnr_3')
// (10, 8, 'sp4_r_v_b_35')
// (10, 9, 'neigh_op_rgt_3')
// (10, 9, 'sp4_r_v_b_22')
// (10, 10, 'neigh_op_bnr_3')
// (10, 10, 'sp4_r_v_b_11')
// (10, 11, 'sp4_r_v_b_39')
// (10, 12, 'sp4_r_v_b_26')
// (10, 13, 'sp4_r_v_b_15')
// (10, 14, 'sp4_r_v_b_2')
// (11, 6, 'sp4_v_t_46')
// (11, 7, 'sp4_v_b_46')
// (11, 8, 'neigh_op_top_3')
// (11, 8, 'sp4_v_b_35')
// (11, 9, 'lutff_3/out')
// (11, 9, 'sp4_v_b_22')
// (11, 10, 'neigh_op_bot_3')
// (11, 10, 'sp4_v_b_11')
// (11, 10, 'sp4_v_t_39')
// (11, 11, 'sp4_v_b_39')
// (11, 12, 'sp4_v_b_26')
// (11, 13, 'sp4_v_b_15')
// (11, 14, 'local_g0_2')
// (11, 14, 'lutff_3/in_1')
// (11, 14, 'sp4_v_b_2')
// (12, 8, 'neigh_op_tnl_3')
// (12, 9, 'neigh_op_lft_3')
// (12, 10, 'neigh_op_bnl_3')

reg n1446 = 0;
// (10, 8, 'neigh_op_tnr_0')
// (10, 9, 'local_g2_0')
// (10, 9, 'lutff_3/in_3')
// (10, 9, 'neigh_op_rgt_0')
// (10, 10, 'neigh_op_bnr_0')
// (11, 8, 'neigh_op_top_0')
// (11, 9, 'local_g1_0')
// (11, 9, 'lutff_0/out')
// (11, 9, 'lutff_2/in_3')
// (11, 9, 'lutff_7/in_2')
// (11, 10, 'neigh_op_bot_0')
// (12, 8, 'neigh_op_tnl_0')
// (12, 9, 'neigh_op_lft_0')
// (12, 10, 'neigh_op_bnl_0')

reg n1447 = 0;
// (10, 8, 'neigh_op_tnr_1')
// (10, 9, 'local_g2_1')
// (10, 9, 'lutff_3/in_0')
// (10, 9, 'neigh_op_rgt_1')
// (10, 10, 'neigh_op_bnr_1')
// (11, 8, 'neigh_op_top_1')
// (11, 9, 'lutff_1/out')
// (11, 10, 'neigh_op_bot_1')
// (12, 8, 'neigh_op_tnl_1')
// (12, 9, 'neigh_op_lft_1')
// (12, 10, 'neigh_op_bnl_1')

wire n1448;
// (10, 8, 'neigh_op_tnr_2')
// (10, 9, 'neigh_op_rgt_2')
// (10, 10, 'neigh_op_bnr_2')
// (11, 8, 'neigh_op_top_2')
// (11, 9, 'lutff_2/out')
// (11, 10, 'local_g1_2')
// (11, 10, 'lutff_5/in_0')
// (11, 10, 'neigh_op_bot_2')
// (12, 8, 'neigh_op_tnl_2')
// (12, 9, 'neigh_op_lft_2')
// (12, 10, 'neigh_op_bnl_2')

reg n1449 = 0;
// (10, 8, 'neigh_op_tnr_4')
// (10, 9, 'neigh_op_rgt_4')
// (10, 10, 'neigh_op_bnr_4')
// (11, 8, 'neigh_op_top_4')
// (11, 9, 'local_g3_4')
// (11, 9, 'lutff_4/out')
// (11, 9, 'lutff_7/in_0')
// (11, 10, 'neigh_op_bot_4')
// (12, 8, 'neigh_op_tnl_4')
// (12, 9, 'neigh_op_lft_4')
// (12, 10, 'neigh_op_bnl_4')

reg n1450 = 0;
// (10, 8, 'neigh_op_tnr_5')
// (10, 9, 'local_g2_5')
// (10, 9, 'lutff_2/in_3')
// (10, 9, 'neigh_op_rgt_5')
// (10, 10, 'neigh_op_bnr_5')
// (11, 8, 'neigh_op_top_5')
// (11, 9, 'lutff_5/out')
// (11, 10, 'neigh_op_bot_5')
// (12, 8, 'neigh_op_tnl_5')
// (12, 9, 'neigh_op_lft_5')
// (12, 10, 'neigh_op_bnl_5')

wire n1451;
// (10, 8, 'neigh_op_tnr_7')
// (10, 9, 'neigh_op_rgt_7')
// (10, 10, 'neigh_op_bnr_7')
// (11, 8, 'neigh_op_top_7')
// (11, 9, 'lutff_7/out')
// (11, 10, 'local_g0_7')
// (11, 10, 'lutff_1/in_0')
// (11, 10, 'neigh_op_bot_7')
// (12, 8, 'neigh_op_tnl_7')
// (12, 9, 'neigh_op_lft_7')
// (12, 10, 'neigh_op_bnl_7')

reg n1452 = 0;
// (10, 8, 'sp4_h_r_11')
// (11, 8, 'sp4_h_r_22')
// (12, 8, 'local_g2_3')
// (12, 8, 'lutff_1/in_0')
// (12, 8, 'sp4_h_r_35')
// (12, 11, 'sp4_h_r_8')
// (13, 5, 'sp4_r_v_b_45')
// (13, 6, 'sp4_r_v_b_32')
// (13, 7, 'sp4_r_v_b_21')
// (13, 8, 'sp4_h_r_46')
// (13, 8, 'sp4_r_v_b_8')
// (13, 9, 'sp4_r_v_b_40')
// (13, 10, 'neigh_op_tnr_0')
// (13, 10, 'sp4_r_v_b_29')
// (13, 11, 'local_g2_0')
// (13, 11, 'lutff_6/in_0')
// (13, 11, 'neigh_op_rgt_0')
// (13, 11, 'sp4_h_r_21')
// (13, 11, 'sp4_r_v_b_16')
// (13, 12, 'neigh_op_bnr_0')
// (13, 12, 'sp4_r_v_b_5')
// (14, 4, 'sp4_v_t_45')
// (14, 5, 'sp4_v_b_45')
// (14, 6, 'sp4_v_b_32')
// (14, 7, 'local_g0_5')
// (14, 7, 'lutff_2/in_1')
// (14, 7, 'sp4_v_b_21')
// (14, 8, 'sp4_h_l_46')
// (14, 8, 'sp4_v_b_8')
// (14, 8, 'sp4_v_t_40')
// (14, 9, 'sp4_v_b_40')
// (14, 10, 'neigh_op_top_0')
// (14, 10, 'sp4_v_b_29')
// (14, 11, 'lutff_0/out')
// (14, 11, 'sp4_h_r_32')
// (14, 11, 'sp4_v_b_16')
// (14, 12, 'local_g1_0')
// (14, 12, 'lutff_2/in_1')
// (14, 12, 'neigh_op_bot_0')
// (14, 12, 'sp4_v_b_5')
// (15, 4, 'sp4_r_v_b_47')
// (15, 5, 'sp4_r_v_b_34')
// (15, 6, 'sp4_r_v_b_23')
// (15, 7, 'sp4_r_v_b_10')
// (15, 8, 'sp4_r_v_b_39')
// (15, 9, 'sp4_r_v_b_26')
// (15, 10, 'neigh_op_tnl_0')
// (15, 10, 'sp4_r_v_b_15')
// (15, 11, 'neigh_op_lft_0')
// (15, 11, 'sp4_h_r_45')
// (15, 11, 'sp4_r_v_b_2')
// (15, 12, 'local_g3_0')
// (15, 12, 'lutff_5/in_0')
// (15, 12, 'neigh_op_bnl_0')
// (16, 3, 'sp4_v_t_47')
// (16, 4, 'sp4_v_b_47')
// (16, 5, 'sp4_v_b_34')
// (16, 6, 'local_g1_7')
// (16, 6, 'lutff_4/in_2')
// (16, 6, 'sp4_v_b_23')
// (16, 7, 'sp4_v_b_10')
// (16, 7, 'sp4_v_t_39')
// (16, 8, 'sp4_v_b_39')
// (16, 9, 'sp4_v_b_26')
// (16, 10, 'sp4_v_b_15')
// (16, 11, 'sp4_h_l_45')
// (16, 11, 'sp4_v_b_2')

reg n1453 = 0;
// (10, 8, 'sp4_h_r_9')
// (11, 8, 'sp4_h_r_20')
// (12, 8, 'local_g3_1')
// (12, 8, 'lutff_3/in_3')
// (12, 8, 'sp4_h_r_33')
// (13, 8, 'sp4_h_r_44')
// (13, 9, 'sp4_r_v_b_38')
// (13, 10, 'neigh_op_tnr_7')
// (13, 10, 'sp4_r_v_b_27')
// (13, 11, 'local_g2_7')
// (13, 11, 'lutff_2/in_1')
// (13, 11, 'neigh_op_rgt_7')
// (13, 11, 'sp4_h_r_3')
// (13, 11, 'sp4_r_v_b_14')
// (13, 12, 'neigh_op_bnr_7')
// (13, 12, 'sp4_r_v_b_3')
// (14, 8, 'sp4_h_l_44')
// (14, 8, 'sp4_v_t_38')
// (14, 9, 'sp4_v_b_38')
// (14, 10, 'neigh_op_top_7')
// (14, 10, 'sp4_v_b_27')
// (14, 11, 'lutff_7/out')
// (14, 11, 'sp4_h_r_14')
// (14, 11, 'sp4_v_b_14')
// (14, 12, 'local_g1_7')
// (14, 12, 'lutff_1/in_3')
// (14, 12, 'neigh_op_bot_7')
// (14, 12, 'sp4_h_r_9')
// (14, 12, 'sp4_v_b_3')
// (15, 10, 'neigh_op_tnl_7')
// (15, 11, 'neigh_op_lft_7')
// (15, 11, 'sp4_h_r_27')
// (15, 12, 'neigh_op_bnl_7')
// (15, 12, 'sp4_h_r_20')
// (16, 4, 'sp4_r_v_b_37')
// (16, 4, 'sp4_r_v_b_40')
// (16, 5, 'local_g0_5')
// (16, 5, 'lutff_6/in_3')
// (16, 5, 'sp4_r_v_b_24')
// (16, 5, 'sp4_r_v_b_29')
// (16, 6, 'local_g2_5')
// (16, 6, 'lutff_2/in_3')
// (16, 6, 'sp4_r_v_b_13')
// (16, 6, 'sp4_r_v_b_16')
// (16, 7, 'sp4_r_v_b_0')
// (16, 7, 'sp4_r_v_b_5')
// (16, 8, 'sp4_r_v_b_44')
// (16, 9, 'sp4_r_v_b_33')
// (16, 10, 'sp4_r_v_b_20')
// (16, 11, 'sp4_h_r_38')
// (16, 11, 'sp4_r_v_b_9')
// (16, 12, 'local_g3_1')
// (16, 12, 'lutff_4/in_2')
// (16, 12, 'sp4_h_r_33')
// (17, 3, 'sp4_v_t_37')
// (17, 3, 'sp4_v_t_40')
// (17, 4, 'sp4_v_b_37')
// (17, 4, 'sp4_v_b_40')
// (17, 5, 'sp4_v_b_24')
// (17, 5, 'sp4_v_b_29')
// (17, 6, 'sp4_v_b_13')
// (17, 6, 'sp4_v_b_16')
// (17, 7, 'sp4_v_b_0')
// (17, 7, 'sp4_v_b_5')
// (17, 7, 'sp4_v_t_44')
// (17, 8, 'sp4_v_b_44')
// (17, 9, 'sp4_v_b_33')
// (17, 10, 'sp4_v_b_20')
// (17, 11, 'sp4_h_l_38')
// (17, 11, 'sp4_v_b_9')
// (17, 12, 'sp4_h_r_44')
// (18, 12, 'sp4_h_l_44')

reg n1454 = 0;
// (10, 8, 'sp4_r_v_b_41')
// (10, 9, 'sp4_r_v_b_28')
// (10, 10, 'sp4_r_v_b_17')
// (10, 11, 'sp4_r_v_b_4')
// (11, 7, 'sp4_h_r_4')
// (11, 7, 'sp4_v_t_41')
// (11, 8, 'sp4_v_b_41')
// (11, 9, 'sp4_v_b_28')
// (11, 10, 'sp4_v_b_17')
// (11, 11, 'sp4_h_r_4')
// (11, 11, 'sp4_v_b_4')
// (12, 7, 'local_g1_1')
// (12, 7, 'lutff_2/in_0')
// (12, 7, 'sp4_h_r_17')
// (12, 10, 'neigh_op_tnr_6')
// (12, 11, 'neigh_op_rgt_6')
// (12, 11, 'sp4_h_r_17')
// (12, 12, 'neigh_op_bnr_6')
// (13, 7, 'sp4_h_r_28')
// (13, 9, 'sp4_r_v_b_37')
// (13, 10, 'local_g0_6')
// (13, 10, 'lutff_7/in_1')
// (13, 10, 'neigh_op_top_6')
// (13, 10, 'sp4_r_v_b_24')
// (13, 11, 'lutff_6/out')
// (13, 11, 'sp4_h_r_28')
// (13, 11, 'sp4_r_v_b_13')
// (13, 12, 'neigh_op_bot_6')
// (13, 12, 'sp4_r_v_b_0')
// (14, 7, 'sp4_h_r_41')
// (14, 8, 'sp4_r_v_b_47')
// (14, 8, 'sp4_v_t_37')
// (14, 9, 'sp4_r_v_b_34')
// (14, 9, 'sp4_v_b_37')
// (14, 10, 'local_g2_6')
// (14, 10, 'lutff_5/in_3')
// (14, 10, 'neigh_op_tnl_6')
// (14, 10, 'sp4_r_v_b_23')
// (14, 10, 'sp4_v_b_24')
// (14, 11, 'neigh_op_lft_6')
// (14, 11, 'sp4_h_r_41')
// (14, 11, 'sp4_r_v_b_10')
// (14, 11, 'sp4_v_b_13')
// (14, 12, 'neigh_op_bnl_6')
// (14, 12, 'sp4_h_r_0')
// (14, 12, 'sp4_r_v_b_41')
// (14, 12, 'sp4_v_b_0')
// (14, 13, 'sp4_r_v_b_28')
// (14, 14, 'local_g3_1')
// (14, 14, 'lutff_5/in_3')
// (14, 14, 'sp4_r_v_b_17')
// (14, 15, 'sp4_r_v_b_4')
// (15, 7, 'local_g1_2')
// (15, 7, 'lutff_3/in_2')
// (15, 7, 'sp4_h_l_41')
// (15, 7, 'sp4_h_r_10')
// (15, 7, 'sp4_v_t_47')
// (15, 8, 'sp4_v_b_47')
// (15, 9, 'sp4_v_b_34')
// (15, 10, 'sp4_v_b_23')
// (15, 11, 'sp4_h_l_41')
// (15, 11, 'sp4_v_b_10')
// (15, 11, 'sp4_v_t_41')
// (15, 12, 'sp4_h_r_13')
// (15, 12, 'sp4_v_b_41')
// (15, 13, 'sp4_v_b_28')
// (15, 14, 'sp4_v_b_17')
// (15, 15, 'sp4_v_b_4')
// (16, 7, 'sp4_h_r_23')
// (16, 12, 'local_g3_0')
// (16, 12, 'lutff_5/in_2')
// (16, 12, 'sp4_h_r_24')
// (17, 7, 'sp4_h_r_34')
// (17, 12, 'sp4_h_r_37')
// (18, 7, 'sp4_h_r_47')
// (18, 12, 'sp4_h_l_37')
// (19, 7, 'sp4_h_l_47')

reg n1455 = 0;
// (10, 9, 'neigh_op_tnr_0')
// (10, 10, 'local_g3_0')
// (10, 10, 'lutff_3/in_0')
// (10, 10, 'neigh_op_rgt_0')
// (10, 11, 'neigh_op_bnr_0')
// (11, 9, 'neigh_op_top_0')
// (11, 10, 'lutff_0/out')
// (11, 11, 'neigh_op_bot_0')
// (12, 9, 'neigh_op_tnl_0')
// (12, 10, 'neigh_op_lft_0')
// (12, 11, 'neigh_op_bnl_0')

wire n1456;
// (10, 9, 'neigh_op_tnr_1')
// (10, 10, 'neigh_op_rgt_1')
// (10, 11, 'local_g0_1')
// (10, 11, 'lutff_3/in_0')
// (10, 11, 'neigh_op_bnr_1')
// (11, 9, 'neigh_op_top_1')
// (11, 10, 'lutff_1/out')
// (11, 11, 'neigh_op_bot_1')
// (12, 9, 'neigh_op_tnl_1')
// (12, 10, 'neigh_op_lft_1')
// (12, 11, 'neigh_op_bnl_1')

wire n1457;
// (10, 9, 'neigh_op_tnr_2')
// (10, 10, 'neigh_op_rgt_2')
// (10, 10, 'sp4_r_v_b_36')
// (10, 11, 'neigh_op_bnr_2')
// (10, 11, 'sp4_r_v_b_25')
// (10, 11, 'sp4_r_v_b_47')
// (10, 12, 'sp4_r_v_b_12')
// (10, 12, 'sp4_r_v_b_34')
// (10, 13, 'sp4_r_v_b_1')
// (10, 13, 'sp4_r_v_b_23')
// (10, 14, 'local_g2_2')
// (10, 14, 'lutff_4/in_0')
// (10, 14, 'sp4_r_v_b_10')
// (10, 14, 'sp4_r_v_b_36')
// (10, 15, 'sp4_r_v_b_25')
// (10, 16, 'local_g2_4')
// (10, 16, 'lutff_7/in_3')
// (10, 16, 'sp4_r_v_b_12')
// (10, 17, 'sp4_r_v_b_1')
// (11, 9, 'neigh_op_top_2')
// (11, 9, 'sp4_v_t_36')
// (11, 10, 'local_g2_2')
// (11, 10, 'lutff_2/out')
// (11, 10, 'lutff_3/in_3')
// (11, 10, 'sp4_h_r_4')
// (11, 10, 'sp4_r_v_b_37')
// (11, 10, 'sp4_v_b_36')
// (11, 10, 'sp4_v_t_47')
// (11, 11, 'neigh_op_bot_2')
// (11, 11, 'sp4_r_v_b_24')
// (11, 11, 'sp4_v_b_25')
// (11, 11, 'sp4_v_b_47')
// (11, 12, 'local_g0_4')
// (11, 12, 'lutff_4/in_0')
// (11, 12, 'sp4_r_v_b_13')
// (11, 12, 'sp4_v_b_12')
// (11, 12, 'sp4_v_b_34')
// (11, 13, 'sp4_r_v_b_0')
// (11, 13, 'sp4_v_b_1')
// (11, 13, 'sp4_v_b_23')
// (11, 13, 'sp4_v_t_36')
// (11, 14, 'sp4_r_v_b_38')
// (11, 14, 'sp4_v_b_10')
// (11, 14, 'sp4_v_b_36')
// (11, 15, 'sp4_r_v_b_27')
// (11, 15, 'sp4_v_b_25')
// (11, 16, 'local_g0_4')
// (11, 16, 'local_g2_6')
// (11, 16, 'lutff_3/in_3')
// (11, 16, 'lutff_6/in_2')
// (11, 16, 'sp4_r_v_b_14')
// (11, 16, 'sp4_v_b_12')
// (11, 17, 'sp4_r_v_b_3')
// (11, 17, 'sp4_v_b_1')
// (12, 9, 'neigh_op_tnl_2')
// (12, 9, 'sp4_v_t_37')
// (12, 10, 'neigh_op_lft_2')
// (12, 10, 'sp4_h_r_17')
// (12, 10, 'sp4_v_b_37')
// (12, 11, 'neigh_op_bnl_2')
// (12, 11, 'sp4_v_b_24')
// (12, 12, 'sp4_v_b_13')
// (12, 13, 'sp4_v_b_0')
// (12, 13, 'sp4_v_t_38')
// (12, 14, 'sp4_v_b_38')
// (12, 15, 'sp4_v_b_27')
// (12, 16, 'sp4_v_b_14')
// (12, 17, 'sp4_v_b_3')
// (13, 10, 'sp4_h_r_28')
// (14, 10, 'sp4_h_r_41')
// (15, 10, 'sp4_h_l_41')

reg n1458 = 0;
// (10, 9, 'neigh_op_tnr_3')
// (10, 10, 'neigh_op_rgt_3')
// (10, 11, 'neigh_op_bnr_3')
// (11, 9, 'neigh_op_top_3')
// (11, 10, 'local_g1_3')
// (11, 10, 'lutff_1/in_1')
// (11, 10, 'lutff_3/out')
// (11, 11, 'neigh_op_bot_3')
// (12, 9, 'neigh_op_tnl_3')
// (12, 10, 'neigh_op_lft_3')
// (12, 11, 'neigh_op_bnl_3')

wire n1459;
// (10, 9, 'neigh_op_tnr_4')
// (10, 9, 'sp4_r_v_b_37')
// (10, 10, 'local_g2_4')
// (10, 10, 'lutff_7/in_3')
// (10, 10, 'neigh_op_rgt_4')
// (10, 10, 'sp4_r_v_b_24')
// (10, 10, 'sp4_r_v_b_40')
// (10, 11, 'local_g0_4')
// (10, 11, 'lutff_0/in_2')
// (10, 11, 'neigh_op_bnr_4')
// (10, 11, 'sp4_r_v_b_13')
// (10, 11, 'sp4_r_v_b_29')
// (10, 11, 'sp4_r_v_b_45')
// (10, 12, 'sp4_r_v_b_0')
// (10, 12, 'sp4_r_v_b_16')
// (10, 12, 'sp4_r_v_b_32')
// (10, 13, 'local_g1_5')
// (10, 13, 'lutff_3/in_3')
// (10, 13, 'lutff_4/in_2')
// (10, 13, 'lutff_6/in_2')
// (10, 13, 'sp4_r_v_b_21')
// (10, 13, 'sp4_r_v_b_37')
// (10, 13, 'sp4_r_v_b_38')
// (10, 13, 'sp4_r_v_b_5')
// (10, 14, 'local_g2_0')
// (10, 14, 'lutff_0/in_0')
// (10, 14, 'lutff_1/in_1')
// (10, 14, 'lutff_6/in_2')
// (10, 14, 'sp4_r_v_b_24')
// (10, 14, 'sp4_r_v_b_27')
// (10, 14, 'sp4_r_v_b_8')
// (10, 15, 'local_g2_5')
// (10, 15, 'lutff_0/in_3')
// (10, 15, 'sp4_r_v_b_13')
// (10, 15, 'sp4_r_v_b_14')
// (10, 16, 'local_g1_0')
// (10, 16, 'lutff_2/in_3')
// (10, 16, 'lutff_3/in_0')
// (10, 16, 'sp4_r_v_b_0')
// (10, 16, 'sp4_r_v_b_3')
// (11, 8, 'sp4_v_t_37')
// (11, 9, 'neigh_op_top_4')
// (11, 9, 'sp4_v_b_37')
// (11, 9, 'sp4_v_t_40')
// (11, 10, 'local_g2_4')
// (11, 10, 'lutff_3/in_1')
// (11, 10, 'lutff_4/out')
// (11, 10, 'lutff_7/in_1')
// (11, 10, 'sp4_h_r_8')
// (11, 10, 'sp4_v_b_24')
// (11, 10, 'sp4_v_b_40')
// (11, 10, 'sp4_v_t_45')
// (11, 11, 'neigh_op_bot_4')
// (11, 11, 'sp4_v_b_13')
// (11, 11, 'sp4_v_b_29')
// (11, 11, 'sp4_v_b_45')
// (11, 12, 'sp4_v_b_0')
// (11, 12, 'sp4_v_b_16')
// (11, 12, 'sp4_v_b_32')
// (11, 12, 'sp4_v_t_37')
// (11, 12, 'sp4_v_t_38')
// (11, 13, 'sp4_v_b_21')
// (11, 13, 'sp4_v_b_37')
// (11, 13, 'sp4_v_b_38')
// (11, 13, 'sp4_v_b_5')
// (11, 14, 'sp4_v_b_24')
// (11, 14, 'sp4_v_b_27')
// (11, 14, 'sp4_v_b_8')
// (11, 15, 'sp4_v_b_13')
// (11, 15, 'sp4_v_b_14')
// (11, 16, 'local_g0_0')
// (11, 16, 'local_g0_3')
// (11, 16, 'lutff_0/in_0')
// (11, 16, 'lutff_1/in_1')
// (11, 16, 'lutff_4/in_0')
// (11, 16, 'lutff_7/in_0')
// (11, 16, 'sp4_v_b_0')
// (11, 16, 'sp4_v_b_3')
// (12, 9, 'neigh_op_tnl_4')
// (12, 10, 'neigh_op_lft_4')
// (12, 10, 'sp4_h_r_21')
// (12, 11, 'neigh_op_bnl_4')
// (13, 10, 'sp4_h_r_32')
// (14, 10, 'sp4_h_r_45')
// (15, 10, 'sp4_h_l_45')

wire n1460;
// (10, 9, 'neigh_op_tnr_5')
// (10, 10, 'neigh_op_rgt_5')
// (10, 11, 'neigh_op_bnr_5')
// (11, 7, 'sp4_r_v_b_46')
// (11, 8, 'sp4_r_v_b_35')
// (11, 9, 'neigh_op_top_5')
// (11, 9, 'sp4_r_v_b_22')
// (11, 10, 'lutff_5/out')
// (11, 10, 'sp4_r_v_b_11')
// (11, 11, 'neigh_op_bot_5')
// (11, 11, 'sp4_r_v_b_46')
// (11, 12, 'sp4_r_v_b_35')
// (11, 13, 'sp4_r_v_b_22')
// (11, 14, 'local_g2_3')
// (11, 14, 'lutff_1/in_2')
// (11, 14, 'sp4_r_v_b_11')
// (12, 6, 'sp4_v_t_46')
// (12, 7, 'sp4_v_b_46')
// (12, 8, 'sp4_v_b_35')
// (12, 9, 'neigh_op_tnl_5')
// (12, 9, 'sp4_v_b_22')
// (12, 10, 'neigh_op_lft_5')
// (12, 10, 'sp4_v_b_11')
// (12, 10, 'sp4_v_t_46')
// (12, 11, 'neigh_op_bnl_5')
// (12, 11, 'sp4_v_b_46')
// (12, 12, 'sp4_v_b_35')
// (12, 13, 'sp4_v_b_22')
// (12, 14, 'sp4_v_b_11')

wire n1461;
// (10, 9, 'neigh_op_tnr_6')
// (10, 9, 'sp4_r_v_b_41')
// (10, 10, 'neigh_op_rgt_6')
// (10, 10, 'sp4_r_v_b_28')
// (10, 11, 'neigh_op_bnr_6')
// (10, 11, 'sp4_r_v_b_17')
// (10, 12, 'sp4_r_v_b_4')
// (10, 13, 'sp4_r_v_b_42')
// (10, 14, 'sp4_r_v_b_31')
// (10, 15, 'sp4_r_v_b_18')
// (10, 16, 'sp4_r_v_b_7')
// (11, 8, 'sp4_v_t_41')
// (11, 9, 'neigh_op_top_6')
// (11, 9, 'sp4_v_b_41')
// (11, 10, 'lutff_6/out')
// (11, 10, 'sp4_v_b_28')
// (11, 11, 'neigh_op_bot_6')
// (11, 11, 'sp4_v_b_17')
// (11, 12, 'sp4_v_b_4')
// (11, 12, 'sp4_v_t_42')
// (11, 13, 'local_g2_2')
// (11, 13, 'lutff_global/cen')
// (11, 13, 'sp4_v_b_42')
// (11, 14, 'sp4_v_b_31')
// (11, 15, 'sp4_v_b_18')
// (11, 16, 'sp4_v_b_7')
// (12, 9, 'neigh_op_tnl_6')
// (12, 10, 'neigh_op_lft_6')
// (12, 11, 'neigh_op_bnl_6')

reg n1462 = 0;
// (10, 9, 'neigh_op_tnr_7')
// (10, 10, 'neigh_op_rgt_7')
// (10, 10, 'sp4_r_v_b_46')
// (10, 11, 'neigh_op_bnr_7')
// (10, 11, 'sp4_r_v_b_35')
// (10, 12, 'local_g3_6')
// (10, 12, 'lutff_6/in_1')
// (10, 12, 'sp4_r_v_b_22')
// (10, 13, 'sp4_r_v_b_11')
// (11, 9, 'neigh_op_top_7')
// (11, 9, 'sp4_v_t_46')
// (11, 10, 'local_g3_7')
// (11, 10, 'lutff_5/in_3')
// (11, 10, 'lutff_7/out')
// (11, 10, 'sp4_v_b_46')
// (11, 11, 'neigh_op_bot_7')
// (11, 11, 'sp4_v_b_35')
// (11, 12, 'sp4_v_b_22')
// (11, 13, 'sp4_v_b_11')
// (12, 9, 'neigh_op_tnl_7')
// (12, 10, 'neigh_op_lft_7')
// (12, 11, 'neigh_op_bnl_7')

reg n1463 = 0;
// (10, 9, 'sp4_h_r_3')
// (11, 9, 'sp4_h_r_14')
// (12, 9, 'local_g2_3')
// (12, 9, 'lutff_7/in_2')
// (12, 9, 'sp4_h_r_27')
// (13, 9, 'neigh_op_tnr_3')
// (13, 9, 'sp4_h_r_38')
// (13, 10, 'neigh_op_rgt_3')
// (13, 10, 'sp4_r_v_b_38')
// (13, 11, 'neigh_op_bnr_3')
// (13, 11, 'sp4_r_v_b_27')
// (13, 11, 'sp4_r_v_b_43')
// (13, 12, 'sp4_r_v_b_14')
// (13, 12, 'sp4_r_v_b_30')
// (13, 13, 'sp4_r_v_b_19')
// (13, 13, 'sp4_r_v_b_3')
// (13, 14, 'sp4_r_v_b_6')
// (14, 3, 'sp4_r_v_b_42')
// (14, 4, 'sp4_r_v_b_31')
// (14, 5, 'sp4_r_v_b_18')
// (14, 6, 'sp4_r_v_b_7')
// (14, 7, 'sp4_r_v_b_42')
// (14, 8, 'sp4_r_v_b_31')
// (14, 9, 'neigh_op_top_3')
// (14, 9, 'sp4_h_l_38')
// (14, 9, 'sp4_r_v_b_18')
// (14, 9, 'sp4_v_t_38')
// (14, 10, 'lutff_3/out')
// (14, 10, 'sp4_h_r_6')
// (14, 10, 'sp4_r_v_b_7')
// (14, 10, 'sp4_v_b_38')
// (14, 10, 'sp4_v_t_43')
// (14, 11, 'local_g1_3')
// (14, 11, 'lutff_0/in_0')
// (14, 11, 'neigh_op_bot_3')
// (14, 11, 'sp4_v_b_27')
// (14, 11, 'sp4_v_b_43')
// (14, 12, 'sp4_v_b_14')
// (14, 12, 'sp4_v_b_30')
// (14, 13, 'sp4_h_r_9')
// (14, 13, 'sp4_v_b_19')
// (14, 13, 'sp4_v_b_3')
// (14, 14, 'local_g0_6')
// (14, 14, 'lutff_6/in_2')
// (14, 14, 'sp4_v_b_6')
// (15, 2, 'sp4_v_t_42')
// (15, 3, 'sp4_v_b_42')
// (15, 4, 'sp4_v_b_31')
// (15, 5, 'sp4_v_b_18')
// (15, 6, 'local_g0_7')
// (15, 6, 'lutff_2/in_1')
// (15, 6, 'sp4_h_r_7')
// (15, 6, 'sp4_v_b_7')
// (15, 6, 'sp4_v_t_42')
// (15, 7, 'sp4_v_b_42')
// (15, 8, 'sp4_v_b_31')
// (15, 9, 'neigh_op_tnl_3')
// (15, 9, 'sp4_v_b_18')
// (15, 10, 'neigh_op_lft_3')
// (15, 10, 'sp4_h_r_19')
// (15, 10, 'sp4_v_b_7')
// (15, 11, 'neigh_op_bnl_3')
// (15, 13, 'sp4_h_r_20')
// (16, 6, 'local_g1_2')
// (16, 6, 'lutff_6/in_1')
// (16, 6, 'sp4_h_r_18')
// (16, 10, 'sp4_h_r_30')
// (16, 13, 'local_g3_1')
// (16, 13, 'lutff_0/in_2')
// (16, 13, 'sp4_h_r_33')
// (17, 6, 'sp4_h_r_31')
// (17, 10, 'sp4_h_r_43')
// (17, 13, 'sp4_h_r_44')
// (18, 6, 'sp4_h_r_42')
// (18, 10, 'sp4_h_l_43')
// (18, 13, 'sp4_h_l_44')
// (19, 6, 'sp4_h_l_42')

reg n1464 = 0;
// (10, 9, 'sp4_r_v_b_36')
// (10, 10, 'local_g1_1')
// (10, 10, 'lutff_0/in_2')
// (10, 10, 'sp4_r_v_b_25')
// (10, 11, 'sp4_r_v_b_12')
// (10, 12, 'sp4_r_v_b_1')
// (10, 13, 'sp4_r_v_b_36')
// (10, 14, 'neigh_op_tnr_6')
// (10, 14, 'sp4_r_v_b_25')
// (10, 15, 'neigh_op_rgt_6')
// (10, 15, 'sp4_r_v_b_12')
// (10, 16, 'neigh_op_bnr_6')
// (10, 16, 'sp4_r_v_b_1')
// (11, 8, 'sp4_v_t_36')
// (11, 9, 'sp4_v_b_36')
// (11, 10, 'sp4_v_b_25')
// (11, 11, 'sp4_v_b_12')
// (11, 12, 'sp4_v_b_1')
// (11, 12, 'sp4_v_t_36')
// (11, 13, 'sp4_v_b_36')
// (11, 14, 'local_g0_6')
// (11, 14, 'lutff_7/in_3')
// (11, 14, 'neigh_op_top_6')
// (11, 14, 'sp4_v_b_25')
// (11, 15, 'local_g3_6')
// (11, 15, 'lutff_6/in_1')
// (11, 15, 'lutff_6/out')
// (11, 15, 'sp4_v_b_12')
// (11, 16, 'neigh_op_bot_6')
// (11, 16, 'sp4_v_b_1')
// (12, 14, 'neigh_op_tnl_6')
// (12, 15, 'neigh_op_lft_6')
// (12, 16, 'neigh_op_bnl_6')

reg n1465 = 0;
// (10, 9, 'sp4_r_v_b_46')
// (10, 10, 'sp4_r_v_b_35')
// (10, 11, 'sp4_r_v_b_22')
// (10, 12, 'neigh_op_tnr_7')
// (10, 12, 'sp4_r_v_b_11')
// (10, 13, 'neigh_op_rgt_7')
// (10, 13, 'sp4_r_v_b_46')
// (10, 14, 'neigh_op_bnr_7')
// (10, 14, 'sp4_r_v_b_35')
// (10, 15, 'local_g3_6')
// (10, 15, 'lutff_0/in_1')
// (10, 15, 'sp4_r_v_b_22')
// (10, 16, 'sp4_r_v_b_11')
// (11, 8, 'sp4_h_r_11')
// (11, 8, 'sp4_v_t_46')
// (11, 9, 'sp4_v_b_46')
// (11, 10, 'sp4_v_b_35')
// (11, 11, 'sp4_v_b_22')
// (11, 12, 'neigh_op_top_7')
// (11, 12, 'sp4_h_r_11')
// (11, 12, 'sp4_v_b_11')
// (11, 12, 'sp4_v_t_46')
// (11, 13, 'lutff_7/out')
// (11, 13, 'sp4_v_b_46')
// (11, 14, 'neigh_op_bot_7')
// (11, 14, 'sp4_v_b_35')
// (11, 15, 'sp4_v_b_22')
// (11, 16, 'sp4_v_b_11')
// (12, 8, 'sp4_h_r_22')
// (12, 12, 'neigh_op_tnl_7')
// (12, 12, 'sp4_h_r_22')
// (12, 13, 'neigh_op_lft_7')
// (12, 14, 'neigh_op_bnl_7')
// (13, 8, 'local_g2_3')
// (13, 8, 'lutff_1/in_2')
// (13, 8, 'lutff_6/in_1')
// (13, 8, 'sp4_h_r_35')
// (13, 12, 'sp4_h_r_35')
// (14, 8, 'sp4_h_r_46')
// (14, 9, 'sp4_r_v_b_40')
// (14, 10, 'sp4_r_v_b_29')
// (14, 11, 'sp4_r_v_b_16')
// (14, 12, 'sp4_h_r_46')
// (14, 12, 'sp4_r_v_b_5')
// (15, 8, 'sp4_h_l_46')
// (15, 8, 'sp4_v_t_40')
// (15, 9, 'local_g2_0')
// (15, 9, 'lutff_1/in_1')
// (15, 9, 'lutff_2/in_2')
// (15, 9, 'sp4_v_b_40')
// (15, 10, 'sp4_v_b_29')
// (15, 11, 'sp4_v_b_16')
// (15, 12, 'sp4_h_l_46')
// (15, 12, 'sp4_v_b_5')

wire n1466;
// (10, 10, 'neigh_op_tnr_2')
// (10, 11, 'neigh_op_rgt_2')
// (10, 12, 'neigh_op_bnr_2')
// (11, 10, 'neigh_op_top_2')
// (11, 11, 'lutff_2/out')
// (11, 12, 'neigh_op_bot_2')
// (12, 10, 'neigh_op_tnl_2')
// (12, 11, 'local_g1_2')
// (12, 11, 'lutff_7/in_2')
// (12, 11, 'neigh_op_lft_2')
// (12, 12, 'neigh_op_bnl_2')

wire n1467;
// (10, 10, 'neigh_op_tnr_4')
// (10, 11, 'neigh_op_rgt_4')
// (10, 12, 'neigh_op_bnr_4')
// (11, 10, 'neigh_op_top_4')
// (11, 11, 'lutff_4/out')
// (11, 11, 'sp4_r_v_b_41')
// (11, 12, 'neigh_op_bot_4')
// (11, 12, 'sp4_r_v_b_28')
// (11, 13, 'sp4_r_v_b_17')
// (11, 14, 'sp4_r_v_b_4')
// (12, 10, 'neigh_op_tnl_4')
// (12, 10, 'sp4_v_t_41')
// (12, 11, 'neigh_op_lft_4')
// (12, 11, 'sp4_v_b_41')
// (12, 12, 'neigh_op_bnl_4')
// (12, 12, 'sp4_v_b_28')
// (12, 13, 'sp4_v_b_17')
// (12, 14, 'local_g0_4')
// (12, 14, 'lutff_4/in_2')
// (12, 14, 'sp4_v_b_4')

reg n1468 = 0;
// (10, 10, 'neigh_op_tnr_5')
// (10, 11, 'neigh_op_rgt_5')
// (10, 12, 'neigh_op_bnr_5')
// (11, 10, 'local_g0_5')
// (11, 10, 'lutff_5/in_2')
// (11, 10, 'neigh_op_top_5')
// (11, 11, 'lutff_5/out')
// (11, 12, 'neigh_op_bot_5')
// (12, 10, 'neigh_op_tnl_5')
// (12, 11, 'neigh_op_lft_5')
// (12, 12, 'neigh_op_bnl_5')

reg n1469 = 0;
// (10, 10, 'sp4_r_v_b_37')
// (10, 11, 'sp4_r_v_b_24')
// (10, 12, 'sp4_r_v_b_13')
// (10, 13, 'sp4_r_v_b_0')
// (10, 14, 'sp4_r_v_b_37')
// (10, 15, 'sp4_r_v_b_24')
// (10, 16, 'neigh_op_tnr_0')
// (10, 16, 'sp4_r_v_b_13')
// (10, 17, 'neigh_op_rgt_0')
// (10, 17, 'sp4_r_v_b_0')
// (10, 18, 'neigh_op_bnr_0')
// (11, 9, 'sp4_v_t_37')
// (11, 10, 'local_g3_5')
// (11, 10, 'lutff_0/in_0')
// (11, 10, 'sp4_v_b_37')
// (11, 11, 'sp4_v_b_24')
// (11, 12, 'sp4_v_b_13')
// (11, 13, 'sp4_v_b_0')
// (11, 13, 'sp4_v_t_37')
// (11, 14, 'sp4_v_b_37')
// (11, 15, 'sp4_v_b_24')
// (11, 16, 'neigh_op_top_0')
// (11, 16, 'sp4_v_b_13')
// (11, 17, 'local_g3_0')
// (11, 17, 'lutff_0/out')
// (11, 17, 'lutff_2/in_1')
// (11, 17, 'sp4_v_b_0')
// (11, 18, 'neigh_op_bot_0')
// (12, 16, 'neigh_op_tnl_0')
// (12, 17, 'neigh_op_lft_0')
// (12, 18, 'neigh_op_bnl_0')

reg n1470 = 0;
// (10, 10, 'sp4_r_v_b_41')
// (10, 11, 'sp4_r_v_b_28')
// (10, 12, 'local_g3_1')
// (10, 12, 'lutff_5/in_1')
// (10, 12, 'sp4_r_v_b_17')
// (10, 13, 'sp4_r_v_b_4')
// (11, 9, 'sp4_v_t_41')
// (11, 10, 'sp4_v_b_41')
// (11, 11, 'sp4_v_b_28')
// (11, 12, 'neigh_op_tnr_3')
// (11, 12, 'sp4_v_b_17')
// (11, 13, 'neigh_op_rgt_3')
// (11, 13, 'sp4_h_r_11')
// (11, 13, 'sp4_v_b_4')
// (11, 14, 'neigh_op_bnr_3')
// (12, 12, 'neigh_op_top_3')
// (12, 13, 'lutff_3/out')
// (12, 13, 'sp4_h_r_22')
// (12, 14, 'neigh_op_bot_3')
// (13, 12, 'neigh_op_tnl_3')
// (13, 13, 'neigh_op_lft_3')
// (13, 13, 'sp4_h_r_35')
// (13, 14, 'neigh_op_bnl_3')
// (14, 13, 'sp4_h_r_46')
// (15, 13, 'sp4_h_l_46')

wire n1471;
// (10, 11, 'local_g3_4')
// (10, 11, 'lutff_0/in_3')
// (10, 11, 'lutff_2/in_3')
// (10, 11, 'neigh_op_tnr_4')
// (10, 12, 'neigh_op_rgt_4')
// (10, 13, 'local_g1_4')
// (10, 13, 'lutff_3/in_2')
// (10, 13, 'neigh_op_bnr_4')
// (11, 11, 'local_g1_4')
// (11, 11, 'lutff_5/in_2')
// (11, 11, 'neigh_op_top_4')
// (11, 12, 'lutff_4/out')
// (11, 13, 'neigh_op_bot_4')
// (12, 11, 'neigh_op_tnl_4')
// (12, 12, 'neigh_op_lft_4')
// (12, 13, 'neigh_op_bnl_4')

wire n1472;
// (10, 11, 'neigh_op_tnr_1')
// (10, 12, 'neigh_op_rgt_1')
// (10, 13, 'neigh_op_bnr_1')
// (11, 11, 'neigh_op_top_1')
// (11, 12, 'local_g0_1')
// (11, 12, 'lutff_1/out')
// (11, 12, 'lutff_5/in_0')
// (11, 13, 'neigh_op_bot_1')
// (12, 11, 'neigh_op_tnl_1')
// (12, 12, 'neigh_op_lft_1')
// (12, 13, 'neigh_op_bnl_1')

reg n1473 = 0;
// (10, 11, 'neigh_op_tnr_3')
// (10, 12, 'local_g3_3')
// (10, 12, 'lutff_2/in_0')
// (10, 12, 'neigh_op_rgt_3')
// (10, 13, 'neigh_op_bnr_3')
// (11, 11, 'local_g1_3')
// (11, 11, 'lutff_1/in_1')
// (11, 11, 'neigh_op_top_3')
// (11, 12, 'local_g1_3')
// (11, 12, 'lutff_0/in_2')
// (11, 12, 'lutff_1/in_1')
// (11, 12, 'lutff_3/out')
// (11, 12, 'sp4_h_r_6')
// (11, 13, 'neigh_op_bot_3')
// (12, 11, 'neigh_op_tnl_3')
// (12, 12, 'local_g0_3')
// (12, 12, 'lutff_4/in_1')
// (12, 12, 'neigh_op_lft_3')
// (12, 12, 'sp4_h_r_19')
// (12, 13, 'neigh_op_bnl_3')
// (13, 12, 'sp4_h_r_30')
// (14, 9, 'sp4_r_v_b_42')
// (14, 10, 'sp4_r_v_b_31')
// (14, 11, 'sp4_r_v_b_18')
// (14, 12, 'sp4_h_r_43')
// (14, 12, 'sp4_r_v_b_7')
// (14, 13, 'sp4_r_v_b_46')
// (14, 14, 'sp4_r_v_b_35')
// (14, 15, 'sp4_r_v_b_22')
// (14, 16, 'sp4_r_v_b_11')
// (15, 8, 'sp4_v_t_42')
// (15, 9, 'sp4_v_b_42')
// (15, 10, 'sp4_v_b_31')
// (15, 11, 'local_g0_2')
// (15, 11, 'lutff_0/in_2')
// (15, 11, 'lutff_4/in_2')
// (15, 11, 'sp4_v_b_18')
// (15, 12, 'sp4_h_l_43')
// (15, 12, 'sp4_h_r_2')
// (15, 12, 'sp4_v_b_7')
// (15, 12, 'sp4_v_t_46')
// (15, 13, 'sp4_v_b_46')
// (15, 14, 'local_g2_3')
// (15, 14, 'lutff_7/in_2')
// (15, 14, 'sp4_v_b_35')
// (15, 15, 'sp4_v_b_22')
// (15, 16, 'sp4_v_b_11')
// (16, 12, 'sp4_h_r_15')
// (17, 12, 'sp4_h_r_26')
// (18, 12, 'sp4_h_r_39')
// (19, 12, 'sp4_h_l_39')

reg n1474 = 0;
// (10, 11, 'neigh_op_tnr_6')
// (10, 12, 'neigh_op_rgt_6')
// (10, 13, 'neigh_op_bnr_6')
// (11, 11, 'local_g0_6')
// (11, 11, 'lutff_0/in_2')
// (11, 11, 'neigh_op_top_6')
// (11, 11, 'sp4_r_v_b_40')
// (11, 12, 'local_g0_6')
// (11, 12, 'lutff_1/in_3')
// (11, 12, 'lutff_3/in_3')
// (11, 12, 'lutff_6/out')
// (11, 12, 'sp4_r_v_b_29')
// (11, 13, 'neigh_op_bot_6')
// (11, 13, 'sp4_r_v_b_16')
// (11, 14, 'sp4_r_v_b_5')
// (12, 10, 'sp4_h_r_10')
// (12, 10, 'sp4_v_t_40')
// (12, 11, 'neigh_op_tnl_6')
// (12, 11, 'sp4_v_b_40')
// (12, 12, 'local_g0_6')
// (12, 12, 'lutff_4/in_0')
// (12, 12, 'lutff_7/in_1')
// (12, 12, 'neigh_op_lft_6')
// (12, 12, 'sp4_v_b_29')
// (12, 13, 'neigh_op_bnl_6')
// (12, 13, 'sp4_v_b_16')
// (12, 14, 'sp4_h_r_11')
// (12, 14, 'sp4_h_r_5')
// (12, 14, 'sp4_v_b_5')
// (13, 10, 'sp4_h_r_23')
// (13, 14, 'local_g1_6')
// (13, 14, 'lutff_4/in_1')
// (13, 14, 'sp4_h_r_16')
// (13, 14, 'sp4_h_r_22')
// (14, 10, 'sp4_h_r_34')
// (14, 14, 'sp4_h_r_29')
// (14, 14, 'sp4_h_r_35')
// (15, 10, 'local_g3_7')
// (15, 10, 'lutff_5/in_1')
// (15, 10, 'sp4_h_r_47')
// (15, 11, 'sp4_r_v_b_46')
// (15, 12, 'sp4_r_v_b_35')
// (15, 13, 'local_g3_6')
// (15, 13, 'lutff_1/in_0')
// (15, 13, 'sp4_r_v_b_22')
// (15, 14, 'sp4_h_r_40')
// (15, 14, 'sp4_h_r_46')
// (15, 14, 'sp4_r_v_b_11')
// (16, 10, 'sp4_h_l_47')
// (16, 10, 'sp4_v_t_46')
// (16, 11, 'sp4_v_b_46')
// (16, 12, 'sp4_v_b_35')
// (16, 13, 'sp4_v_b_22')
// (16, 14, 'sp4_h_l_40')
// (16, 14, 'sp4_h_l_46')
// (16, 14, 'sp4_v_b_11')

wire n1475;
// (10, 11, 'sp4_h_r_8')
// (11, 11, 'local_g1_5')
// (11, 11, 'lutff_4/in_2')
// (11, 11, 'sp4_h_r_21')
// (11, 12, 'local_g1_4')
// (11, 12, 'lutff_5/in_2')
// (11, 12, 'sp4_h_r_4')
// (12, 11, 'local_g3_6')
// (12, 11, 'lutff_7/in_0')
// (12, 11, 'neigh_op_tnr_6')
// (12, 11, 'sp4_h_r_32')
// (12, 12, 'local_g2_6')
// (12, 12, 'lutff_4/in_2')
// (12, 12, 'lutff_6/in_0')
// (12, 12, 'neigh_op_rgt_6')
// (12, 12, 'sp4_h_r_17')
// (12, 13, 'neigh_op_bnr_6')
// (13, 11, 'neigh_op_top_6')
// (13, 11, 'sp4_h_r_45')
// (13, 12, 'lutff_6/out')
// (13, 12, 'sp4_h_r_28')
// (13, 12, 'sp4_r_v_b_45')
// (13, 13, 'neigh_op_bot_6')
// (13, 13, 'sp4_r_v_b_32')
// (13, 14, 'sp4_r_v_b_21')
// (13, 15, 'sp4_r_v_b_8')
// (14, 11, 'neigh_op_tnl_6')
// (14, 11, 'sp4_h_l_45')
// (14, 11, 'sp4_v_t_45')
// (14, 12, 'neigh_op_lft_6')
// (14, 12, 'sp4_h_r_41')
// (14, 12, 'sp4_v_b_45')
// (14, 13, 'neigh_op_bnl_6')
// (14, 13, 'sp4_v_b_32')
// (14, 14, 'sp4_v_b_21')
// (14, 15, 'sp4_v_b_8')
// (15, 12, 'sp4_h_l_41')

wire n1476;
// (10, 12, 'neigh_op_tnr_5')
// (10, 13, 'neigh_op_rgt_5')
// (10, 14, 'neigh_op_bnr_5')
// (11, 12, 'neigh_op_top_5')
// (11, 12, 'sp4_r_v_b_38')
// (11, 13, 'lutff_5/out')
// (11, 13, 'sp4_r_v_b_27')
// (11, 14, 'neigh_op_bot_5')
// (11, 14, 'sp4_r_v_b_14')
// (11, 15, 'sp4_r_v_b_3')
// (12, 11, 'sp4_v_t_38')
// (12, 12, 'neigh_op_tnl_5')
// (12, 12, 'sp4_v_b_38')
// (12, 13, 'neigh_op_lft_5')
// (12, 13, 'sp4_v_b_27')
// (12, 14, 'neigh_op_bnl_5')
// (12, 14, 'sp4_v_b_14')
// (12, 15, 'local_g0_3')
// (12, 15, 'lutff_1/in_0')
// (12, 15, 'sp4_v_b_3')

reg n1477 = 0;
// (10, 12, 'sp4_r_v_b_36')
// (10, 13, 'sp4_r_v_b_25')
// (10, 14, 'local_g2_4')
// (10, 14, 'lutff_1/in_3')
// (10, 14, 'sp4_r_v_b_12')
// (10, 15, 'local_g1_1')
// (10, 15, 'lutff_4/in_0')
// (10, 15, 'sp4_r_v_b_1')
// (10, 16, 'sp4_r_v_b_47')
// (10, 17, 'sp4_r_v_b_34')
// (10, 18, 'neigh_op_tnr_5')
// (10, 18, 'sp4_r_v_b_23')
// (10, 19, 'neigh_op_rgt_5')
// (10, 19, 'sp4_r_v_b_10')
// (10, 20, 'neigh_op_bnr_5')
// (11, 11, 'sp4_v_t_36')
// (11, 12, 'sp4_r_v_b_39')
// (11, 12, 'sp4_v_b_36')
// (11, 13, 'sp4_r_v_b_26')
// (11, 13, 'sp4_v_b_25')
// (11, 14, 'sp4_r_v_b_15')
// (11, 14, 'sp4_v_b_12')
// (11, 15, 'sp4_r_v_b_2')
// (11, 15, 'sp4_v_b_1')
// (11, 15, 'sp4_v_t_47')
// (11, 16, 'sp4_r_v_b_46')
// (11, 16, 'sp4_v_b_47')
// (11, 17, 'sp4_r_v_b_35')
// (11, 17, 'sp4_v_b_34')
// (11, 18, 'local_g0_5')
// (11, 18, 'lutff_1/in_0')
// (11, 18, 'neigh_op_top_5')
// (11, 18, 'sp4_r_v_b_22')
// (11, 18, 'sp4_v_b_23')
// (11, 19, 'local_g2_5')
// (11, 19, 'lutff_5/in_0')
// (11, 19, 'lutff_5/out')
// (11, 19, 'sp4_r_v_b_11')
// (11, 19, 'sp4_v_b_10')
// (11, 20, 'neigh_op_bot_5')
// (12, 11, 'local_g0_7')
// (12, 11, 'lutff_0/in_1')
// (12, 11, 'sp4_h_r_7')
// (12, 11, 'sp4_v_t_39')
// (12, 12, 'sp4_v_b_39')
// (12, 13, 'sp4_v_b_26')
// (12, 14, 'sp4_v_b_15')
// (12, 15, 'sp4_v_b_2')
// (12, 15, 'sp4_v_t_46')
// (12, 16, 'sp4_v_b_46')
// (12, 17, 'sp4_v_b_35')
// (12, 18, 'neigh_op_tnl_5')
// (12, 18, 'sp4_v_b_22')
// (12, 19, 'neigh_op_lft_5')
// (12, 19, 'sp4_v_b_11')
// (12, 20, 'neigh_op_bnl_5')
// (13, 11, 'sp4_h_r_18')
// (14, 11, 'sp4_h_r_31')
// (15, 11, 'sp4_h_r_42')
// (16, 11, 'sp4_h_l_42')

wire n1478;
// (10, 12, 'sp4_r_v_b_45')
// (10, 13, 'sp4_r_v_b_32')
// (10, 14, 'sp4_r_v_b_21')
// (10, 15, 'sp4_r_v_b_8')
// (10, 16, 'sp4_h_r_11')
// (11, 11, 'sp4_v_t_45')
// (11, 12, 'sp4_v_b_45')
// (11, 13, 'sp4_v_b_32')
// (11, 14, 'local_g1_5')
// (11, 14, 'lutff_2/in_2')
// (11, 14, 'sp4_v_b_21')
// (11, 15, 'sp4_h_r_3')
// (11, 15, 'sp4_v_b_8')
// (11, 16, 'local_g0_6')
// (11, 16, 'lutff_6/in_0')
// (11, 16, 'lutff_7/in_1')
// (11, 16, 'sp4_h_r_22')
// (12, 15, 'sp4_h_r_14')
// (12, 16, 'sp4_h_r_35')
// (13, 1, 'sp4_r_v_b_29')
// (13, 2, 'local_g3_0')
// (13, 2, 'lutff_4/in_3')
// (13, 2, 'sp4_r_v_b_16')
// (13, 3, 'sp4_r_v_b_5')
// (13, 4, 'sp4_r_v_b_40')
// (13, 5, 'sp4_r_v_b_29')
// (13, 6, 'sp4_r_v_b_16')
// (13, 7, 'sp4_r_v_b_5')
// (13, 8, 'sp4_r_v_b_44')
// (13, 9, 'sp4_r_v_b_33')
// (13, 10, 'sp4_r_v_b_20')
// (13, 11, 'sp4_r_v_b_9')
// (13, 12, 'sp4_r_v_b_43')
// (13, 13, 'sp4_r_v_b_30')
// (13, 13, 'sp4_r_v_b_46')
// (13, 14, 'neigh_op_tnr_3')
// (13, 14, 'sp4_r_v_b_19')
// (13, 14, 'sp4_r_v_b_35')
// (13, 15, 'neigh_op_rgt_3')
// (13, 15, 'sp4_h_r_27')
// (13, 15, 'sp4_r_v_b_22')
// (13, 15, 'sp4_r_v_b_6')
// (13, 16, 'neigh_op_bnr_3')
// (13, 16, 'sp4_h_r_46')
// (13, 16, 'sp4_r_v_b_11')
// (14, 0, 'span4_vert_29')
// (14, 1, 'sp4_v_b_29')
// (14, 2, 'sp4_v_b_16')
// (14, 3, 'sp4_v_b_5')
// (14, 3, 'sp4_v_t_40')
// (14, 4, 'sp4_v_b_40')
// (14, 5, 'sp4_v_b_29')
// (14, 6, 'sp4_v_b_16')
// (14, 7, 'sp4_v_b_5')
// (14, 7, 'sp4_v_t_44')
// (14, 8, 'sp4_v_b_44')
// (14, 9, 'sp4_v_b_33')
// (14, 10, 'sp4_v_b_20')
// (14, 11, 'sp4_v_b_9')
// (14, 11, 'sp4_v_t_43')
// (14, 12, 'sp4_v_b_43')
// (14, 12, 'sp4_v_t_46')
// (14, 13, 'sp4_v_b_30')
// (14, 13, 'sp4_v_b_46')
// (14, 14, 'neigh_op_top_3')
// (14, 14, 'sp4_v_b_19')
// (14, 14, 'sp4_v_b_35')
// (14, 15, 'lutff_3/out')
// (14, 15, 'sp4_h_r_38')
// (14, 15, 'sp4_v_b_22')
// (14, 15, 'sp4_v_b_6')
// (14, 16, 'neigh_op_bot_3')
// (14, 16, 'sp4_h_l_46')
// (14, 16, 'sp4_v_b_11')
// (15, 14, 'neigh_op_tnl_3')
// (15, 15, 'neigh_op_lft_3')
// (15, 15, 'sp4_h_l_38')
// (15, 16, 'neigh_op_bnl_3')

reg n1479 = 0;
// (10, 12, 'sp4_r_v_b_47')
// (10, 13, 'local_g2_2')
// (10, 13, 'lutff_2/in_0')
// (10, 13, 'sp4_r_v_b_34')
// (10, 14, 'sp4_r_v_b_23')
// (10, 15, 'sp4_r_v_b_10')
// (10, 16, 'neigh_op_tnr_5')
// (10, 16, 'sp4_r_v_b_39')
// (10, 17, 'neigh_op_rgt_5')
// (10, 17, 'sp4_r_v_b_26')
// (10, 18, 'neigh_op_bnr_5')
// (10, 18, 'sp4_r_v_b_15')
// (10, 19, 'sp4_r_v_b_2')
// (11, 11, 'sp4_v_t_47')
// (11, 12, 'sp4_v_b_47')
// (11, 13, 'sp4_v_b_34')
// (11, 14, 'sp4_v_b_23')
// (11, 15, 'sp4_v_b_10')
// (11, 15, 'sp4_v_t_39')
// (11, 16, 'neigh_op_top_5')
// (11, 16, 'sp4_v_b_39')
// (11, 17, 'local_g2_5')
// (11, 17, 'lutff_5/out')
// (11, 17, 'lutff_6/in_3')
// (11, 17, 'sp4_v_b_26')
// (11, 18, 'neigh_op_bot_5')
// (11, 18, 'sp4_v_b_15')
// (11, 19, 'sp4_v_b_2')
// (12, 16, 'neigh_op_tnl_5')
// (12, 17, 'neigh_op_lft_5')
// (12, 18, 'neigh_op_bnl_5')

reg n1480 = 0;
// (10, 13, 'neigh_op_tnr_1')
// (10, 13, 'sp4_r_v_b_47')
// (10, 14, 'neigh_op_rgt_1')
// (10, 14, 'sp4_r_v_b_34')
// (10, 15, 'neigh_op_bnr_1')
// (10, 15, 'sp4_r_v_b_23')
// (10, 16, 'sp4_r_v_b_10')
// (11, 12, 'sp4_v_t_47')
// (11, 13, 'neigh_op_top_1')
// (11, 13, 'sp4_v_b_47')
// (11, 14, 'lutff_1/out')
// (11, 14, 'sp4_v_b_34')
// (11, 15, 'neigh_op_bot_1')
// (11, 15, 'sp4_v_b_23')
// (11, 16, 'sp4_h_r_10')
// (11, 16, 'sp4_v_b_10')
// (12, 13, 'neigh_op_tnl_1')
// (12, 14, 'neigh_op_lft_1')
// (12, 15, 'neigh_op_bnl_1')
// (12, 16, 'sp4_h_r_23')
// (13, 16, 'sp4_h_r_34')
// (14, 16, 'sp4_h_r_47')
// (15, 16, 'sp4_h_l_47')
// (15, 16, 'sp4_h_r_10')
// (16, 16, 'sp4_h_r_23')
// (17, 16, 'local_g2_2')
// (17, 16, 'lutff_6/in_0')
// (17, 16, 'sp4_h_r_34')
// (18, 16, 'sp4_h_r_47')
// (19, 16, 'sp4_h_l_47')

wire n1481;
// (10, 13, 'neigh_op_tnr_3')
// (10, 14, 'neigh_op_rgt_3')
// (10, 15, 'neigh_op_bnr_3')
// (11, 13, 'neigh_op_top_3')
// (11, 14, 'lutff_3/out')
// (11, 15, 'local_g0_3')
// (11, 15, 'lutff_7/in_2')
// (11, 15, 'neigh_op_bot_3')
// (12, 13, 'neigh_op_tnl_3')
// (12, 14, 'neigh_op_lft_3')
// (12, 15, 'neigh_op_bnl_3')

reg n1482 = 0;
// (10, 13, 'neigh_op_tnr_4')
// (10, 14, 'neigh_op_rgt_4')
// (10, 15, 'neigh_op_bnr_4')
// (11, 13, 'neigh_op_top_4')
// (11, 13, 'sp4_r_v_b_36')
// (11, 14, 'lutff_4/out')
// (11, 14, 'sp4_r_v_b_25')
// (11, 15, 'neigh_op_bot_4')
// (11, 15, 'sp4_r_v_b_12')
// (11, 16, 'sp4_r_v_b_1')
// (12, 12, 'sp4_v_t_36')
// (12, 13, 'neigh_op_tnl_4')
// (12, 13, 'sp4_v_b_36')
// (12, 14, 'neigh_op_lft_4')
// (12, 14, 'sp4_v_b_25')
// (12, 15, 'neigh_op_bnl_4')
// (12, 15, 'sp4_v_b_12')
// (12, 16, 'sp4_h_r_7')
// (12, 16, 'sp4_v_b_1')
// (13, 16, 'sp4_h_r_18')
// (14, 16, 'sp4_h_r_31')
// (15, 13, 'sp4_r_v_b_36')
// (15, 14, 'sp4_r_v_b_25')
// (15, 15, 'sp4_r_v_b_12')
// (15, 16, 'sp4_h_r_42')
// (15, 16, 'sp4_r_v_b_1')
// (16, 12, 'sp4_v_t_36')
// (16, 13, 'sp4_v_b_36')
// (16, 14, 'sp4_v_b_25')
// (16, 15, 'local_g1_4')
// (16, 15, 'lutff_6/in_1')
// (16, 15, 'sp4_v_b_12')
// (16, 16, 'sp4_h_l_42')
// (16, 16, 'sp4_v_b_1')

wire n1483;
// (10, 13, 'neigh_op_tnr_5')
// (10, 14, 'neigh_op_rgt_5')
// (10, 15, 'neigh_op_bnr_5')
// (11, 13, 'neigh_op_top_5')
// (11, 13, 'sp4_r_v_b_38')
// (11, 14, 'lutff_5/out')
// (11, 14, 'sp4_r_v_b_27')
// (11, 14, 'sp4_r_v_b_43')
// (11, 15, 'local_g1_5')
// (11, 15, 'lutff_1/in_3')
// (11, 15, 'neigh_op_bot_5')
// (11, 15, 'sp4_r_v_b_14')
// (11, 15, 'sp4_r_v_b_30')
// (11, 16, 'sp4_r_v_b_19')
// (11, 16, 'sp4_r_v_b_3')
// (11, 17, 'sp4_r_v_b_6')
// (12, 12, 'sp4_v_t_38')
// (12, 13, 'neigh_op_tnl_5')
// (12, 13, 'sp4_v_b_38')
// (12, 13, 'sp4_v_t_43')
// (12, 14, 'neigh_op_lft_5')
// (12, 14, 'sp4_v_b_27')
// (12, 14, 'sp4_v_b_43')
// (12, 15, 'neigh_op_bnl_5')
// (12, 15, 'sp4_v_b_14')
// (12, 15, 'sp4_v_b_30')
// (12, 16, 'local_g0_3')
// (12, 16, 'lutff_2/in_3')
// (12, 16, 'sp4_v_b_19')
// (12, 16, 'sp4_v_b_3')
// (12, 17, 'local_g0_6')
// (12, 17, 'lutff_2/in_0')
// (12, 17, 'sp4_v_b_6')

wire n1484;
// (10, 13, 'neigh_op_tnr_6')
// (10, 14, 'neigh_op_rgt_6')
// (10, 15, 'neigh_op_bnr_6')
// (11, 13, 'neigh_op_top_6')
// (11, 14, 'local_g1_6')
// (11, 14, 'lutff_4/in_3')
// (11, 14, 'lutff_6/out')
// (11, 15, 'neigh_op_bot_6')
// (12, 13, 'neigh_op_tnl_6')
// (12, 14, 'neigh_op_lft_6')
// (12, 15, 'neigh_op_bnl_6')

wire n1485;
// (10, 13, 'neigh_op_tnr_7')
// (10, 14, 'neigh_op_rgt_7')
// (10, 15, 'neigh_op_bnr_7')
// (11, 13, 'neigh_op_top_7')
// (11, 14, 'lutff_7/out')
// (11, 14, 'sp4_r_v_b_47')
// (11, 15, 'neigh_op_bot_7')
// (11, 15, 'sp4_r_v_b_34')
// (11, 16, 'sp4_r_v_b_23')
// (11, 17, 'sp4_r_v_b_10')
// (12, 13, 'neigh_op_tnl_7')
// (12, 13, 'sp4_v_t_47')
// (12, 14, 'neigh_op_lft_7')
// (12, 14, 'sp4_v_b_47')
// (12, 15, 'neigh_op_bnl_7')
// (12, 15, 'sp4_v_b_34')
// (12, 16, 'sp4_v_b_23')
// (12, 17, 'local_g1_2')
// (12, 17, 'lutff_2/in_3')
// (12, 17, 'sp4_v_b_10')

reg n1486 = 0;
// (10, 13, 'sp4_r_v_b_43')
// (10, 14, 'sp4_r_v_b_30')
// (10, 15, 'neigh_op_tnr_3')
// (10, 15, 'sp4_r_v_b_19')
// (10, 16, 'neigh_op_rgt_3')
// (10, 16, 'sp4_r_v_b_6')
// (10, 17, 'neigh_op_bnr_3')
// (11, 12, 'sp4_v_t_43')
// (11, 13, 'sp4_v_b_43')
// (11, 14, 'local_g2_6')
// (11, 14, 'lutff_3/in_3')
// (11, 14, 'sp4_v_b_30')
// (11, 15, 'neigh_op_top_3')
// (11, 15, 'sp4_v_b_19')
// (11, 16, 'lutff_3/out')
// (11, 16, 'sp4_v_b_6')
// (11, 17, 'neigh_op_bot_3')
// (12, 15, 'neigh_op_tnl_3')
// (12, 16, 'neigh_op_lft_3')
// (12, 17, 'neigh_op_bnl_3')

reg n1487 = 0;
// (10, 14, 'local_g3_0')
// (10, 14, 'lutff_7/in_2')
// (10, 14, 'neigh_op_tnr_0')
// (10, 15, 'neigh_op_rgt_0')
// (10, 16, 'neigh_op_bnr_0')
// (11, 14, 'local_g1_0')
// (11, 14, 'lutff_7/in_2')
// (11, 14, 'neigh_op_top_0')
// (11, 15, 'local_g3_0')
// (11, 15, 'lutff_0/in_1')
// (11, 15, 'lutff_0/out')
// (11, 16, 'neigh_op_bot_0')
// (12, 14, 'neigh_op_tnl_0')
// (12, 15, 'neigh_op_lft_0')
// (12, 16, 'neigh_op_bnl_0')

reg n1488 = 0;
// (10, 14, 'neigh_op_tnr_1')
// (10, 15, 'local_g2_1')
// (10, 15, 'lutff_2/in_1')
// (10, 15, 'neigh_op_rgt_1')
// (10, 16, 'neigh_op_bnr_1')
// (11, 14, 'neigh_op_top_1')
// (11, 14, 'sp4_r_v_b_46')
// (11, 15, 'local_g0_1')
// (11, 15, 'lutff_1/in_2')
// (11, 15, 'lutff_1/out')
// (11, 15, 'sp4_r_v_b_35')
// (11, 16, 'neigh_op_bot_1')
// (11, 16, 'sp4_r_v_b_22')
// (11, 17, 'sp4_r_v_b_11')
// (12, 13, 'sp4_v_t_46')
// (12, 14, 'neigh_op_tnl_1')
// (12, 14, 'sp4_v_b_46')
// (12, 15, 'neigh_op_lft_1')
// (12, 15, 'sp4_v_b_35')
// (12, 16, 'neigh_op_bnl_1')
// (12, 16, 'sp4_v_b_22')
// (12, 17, 'local_g0_3')
// (12, 17, 'lutff_7/in_2')
// (12, 17, 'sp4_v_b_11')

wire n1489;
// (10, 14, 'neigh_op_tnr_2')
// (10, 15, 'neigh_op_rgt_2')
// (10, 16, 'neigh_op_bnr_2')
// (11, 14, 'neigh_op_top_2')
// (11, 15, 'lutff_2/out')
// (11, 16, 'neigh_op_bot_2')
// (12, 14, 'neigh_op_tnl_2')
// (12, 15, 'local_g1_2')
// (12, 15, 'lutff_6/in_1')
// (12, 15, 'neigh_op_lft_2')
// (12, 16, 'neigh_op_bnl_2')

reg n1490 = 0;
// (10, 14, 'neigh_op_tnr_3')
// (10, 15, 'neigh_op_rgt_3')
// (10, 15, 'sp4_r_v_b_38')
// (10, 16, 'neigh_op_bnr_3')
// (10, 16, 'sp4_r_v_b_27')
// (10, 17, 'sp4_r_v_b_14')
// (10, 18, 'sp4_r_v_b_3')
// (11, 14, 'neigh_op_top_3')
// (11, 14, 'sp4_v_t_38')
// (11, 15, 'lutff_3/out')
// (11, 15, 'sp4_v_b_38')
// (11, 16, 'neigh_op_bot_3')
// (11, 16, 'sp4_v_b_27')
// (11, 17, 'sp4_v_b_14')
// (11, 18, 'local_g1_3')
// (11, 18, 'lutff_5/in_3')
// (11, 18, 'sp4_v_b_3')
// (12, 14, 'neigh_op_tnl_3')
// (12, 15, 'neigh_op_lft_3')
// (12, 16, 'neigh_op_bnl_3')

reg n1491 = 0;
// (10, 14, 'neigh_op_tnr_4')
// (10, 15, 'neigh_op_rgt_4')
// (10, 15, 'sp4_r_v_b_40')
// (10, 16, 'neigh_op_bnr_4')
// (10, 16, 'sp4_r_v_b_29')
// (10, 17, 'sp4_r_v_b_16')
// (10, 18, 'sp4_r_v_b_5')
// (11, 14, 'neigh_op_top_4')
// (11, 14, 'sp4_r_v_b_36')
// (11, 14, 'sp4_v_t_40')
// (11, 15, 'local_g2_4')
// (11, 15, 'lutff_4/in_2')
// (11, 15, 'lutff_4/out')
// (11, 15, 'sp4_h_r_8')
// (11, 15, 'sp4_r_v_b_25')
// (11, 15, 'sp4_r_v_b_41')
// (11, 15, 'sp4_v_b_40')
// (11, 16, 'neigh_op_bot_4')
// (11, 16, 'sp4_r_v_b_12')
// (11, 16, 'sp4_r_v_b_28')
// (11, 16, 'sp4_v_b_29')
// (11, 17, 'sp4_r_v_b_1')
// (11, 17, 'sp4_r_v_b_17')
// (11, 17, 'sp4_v_b_16')
// (11, 18, 'sp4_h_r_11')
// (11, 18, 'sp4_r_v_b_4')
// (11, 18, 'sp4_r_v_b_44')
// (11, 18, 'sp4_v_b_5')
// (11, 19, 'sp4_r_v_b_33')
// (11, 19, 'sp4_r_v_b_42')
// (11, 20, 'sp4_r_v_b_20')
// (11, 20, 'sp4_r_v_b_31')
// (11, 21, 'sp4_r_v_b_18')
// (11, 21, 'sp4_r_v_b_9')
// (11, 22, 'sp4_r_v_b_7')
// (12, 13, 'sp4_v_t_36')
// (12, 14, 'neigh_op_tnl_4')
// (12, 14, 'sp4_v_b_36')
// (12, 14, 'sp4_v_t_41')
// (12, 15, 'local_g0_4')
// (12, 15, 'lutff_4/in_2')
// (12, 15, 'neigh_op_lft_4')
// (12, 15, 'sp4_h_r_21')
// (12, 15, 'sp4_v_b_25')
// (12, 15, 'sp4_v_b_41')
// (12, 16, 'neigh_op_bnl_4')
// (12, 16, 'sp4_v_b_12')
// (12, 16, 'sp4_v_b_28')
// (12, 17, 'sp4_h_r_7')
// (12, 17, 'sp4_v_b_1')
// (12, 17, 'sp4_v_b_17')
// (12, 17, 'sp4_v_t_44')
// (12, 18, 'sp4_h_r_22')
// (12, 18, 'sp4_v_b_4')
// (12, 18, 'sp4_v_b_44')
// (12, 18, 'sp4_v_t_42')
// (12, 19, 'sp4_v_b_33')
// (12, 19, 'sp4_v_b_42')
// (12, 20, 'sp4_v_b_20')
// (12, 20, 'sp4_v_b_31')
// (12, 21, 'sp4_h_r_3')
// (12, 21, 'sp4_v_b_18')
// (12, 21, 'sp4_v_b_9')
// (12, 22, 'sp4_h_r_1')
// (12, 22, 'sp4_v_b_7')
// (13, 15, 'sp4_h_r_32')
// (13, 17, 'sp4_h_r_18')
// (13, 18, 'sp4_h_r_35')
// (13, 21, 'local_g0_6')
// (13, 21, 'lutff_0/in_0')
// (13, 21, 'lutff_1/in_1')
// (13, 21, 'lutff_2/in_0')
// (13, 21, 'lutff_3/in_3')
// (13, 21, 'lutff_6/in_0')
// (13, 21, 'sp4_h_r_14')
// (13, 22, 'local_g0_4')
// (13, 22, 'lutff_1/in_1')
// (13, 22, 'lutff_3/in_3')
// (13, 22, 'sp4_h_r_12')
// (14, 15, 'sp4_h_r_45')
// (14, 16, 'sp4_r_v_b_36')
// (14, 17, 'sp4_h_r_31')
// (14, 17, 'sp4_r_v_b_25')
// (14, 18, 'sp4_h_r_46')
// (14, 18, 'sp4_r_v_b_12')
// (14, 19, 'sp4_r_v_b_1')
// (14, 19, 'sp4_r_v_b_46')
// (14, 20, 'sp4_r_v_b_35')
// (14, 21, 'local_g3_6')
// (14, 21, 'lutff_1/in_0')
// (14, 21, 'lutff_3/in_0')
// (14, 21, 'lutff_5/in_2')
// (14, 21, 'lutff_7/in_0')
// (14, 21, 'sp4_h_r_27')
// (14, 21, 'sp4_r_v_b_22')
// (14, 22, 'sp4_h_r_25')
// (14, 22, 'sp4_r_v_b_11')
// (15, 15, 'sp4_h_l_45')
// (15, 15, 'sp4_v_t_36')
// (15, 16, 'local_g3_4')
// (15, 16, 'lutff_6/in_3')
// (15, 16, 'sp4_v_b_36')
// (15, 17, 'sp4_h_r_42')
// (15, 17, 'sp4_v_b_25')
// (15, 18, 'sp4_h_l_46')
// (15, 18, 'sp4_r_v_b_37')
// (15, 18, 'sp4_v_b_12')
// (15, 18, 'sp4_v_t_46')
// (15, 19, 'sp4_r_v_b_24')
// (15, 19, 'sp4_v_b_1')
// (15, 19, 'sp4_v_b_46')
// (15, 20, 'local_g2_5')
// (15, 20, 'lutff_0/in_1')
// (15, 20, 'lutff_5/in_2')
// (15, 20, 'sp4_r_v_b_13')
// (15, 20, 'sp4_v_b_35')
// (15, 21, 'sp4_h_r_38')
// (15, 21, 'sp4_r_v_b_0')
// (15, 21, 'sp4_v_b_22')
// (15, 22, 'sp4_h_r_36')
// (15, 22, 'sp4_v_b_11')
// (16, 17, 'sp4_h_l_42')
// (16, 17, 'sp4_v_t_37')
// (16, 18, 'sp4_v_b_37')
// (16, 19, 'sp4_v_b_24')
// (16, 20, 'sp4_v_b_13')
// (16, 21, 'sp4_h_l_38')
// (16, 21, 'sp4_v_b_0')
// (16, 22, 'sp4_h_l_36')

wire n1492;
// (10, 14, 'neigh_op_tnr_5')
// (10, 15, 'neigh_op_rgt_5')
// (10, 16, 'neigh_op_bnr_5')
// (11, 14, 'neigh_op_top_5')
// (11, 15, 'lutff_5/out')
// (11, 16, 'neigh_op_bot_5')
// (12, 14, 'neigh_op_tnl_5')
// (12, 15, 'local_g0_5')
// (12, 15, 'lutff_7/in_0')
// (12, 15, 'neigh_op_lft_5')
// (12, 16, 'neigh_op_bnl_5')

wire n1493;
// (10, 14, 'neigh_op_tnr_7')
// (10, 15, 'neigh_op_rgt_7')
// (10, 16, 'neigh_op_bnr_7')
// (11, 14, 'neigh_op_top_7')
// (11, 15, 'lutff_7/out')
// (11, 16, 'neigh_op_bot_7')
// (12, 14, 'neigh_op_tnl_7')
// (12, 15, 'local_g0_7')
// (12, 15, 'lutff_6/in_3')
// (12, 15, 'neigh_op_lft_7')
// (12, 16, 'neigh_op_bnl_7')

wire n1494;
// (10, 14, 'sp4_h_r_1')
// (11, 14, 'sp4_h_r_12')
// (12, 12, 'sp4_r_v_b_44')
// (12, 13, 'neigh_op_tnr_2')
// (12, 13, 'sp4_r_v_b_33')
// (12, 14, 'neigh_op_rgt_2')
// (12, 14, 'sp4_h_r_25')
// (12, 14, 'sp4_r_v_b_20')
// (12, 15, 'neigh_op_bnr_2')
// (12, 15, 'sp4_r_v_b_9')
// (13, 11, 'sp4_v_t_44')
// (13, 12, 'local_g2_4')
// (13, 12, 'local_g3_4')
// (13, 12, 'lutff_0/in_1')
// (13, 12, 'lutff_3/in_2')
// (13, 12, 'lutff_4/in_2')
// (13, 12, 'sp4_v_b_44')
// (13, 13, 'neigh_op_top_2')
// (13, 13, 'sp4_v_b_33')
// (13, 14, 'local_g3_2')
// (13, 14, 'lutff_0/in_1')
// (13, 14, 'lutff_2/out')
// (13, 14, 'lutff_3/in_2')
// (13, 14, 'sp4_h_r_36')
// (13, 14, 'sp4_r_v_b_37')
// (13, 14, 'sp4_v_b_20')
// (13, 15, 'neigh_op_bot_2')
// (13, 15, 'sp4_r_v_b_24')
// (13, 15, 'sp4_v_b_9')
// (13, 16, 'sp4_r_v_b_13')
// (13, 17, 'sp4_r_v_b_0')
// (14, 13, 'local_g2_2')
// (14, 13, 'local_g3_2')
// (14, 13, 'lutff_1/in_0')
// (14, 13, 'lutff_5/in_1')
// (14, 13, 'lutff_6/in_2')
// (14, 13, 'neigh_op_tnl_2')
// (14, 13, 'sp4_h_r_5')
// (14, 13, 'sp4_v_t_37')
// (14, 14, 'local_g1_2')
// (14, 14, 'lutff_2/in_3')
// (14, 14, 'lutff_4/in_1')
// (14, 14, 'lutff_7/in_2')
// (14, 14, 'neigh_op_lft_2')
// (14, 14, 'sp4_h_l_36')
// (14, 14, 'sp4_h_r_9')
// (14, 14, 'sp4_v_b_37')
// (14, 15, 'neigh_op_bnl_2')
// (14, 15, 'sp4_v_b_24')
// (14, 16, 'sp4_v_b_13')
// (14, 17, 'sp4_v_b_0')
// (15, 13, 'local_g0_0')
// (15, 13, 'lutff_6/in_2')
// (15, 13, 'sp4_h_r_16')
// (15, 14, 'local_g0_4')
// (15, 14, 'lutff_0/in_2')
// (15, 14, 'lutff_7/in_1')
// (15, 14, 'sp4_h_r_20')
// (16, 13, 'sp4_h_r_29')
// (16, 14, 'sp4_h_r_33')
// (17, 13, 'sp4_h_r_40')
// (17, 14, 'sp4_h_r_44')
// (18, 13, 'sp4_h_l_40')
// (18, 14, 'sp4_h_l_44')

reg n1495 = 0;
// (10, 14, 'sp4_r_v_b_41')
// (10, 15, 'local_g1_4')
// (10, 15, 'lutff_1/in_2')
// (10, 15, 'sp4_r_v_b_28')
// (10, 16, 'sp4_r_v_b_17')
// (10, 17, 'sp4_r_v_b_4')
// (11, 13, 'sp4_v_t_41')
// (11, 14, 'sp4_v_b_41')
// (11, 15, 'sp4_v_b_28')
// (11, 16, 'neigh_op_tnr_3')
// (11, 16, 'sp4_v_b_17')
// (11, 17, 'neigh_op_rgt_3')
// (11, 17, 'sp4_h_r_11')
// (11, 17, 'sp4_v_b_4')
// (11, 18, 'neigh_op_bnr_3')
// (12, 16, 'neigh_op_top_3')
// (12, 17, 'local_g2_3')
// (12, 17, 'lutff_3/in_0')
// (12, 17, 'lutff_3/out')
// (12, 17, 'lutff_7/in_0')
// (12, 17, 'sp4_h_r_22')
// (12, 18, 'neigh_op_bot_3')
// (13, 16, 'neigh_op_tnl_3')
// (13, 17, 'neigh_op_lft_3')
// (13, 17, 'sp4_h_r_35')
// (13, 18, 'neigh_op_bnl_3')
// (14, 17, 'sp4_h_r_46')
// (15, 17, 'sp4_h_l_46')

reg n1496 = 0;
// (10, 15, 'neigh_op_tnr_0')
// (10, 16, 'neigh_op_rgt_0')
// (10, 17, 'neigh_op_bnr_0')
// (11, 15, 'local_g1_0')
// (11, 15, 'lutff_7/in_0')
// (11, 15, 'neigh_op_top_0')
// (11, 16, 'lutff_0/out')
// (11, 17, 'neigh_op_bot_0')
// (12, 15, 'neigh_op_tnl_0')
// (12, 16, 'neigh_op_lft_0')
// (12, 17, 'neigh_op_bnl_0')

wire n1497;
// (10, 15, 'neigh_op_tnr_1')
// (10, 16, 'neigh_op_rgt_1')
// (10, 17, 'neigh_op_bnr_1')
// (11, 15, 'neigh_op_top_1')
// (11, 16, 'local_g2_1')
// (11, 16, 'lutff_1/out')
// (11, 16, 'lutff_2/in_3')
// (11, 16, 'lutff_3/in_2')
// (11, 17, 'neigh_op_bot_1')
// (12, 15, 'neigh_op_tnl_1')
// (12, 16, 'neigh_op_lft_1')
// (12, 17, 'neigh_op_bnl_1')

reg n1498 = 0;
// (10, 15, 'neigh_op_tnr_2')
// (10, 16, 'neigh_op_rgt_2')
// (10, 17, 'neigh_op_bnr_2')
// (11, 15, 'local_g0_2')
// (11, 15, 'lutff_2/in_2')
// (11, 15, 'neigh_op_top_2')
// (11, 16, 'lutff_2/out')
// (11, 17, 'neigh_op_bot_2')
// (12, 15, 'neigh_op_tnl_2')
// (12, 16, 'neigh_op_lft_2')
// (12, 17, 'neigh_op_bnl_2')

reg n1499 = 0;
// (10, 15, 'neigh_op_tnr_4')
// (10, 16, 'neigh_op_rgt_4')
// (10, 17, 'neigh_op_bnr_4')
// (11, 15, 'local_g1_4')
// (11, 15, 'lutff_2/in_1')
// (11, 15, 'neigh_op_top_4')
// (11, 16, 'lutff_4/out')
// (11, 17, 'neigh_op_bot_4')
// (12, 15, 'neigh_op_tnl_4')
// (12, 16, 'neigh_op_lft_4')
// (12, 17, 'neigh_op_bnl_4')

wire n1500;
// (10, 15, 'neigh_op_tnr_5')
// (10, 16, 'neigh_op_rgt_5')
// (10, 17, 'neigh_op_bnr_5')
// (11, 15, 'local_g0_5')
// (11, 15, 'lutff_4/in_1')
// (11, 15, 'neigh_op_top_5')
// (11, 16, 'lutff_5/out')
// (11, 17, 'neigh_op_bot_5')
// (12, 15, 'neigh_op_tnl_5')
// (12, 16, 'neigh_op_lft_5')
// (12, 17, 'neigh_op_bnl_5')

wire n1501;
// (10, 15, 'neigh_op_tnr_6')
// (10, 16, 'neigh_op_rgt_6')
// (10, 17, 'neigh_op_bnr_6')
// (11, 10, 'sp12_v_t_23')
// (11, 11, 'sp12_v_b_23')
// (11, 12, 'sp12_v_b_20')
// (11, 13, 'sp12_v_b_19')
// (11, 14, 'sp12_v_b_16')
// (11, 14, 'sp4_r_v_b_37')
// (11, 15, 'neigh_op_top_6')
// (11, 15, 'sp12_v_b_15')
// (11, 15, 'sp4_r_v_b_24')
// (11, 16, 'lutff_6/out')
// (11, 16, 'sp12_v_b_12')
// (11, 16, 'sp4_r_v_b_13')
// (11, 17, 'neigh_op_bot_6')
// (11, 17, 'sp12_v_b_11')
// (11, 17, 'sp4_r_v_b_0')
// (11, 18, 'sp12_v_b_8')
// (11, 18, 'sp4_r_v_b_45')
// (11, 19, 'sp12_v_b_7')
// (11, 19, 'sp4_r_v_b_32')
// (11, 20, 'local_g2_4')
// (11, 20, 'lutff_4/in_0')
// (11, 20, 'lutff_6/in_0')
// (11, 20, 'sp12_v_b_4')
// (11, 20, 'sp4_r_v_b_21')
// (11, 21, 'sp12_v_b_3')
// (11, 21, 'sp4_r_v_b_8')
// (11, 22, 'sp12_v_b_0')
// (12, 13, 'sp4_v_t_37')
// (12, 14, 'sp4_v_b_37')
// (12, 15, 'neigh_op_tnl_6')
// (12, 15, 'sp4_v_b_24')
// (12, 16, 'neigh_op_lft_6')
// (12, 16, 'sp4_v_b_13')
// (12, 17, 'neigh_op_bnl_6')
// (12, 17, 'sp4_v_b_0')
// (12, 17, 'sp4_v_t_45')
// (12, 18, 'sp4_v_b_45')
// (12, 19, 'sp4_v_b_32')
// (12, 20, 'local_g0_5')
// (12, 20, 'lutff_1/in_0')
// (12, 20, 'sp4_v_b_21')
// (12, 21, 'local_g0_0')
// (12, 21, 'lutff_7/in_1')
// (12, 21, 'sp4_v_b_8')

wire n1502;
// (10, 15, 'neigh_op_tnr_7')
// (10, 15, 'sp4_r_v_b_43')
// (10, 16, 'neigh_op_rgt_7')
// (10, 16, 'sp4_r_v_b_30')
// (10, 17, 'local_g3_3')
// (10, 17, 'lutff_global/cen')
// (10, 17, 'neigh_op_bnr_7')
// (10, 17, 'sp4_r_v_b_19')
// (10, 18, 'sp4_r_v_b_6')
// (11, 11, 'sp12_v_t_22')
// (11, 12, 'sp12_v_b_22')
// (11, 13, 'sp12_v_b_21')
// (11, 14, 'sp12_v_b_18')
// (11, 14, 'sp4_v_t_43')
// (11, 15, 'neigh_op_top_7')
// (11, 15, 'sp12_v_b_17')
// (11, 15, 'sp4_v_b_43')
// (11, 16, 'lutff_7/out')
// (11, 16, 'sp12_v_b_14')
// (11, 16, 'sp4_v_b_30')
// (11, 17, 'neigh_op_bot_7')
// (11, 17, 'sp12_v_b_13')
// (11, 17, 'sp4_v_b_19')
// (11, 18, 'sp12_v_b_10')
// (11, 18, 'sp4_v_b_6')
// (11, 19, 'sp12_v_b_9')
// (11, 20, 'sp12_v_b_6')
// (11, 21, 'sp12_v_b_5')
// (11, 22, 'sp12_v_b_2')
// (11, 23, 'sp12_v_b_1')
// (11, 23, 'sp12_v_t_22')
// (11, 24, 'sp12_v_b_22')
// (11, 25, 'sp12_v_b_21')
// (11, 26, 'sp12_v_b_18')
// (11, 27, 'sp12_v_b_17')
// (11, 28, 'sp12_v_b_14')
// (11, 29, 'sp12_v_b_13')
// (11, 30, 'local_g3_2')
// (11, 30, 'lutff_0/in_3')
// (11, 30, 'sp12_v_b_10')
// (11, 31, 'span12_vert_9')
// (12, 15, 'neigh_op_tnl_7')
// (12, 16, 'neigh_op_lft_7')
// (12, 17, 'neigh_op_bnl_7')

reg n1503 = 0;
// (10, 15, 'sp4_h_r_10')
// (11, 15, 'sp4_h_r_23')
// (12, 15, 'sp4_h_r_34')
// (13, 15, 'local_g2_7')
// (13, 15, 'lutff_5/in_0')
// (13, 15, 'sp4_h_r_47')
// (13, 16, 'sp4_r_v_b_47')
// (13, 17, 'sp4_r_v_b_34')
// (13, 18, 'local_g2_5')
// (13, 18, 'lutff_0/in_1')
// (13, 18, 'neigh_op_tnr_5')
// (13, 18, 'sp4_r_v_b_23')
// (13, 19, 'neigh_op_rgt_5')
// (13, 19, 'sp4_r_v_b_10')
// (13, 20, 'neigh_op_bnr_5')
// (14, 15, 'sp4_h_l_47')
// (14, 15, 'sp4_v_t_47')
// (14, 16, 'sp4_v_b_47')
// (14, 17, 'sp4_v_b_34')
// (14, 18, 'neigh_op_top_5')
// (14, 18, 'sp4_v_b_23')
// (14, 19, 'local_g2_5')
// (14, 19, 'lutff_5/in_2')
// (14, 19, 'lutff_5/out')
// (14, 19, 'sp4_v_b_10')
// (14, 20, 'neigh_op_bot_5')
// (15, 18, 'neigh_op_tnl_5')
// (15, 19, 'neigh_op_lft_5')
// (15, 20, 'neigh_op_bnl_5')

reg n1504 = 0;
// (10, 15, 'sp4_r_v_b_39')
// (10, 16, 'sp4_r_v_b_26')
// (10, 17, 'neigh_op_tnr_1')
// (10, 17, 'sp4_r_v_b_15')
// (10, 18, 'neigh_op_rgt_1')
// (10, 18, 'sp4_r_v_b_2')
// (10, 19, 'neigh_op_bnr_1')
// (11, 14, 'sp4_v_t_39')
// (11, 15, 'local_g2_7')
// (11, 15, 'lutff_0/in_3')
// (11, 15, 'sp4_v_b_39')
// (11, 16, 'sp4_v_b_26')
// (11, 17, 'neigh_op_top_1')
// (11, 17, 'sp4_v_b_15')
// (11, 18, 'lutff_1/out')
// (11, 18, 'sp4_v_b_2')
// (11, 19, 'neigh_op_bot_1')
// (12, 17, 'neigh_op_tnl_1')
// (12, 18, 'neigh_op_lft_1')
// (12, 19, 'neigh_op_bnl_1')

wire n1505;
// (10, 16, 'neigh_op_tnr_2')
// (10, 17, 'neigh_op_rgt_2')
// (10, 18, 'neigh_op_bnr_2')
// (11, 16, 'neigh_op_top_2')
// (11, 17, 'lutff_2/out')
// (11, 17, 'sp4_h_r_4')
// (11, 18, 'neigh_op_bot_2')
// (12, 16, 'neigh_op_tnl_2')
// (12, 17, 'local_g0_1')
// (12, 17, 'lutff_4/in_1')
// (12, 17, 'neigh_op_lft_2')
// (12, 17, 'sp4_h_r_17')
// (12, 18, 'neigh_op_bnl_2')
// (13, 17, 'sp4_h_r_28')
// (14, 17, 'sp4_h_r_41')
// (15, 17, 'sp4_h_l_41')

wire n1506;
// (10, 16, 'neigh_op_tnr_6')
// (10, 17, 'neigh_op_rgt_6')
// (10, 18, 'neigh_op_bnr_6')
// (11, 16, 'neigh_op_top_6')
// (11, 17, 'lutff_6/out')
// (11, 18, 'neigh_op_bot_6')
// (12, 16, 'neigh_op_tnl_6')
// (12, 17, 'local_g1_6')
// (12, 17, 'lutff_1/in_0')
// (12, 17, 'neigh_op_lft_6')
// (12, 18, 'neigh_op_bnl_6')

wire n1507;
// (10, 16, 'neigh_op_tnr_7')
// (10, 17, 'neigh_op_rgt_7')
// (10, 18, 'neigh_op_bnr_7')
// (11, 16, 'neigh_op_top_7')
// (11, 17, 'lutff_7/out')
// (11, 18, 'neigh_op_bot_7')
// (12, 16, 'neigh_op_tnl_7')
// (12, 17, 'local_g1_7')
// (12, 17, 'lutff_3/in_1')
// (12, 17, 'neigh_op_lft_7')
// (12, 18, 'neigh_op_bnl_7')

reg n1508 = 0;
// (10, 16, 'sp4_r_v_b_45')
// (10, 17, 'sp4_r_v_b_32')
// (10, 18, 'neigh_op_tnr_4')
// (10, 18, 'sp4_r_v_b_21')
// (10, 19, 'neigh_op_rgt_4')
// (10, 19, 'sp4_r_v_b_8')
// (10, 20, 'neigh_op_bnr_4')
// (11, 15, 'sp4_v_t_45')
// (11, 16, 'local_g2_5')
// (11, 16, 'lutff_1/in_2')
// (11, 16, 'sp4_v_b_45')
// (11, 17, 'sp4_v_b_32')
// (11, 18, 'neigh_op_top_4')
// (11, 18, 'sp4_v_b_21')
// (11, 19, 'local_g0_4')
// (11, 19, 'lutff_4/in_0')
// (11, 19, 'lutff_4/out')
// (11, 19, 'sp4_v_b_8')
// (11, 20, 'neigh_op_bot_4')
// (12, 18, 'neigh_op_tnl_4')
// (12, 19, 'neigh_op_lft_4')
// (12, 20, 'neigh_op_bnl_4')

reg n1509 = 0;
// (10, 17, 'neigh_op_tnr_2')
// (10, 18, 'neigh_op_rgt_2')
// (10, 19, 'neigh_op_bnr_2')
// (11, 17, 'neigh_op_top_2')
// (11, 18, 'local_g0_2')
// (11, 18, 'lutff_2/out')
// (11, 18, 'lutff_3/in_1')
// (11, 19, 'neigh_op_bot_2')
// (12, 17, 'neigh_op_tnl_2')
// (12, 18, 'neigh_op_lft_2')
// (12, 19, 'neigh_op_bnl_2')

wire n1510;
// (10, 17, 'neigh_op_tnr_3')
// (10, 18, 'neigh_op_rgt_3')
// (10, 19, 'neigh_op_bnr_3')
// (11, 17, 'local_g1_3')
// (11, 17, 'lutff_7/in_1')
// (11, 17, 'neigh_op_top_3')
// (11, 18, 'lutff_3/out')
// (11, 19, 'local_g1_3')
// (11, 19, 'lutff_4/in_2')
// (11, 19, 'neigh_op_bot_3')
// (12, 17, 'neigh_op_tnl_3')
// (12, 18, 'neigh_op_lft_3')
// (12, 19, 'neigh_op_bnl_3')

wire n1511;
// (10, 17, 'neigh_op_tnr_5')
// (10, 18, 'neigh_op_rgt_5')
// (10, 19, 'neigh_op_bnr_5')
// (11, 17, 'neigh_op_top_5')
// (11, 18, 'lutff_5/out')
// (11, 18, 'sp4_r_v_b_43')
// (11, 19, 'local_g1_5')
// (11, 19, 'lutff_7/in_3')
// (11, 19, 'neigh_op_bot_5')
// (11, 19, 'sp4_r_v_b_30')
// (11, 20, 'sp4_r_v_b_19')
// (11, 21, 'local_g1_6')
// (11, 21, 'lutff_1/in_2')
// (11, 21, 'lutff_5/in_0')
// (11, 21, 'sp4_r_v_b_6')
// (12, 17, 'neigh_op_tnl_5')
// (12, 17, 'sp4_v_t_43')
// (12, 18, 'neigh_op_lft_5')
// (12, 18, 'sp4_v_b_43')
// (12, 19, 'neigh_op_bnl_5')
// (12, 19, 'sp4_v_b_30')
// (12, 20, 'sp4_v_b_19')
// (12, 21, 'sp4_v_b_6')

reg n1512 = 0;
// (10, 17, 'neigh_op_tnr_6')
// (10, 18, 'neigh_op_rgt_6')
// (10, 19, 'neigh_op_bnr_6')
// (11, 17, 'local_g0_6')
// (11, 17, 'lutff_2/in_2')
// (11, 17, 'neigh_op_top_6')
// (11, 18, 'lutff_6/out')
// (11, 19, 'neigh_op_bot_6')
// (12, 17, 'neigh_op_tnl_6')
// (12, 18, 'neigh_op_lft_6')
// (12, 19, 'neigh_op_bnl_6')

wire n1513;
// (10, 17, 'sp4_h_r_2')
// (11, 17, 'sp4_h_r_15')
// (12, 17, 'sp4_h_r_26')
// (13, 17, 'sp4_h_r_39')
// (13, 18, 'sp4_r_v_b_42')
// (13, 19, 'sp4_r_v_b_31')
// (13, 20, 'sp4_r_v_b_18')
// (13, 21, 'sp4_r_v_b_7')
// (14, 17, 'sp4_h_l_39')
// (14, 17, 'sp4_h_r_2')
// (14, 17, 'sp4_v_t_42')
// (14, 18, 'local_g2_2')
// (14, 18, 'lutff_global/cen')
// (14, 18, 'sp4_v_b_42')
// (14, 19, 'sp4_v_b_31')
// (14, 20, 'sp4_v_b_18')
// (14, 21, 'sp4_v_b_7')
// (15, 14, 'sp4_r_v_b_47')
// (15, 15, 'sp4_r_v_b_34')
// (15, 16, 'neigh_op_tnr_5')
// (15, 16, 'sp4_r_v_b_23')
// (15, 17, 'neigh_op_rgt_5')
// (15, 17, 'sp4_h_r_15')
// (15, 17, 'sp4_r_v_b_10')
// (15, 18, 'neigh_op_bnr_5')
// (15, 18, 'sp4_r_v_b_43')
// (15, 19, 'sp4_r_v_b_30')
// (15, 20, 'sp4_r_v_b_19')
// (15, 21, 'sp4_r_v_b_6')
// (16, 13, 'sp4_v_t_47')
// (16, 14, 'sp4_v_b_47')
// (16, 15, 'sp4_v_b_34')
// (16, 16, 'neigh_op_top_5')
// (16, 16, 'sp4_v_b_23')
// (16, 17, 'lutff_5/out')
// (16, 17, 'sp4_h_r_26')
// (16, 17, 'sp4_r_v_b_43')
// (16, 17, 'sp4_v_b_10')
// (16, 17, 'sp4_v_t_43')
// (16, 18, 'local_g3_3')
// (16, 18, 'lutff_global/cen')
// (16, 18, 'neigh_op_bot_5')
// (16, 18, 'sp4_r_v_b_30')
// (16, 18, 'sp4_v_b_43')
// (16, 19, 'local_g3_3')
// (16, 19, 'lutff_global/cen')
// (16, 19, 'sp4_r_v_b_19')
// (16, 19, 'sp4_v_b_30')
// (16, 20, 'sp4_r_v_b_6')
// (16, 20, 'sp4_v_b_19')
// (16, 21, 'sp4_v_b_6')
// (17, 16, 'neigh_op_tnl_5')
// (17, 16, 'sp4_v_t_43')
// (17, 17, 'neigh_op_lft_5')
// (17, 17, 'sp4_h_r_39')
// (17, 17, 'sp4_v_b_43')
// (17, 18, 'neigh_op_bnl_5')
// (17, 18, 'sp4_v_b_30')
// (17, 19, 'sp4_v_b_19')
// (17, 20, 'sp4_v_b_6')
// (18, 17, 'sp4_h_l_39')

reg n1514 = 0;
// (10, 17, 'sp4_r_v_b_38')
// (10, 18, 'neigh_op_tnr_7')
// (10, 18, 'sp4_r_v_b_27')
// (10, 19, 'neigh_op_rgt_7')
// (10, 19, 'sp4_r_v_b_14')
// (10, 20, 'neigh_op_bnr_7')
// (10, 20, 'sp4_r_v_b_3')
// (11, 16, 'local_g1_0')
// (11, 16, 'lutff_5/in_2')
// (11, 16, 'sp4_h_r_8')
// (11, 16, 'sp4_v_t_38')
// (11, 17, 'sp4_v_b_38')
// (11, 18, 'neigh_op_top_7')
// (11, 18, 'sp4_v_b_27')
// (11, 19, 'local_g2_7')
// (11, 19, 'lutff_7/in_2')
// (11, 19, 'lutff_7/out')
// (11, 19, 'sp4_v_b_14')
// (11, 20, 'neigh_op_bot_7')
// (11, 20, 'sp4_v_b_3')
// (12, 16, 'sp4_h_r_21')
// (12, 18, 'neigh_op_tnl_7')
// (12, 19, 'neigh_op_lft_7')
// (12, 20, 'neigh_op_bnl_7')
// (13, 16, 'sp4_h_r_32')
// (14, 16, 'sp4_h_r_45')
// (15, 16, 'sp4_h_l_45')

wire n1515;
// (10, 17, 'sp4_r_v_b_45')
// (10, 18, 'sp4_r_v_b_32')
// (10, 19, 'neigh_op_tnr_4')
// (10, 19, 'sp4_r_v_b_21')
// (10, 20, 'neigh_op_rgt_4')
// (10, 20, 'sp4_r_v_b_8')
// (10, 21, 'neigh_op_bnr_4')
// (11, 16, 'sp4_v_t_45')
// (11, 17, 'sp4_v_b_45')
// (11, 18, 'sp4_v_b_32')
// (11, 19, 'neigh_op_top_4')
// (11, 19, 'sp4_v_b_21')
// (11, 20, 'local_g0_2')
// (11, 20, 'lutff_4/out')
// (11, 20, 'lutff_global/cen')
// (11, 20, 'sp4_h_r_2')
// (11, 20, 'sp4_v_b_8')
// (11, 21, 'neigh_op_bot_4')
// (12, 19, 'neigh_op_tnl_4')
// (12, 20, 'neigh_op_lft_4')
// (12, 20, 'sp4_h_r_15')
// (12, 21, 'neigh_op_bnl_4')
// (13, 20, 'sp4_h_r_26')
// (14, 20, 'sp4_h_r_39')
// (15, 20, 'sp4_h_l_39')

wire n1516;
// (10, 18, 'lutff_7/cout')
// (10, 19, 'carry_in')
// (10, 19, 'carry_in_mux')
// (10, 19, 'lutff_0/in_3')

reg n1517 = 0;
// (10, 18, 'sp4_h_r_4')
// (11, 17, 'neigh_op_tnr_6')
// (11, 18, 'neigh_op_rgt_6')
// (11, 18, 'sp4_h_r_17')
// (11, 19, 'neigh_op_bnr_6')
// (12, 12, 'sp4_r_v_b_45')
// (12, 13, 'sp4_r_v_b_32')
// (12, 14, 'sp4_r_v_b_21')
// (12, 15, 'local_g2_0')
// (12, 15, 'lutff_3/in_3')
// (12, 15, 'sp4_r_v_b_8')
// (12, 16, 'sp4_r_v_b_37')
// (12, 17, 'neigh_op_top_6')
// (12, 17, 'sp4_r_v_b_24')
// (12, 18, 'lutff_6/out')
// (12, 18, 'sp4_h_r_28')
// (12, 18, 'sp4_r_v_b_13')
// (12, 18, 'sp4_r_v_b_45')
// (12, 19, 'neigh_op_bot_6')
// (12, 19, 'sp4_r_v_b_0')
// (12, 19, 'sp4_r_v_b_32')
// (12, 20, 'sp4_r_v_b_21')
// (12, 21, 'sp4_r_v_b_8')
// (13, 11, 'sp4_v_t_45')
// (13, 12, 'sp4_v_b_45')
// (13, 13, 'sp4_v_b_32')
// (13, 14, 'sp4_v_b_21')
// (13, 15, 'sp4_h_r_0')
// (13, 15, 'sp4_r_v_b_41')
// (13, 15, 'sp4_v_b_8')
// (13, 15, 'sp4_v_t_37')
// (13, 16, 'sp4_r_v_b_28')
// (13, 16, 'sp4_v_b_37')
// (13, 17, 'neigh_op_tnl_6')
// (13, 17, 'sp4_h_r_1')
// (13, 17, 'sp4_r_v_b_17')
// (13, 17, 'sp4_v_b_24')
// (13, 17, 'sp4_v_t_45')
// (13, 18, 'neigh_op_lft_6')
// (13, 18, 'sp4_h_r_41')
// (13, 18, 'sp4_r_v_b_4')
// (13, 18, 'sp4_v_b_13')
// (13, 18, 'sp4_v_b_45')
// (13, 19, 'neigh_op_bnl_6')
// (13, 19, 'sp4_v_b_0')
// (13, 19, 'sp4_v_b_32')
// (13, 20, 'sp4_v_b_21')
// (13, 21, 'sp4_v_b_8')
// (14, 14, 'sp4_v_t_41')
// (14, 15, 'local_g3_1')
// (14, 15, 'lutff_4/in_2')
// (14, 15, 'sp4_h_r_13')
// (14, 15, 'sp4_v_b_41')
// (14, 16, 'sp4_v_b_28')
// (14, 17, 'sp4_h_r_12')
// (14, 17, 'sp4_v_b_17')
// (14, 18, 'sp4_h_l_41')
// (14, 18, 'sp4_v_b_4')
// (15, 15, 'local_g2_0')
// (15, 15, 'lutff_7/in_1')
// (15, 15, 'sp4_h_r_24')
// (15, 17, 'sp4_h_r_25')
// (16, 15, 'sp4_h_r_37')
// (16, 17, 'local_g2_4')
// (16, 17, 'lutff_1/in_3')
// (16, 17, 'sp4_h_r_36')
// (17, 15, 'sp4_h_l_37')
// (17, 17, 'sp4_h_l_36')

wire n1518;
// (10, 18, 'sp4_h_r_7')
// (11, 18, 'local_g1_2')
// (11, 18, 'lutff_2/in_3')
// (11, 18, 'lutff_3/in_0')
// (11, 18, 'sp4_h_r_18')
// (12, 18, 'sp4_h_r_31')
// (13, 18, 'sp4_h_r_42')
// (14, 18, 'sp4_h_l_42')
// (14, 18, 'sp4_h_r_11')
// (15, 18, 'sp4_h_r_22')
// (16, 18, 'sp4_h_r_35')
// (17, 18, 'sp4_h_r_46')
// (18, 18, 'sp4_h_l_46')
// (18, 18, 'sp4_h_r_8')
// (19, 17, 'neigh_op_tnr_0')
// (19, 18, 'neigh_op_rgt_0')
// (19, 18, 'sp4_h_r_21')
// (19, 19, 'neigh_op_bnr_0')
// (20, 17, 'neigh_op_top_0')
// (20, 18, 'lutff_0/out')
// (20, 18, 'sp4_h_r_32')
// (20, 19, 'neigh_op_bot_0')
// (21, 17, 'neigh_op_tnl_0')
// (21, 18, 'neigh_op_lft_0')
// (21, 18, 'sp4_h_r_45')
// (21, 19, 'neigh_op_bnl_0')
// (22, 18, 'sp4_h_l_45')

wire n1519;
// (10, 19, 'neigh_op_tnr_1')
// (10, 20, 'neigh_op_rgt_1')
// (10, 21, 'local_g0_1')
// (10, 21, 'lutff_4/in_1')
// (10, 21, 'neigh_op_bnr_1')
// (11, 19, 'local_g1_1')
// (11, 19, 'lutff_5/in_1')
// (11, 19, 'neigh_op_top_1')
// (11, 20, 'lutff_1/out')
// (11, 21, 'local_g0_1')
// (11, 21, 'lutff_2/in_1')
// (11, 21, 'lutff_4/in_1')
// (11, 21, 'lutff_6/in_1')
// (11, 21, 'neigh_op_bot_1')
// (12, 19, 'neigh_op_tnl_1')
// (12, 20, 'neigh_op_lft_1')
// (12, 21, 'neigh_op_bnl_1')

reg n1520 = 0;
// (10, 19, 'neigh_op_tnr_3')
// (10, 20, 'neigh_op_rgt_3')
// (10, 21, 'neigh_op_bnr_3')
// (11, 19, 'local_g0_3')
// (11, 19, 'lutff_7/in_0')
// (11, 19, 'neigh_op_top_3')
// (11, 20, 'local_g2_3')
// (11, 20, 'local_g3_3')
// (11, 20, 'lutff_1/in_3')
// (11, 20, 'lutff_3/in_1')
// (11, 20, 'lutff_3/out')
// (11, 20, 'lutff_4/in_3')
// (11, 21, 'neigh_op_bot_3')
// (12, 19, 'neigh_op_tnl_3')
// (12, 20, 'neigh_op_lft_3')
// (12, 21, 'neigh_op_bnl_3')

reg n1521 = 0;
// (10, 20, 'neigh_op_tnr_1')
// (10, 21, 'neigh_op_rgt_1')
// (10, 22, 'neigh_op_bnr_1')
// (11, 20, 'neigh_op_top_1')
// (11, 21, 'local_g3_1')
// (11, 21, 'lutff_1/in_1')
// (11, 21, 'lutff_1/out')
// (11, 21, 'lutff_5/in_3')
// (11, 22, 'neigh_op_bot_1')
// (12, 20, 'neigh_op_tnl_1')
// (12, 21, 'neigh_op_lft_1')
// (12, 22, 'neigh_op_bnl_1')

wire n1522;
// (10, 20, 'neigh_op_tnr_2')
// (10, 21, 'neigh_op_rgt_2')
// (10, 22, 'neigh_op_bnr_2')
// (11, 20, 'neigh_op_top_2')
// (11, 21, 'local_g1_2')
// (11, 21, 'local_g2_2')
// (11, 21, 'lutff_1/in_0')
// (11, 21, 'lutff_2/out')
// (11, 21, 'lutff_3/in_1')
// (11, 22, 'neigh_op_bot_2')
// (12, 20, 'neigh_op_tnl_2')
// (12, 21, 'neigh_op_lft_2')
// (12, 22, 'neigh_op_bnl_2')

wire n1523;
// (10, 20, 'neigh_op_tnr_4')
// (10, 21, 'neigh_op_rgt_4')
// (10, 22, 'neigh_op_bnr_4')
// (11, 20, 'neigh_op_top_4')
// (11, 21, 'lutff_4/out')
// (11, 22, 'neigh_op_bot_4')
// (12, 20, 'neigh_op_tnl_4')
// (12, 21, 'local_g1_4')
// (12, 21, 'lutff_5/in_0')
// (12, 21, 'lutff_7/in_2')
// (12, 21, 'neigh_op_lft_4')
// (12, 22, 'neigh_op_bnl_4')

wire n1524;
// (10, 20, 'neigh_op_tnr_5')
// (10, 21, 'neigh_op_rgt_5')
// (10, 22, 'neigh_op_bnr_5')
// (11, 20, 'neigh_op_top_5')
// (11, 21, 'local_g0_5')
// (11, 21, 'lutff_3/in_0')
// (11, 21, 'lutff_5/out')
// (11, 22, 'neigh_op_bot_5')
// (12, 20, 'neigh_op_tnl_5')
// (12, 21, 'neigh_op_lft_5')
// (12, 22, 'neigh_op_bnl_5')

wire n1525;
// (10, 20, 'neigh_op_tnr_6')
// (10, 21, 'neigh_op_rgt_6')
// (10, 22, 'neigh_op_bnr_6')
// (11, 20, 'neigh_op_top_6')
// (11, 21, 'local_g0_6')
// (11, 21, 'lutff_4/in_0')
// (11, 21, 'lutff_5/in_1')
// (11, 21, 'lutff_6/out')
// (11, 22, 'neigh_op_bot_6')
// (12, 20, 'neigh_op_tnl_6')
// (12, 21, 'neigh_op_lft_6')
// (12, 22, 'neigh_op_bnl_6')

wire n1526;
// (10, 21, 'sp4_h_r_4')
// (11, 21, 'sp4_h_r_17')
// (12, 21, 'sp4_h_r_28')
// (13, 21, 'sp4_h_r_41')
// (14, 21, 'sp4_h_l_41')
// (14, 21, 'sp4_h_r_1')
// (14, 21, 'sp4_h_r_7')
// (15, 21, 'local_g0_2')
// (15, 21, 'lutff_global/cen')
// (15, 21, 'sp4_h_r_12')
// (15, 21, 'sp4_h_r_18')
// (16, 20, 'neigh_op_tnr_2')
// (16, 21, 'local_g2_2')
// (16, 21, 'lutff_1/in_3')
// (16, 21, 'neigh_op_rgt_2')
// (16, 21, 'sp4_h_r_25')
// (16, 21, 'sp4_h_r_31')
// (16, 22, 'neigh_op_bnr_2')
// (17, 20, 'neigh_op_top_2')
// (17, 21, 'lutff_2/out')
// (17, 21, 'sp4_h_r_36')
// (17, 21, 'sp4_h_r_42')
// (17, 22, 'neigh_op_bot_2')
// (18, 20, 'neigh_op_tnl_2')
// (18, 21, 'neigh_op_lft_2')
// (18, 21, 'sp4_h_l_36')
// (18, 21, 'sp4_h_l_42')
// (18, 22, 'neigh_op_bnl_2')

wire n1527;
// (10, 21, 'sp4_h_r_5')
// (11, 21, 'sp4_h_r_16')
// (12, 20, 'neigh_op_tnr_4')
// (12, 21, 'neigh_op_rgt_4')
// (12, 21, 'sp4_h_r_29')
// (12, 22, 'neigh_op_bnr_4')
// (13, 18, 'sp4_r_v_b_46')
// (13, 19, 'sp4_r_v_b_35')
// (13, 20, 'neigh_op_top_4')
// (13, 20, 'sp4_r_v_b_22')
// (13, 21, 'lutff_4/out')
// (13, 21, 'sp4_h_r_40')
// (13, 21, 'sp4_r_v_b_11')
// (13, 22, 'local_g1_4')
// (13, 22, 'lutff_1/in_0')
// (13, 22, 'neigh_op_bot_4')
// (14, 17, 'sp4_v_t_46')
// (14, 18, 'sp4_v_b_46')
// (14, 19, 'local_g3_3')
// (14, 19, 'lutff_global/cen')
// (14, 19, 'sp4_v_b_35')
// (14, 20, 'neigh_op_tnl_4')
// (14, 20, 'sp4_v_b_22')
// (14, 21, 'neigh_op_lft_4')
// (14, 21, 'sp4_h_l_40')
// (14, 21, 'sp4_v_b_11')
// (14, 22, 'neigh_op_bnl_4')

reg n1528 = 0;
// (10, 23, 'sp4_h_r_0')
// (11, 22, 'neigh_op_tnr_4')
// (11, 23, 'neigh_op_rgt_4')
// (11, 23, 'sp4_h_r_13')
// (11, 24, 'neigh_op_bnr_4')
// (12, 22, 'local_g1_4')
// (12, 22, 'lutff_1/in_2')
// (12, 22, 'neigh_op_top_4')
// (12, 23, 'lutff_4/out')
// (12, 23, 'sp4_h_r_24')
// (12, 23, 'sp4_h_r_8')
// (12, 24, 'neigh_op_bot_4')
// (13, 20, 'sp4_r_v_b_37')
// (13, 21, 'sp4_r_v_b_24')
// (13, 22, 'neigh_op_tnl_4')
// (13, 22, 'sp4_r_v_b_13')
// (13, 23, 'neigh_op_lft_4')
// (13, 23, 'sp4_h_r_21')
// (13, 23, 'sp4_h_r_37')
// (13, 23, 'sp4_r_v_b_0')
// (13, 24, 'neigh_op_bnl_4')
// (14, 19, 'sp4_v_t_37')
// (14, 20, 'sp4_v_b_37')
// (14, 21, 'sp4_v_b_24')
// (14, 22, 'local_g0_5')
// (14, 22, 'lutff_5/in_2')
// (14, 22, 'sp4_v_b_13')
// (14, 23, 'local_g2_0')
// (14, 23, 'lutff_1/in_1')
// (14, 23, 'sp4_h_l_37')
// (14, 23, 'sp4_h_r_32')
// (14, 23, 'sp4_v_b_0')
// (15, 23, 'sp4_h_r_45')
// (16, 23, 'sp4_h_l_45')

wire n1529;
// (11, 1, 'local_g1_4')
// (11, 1, 'lutff_7/in_2')
// (11, 1, 'sp4_r_v_b_4')
// (11, 3, 'sp4_h_r_3')
// (12, 0, 'span4_vert_4')
// (12, 1, 'local_g0_4')
// (12, 1, 'lutff_7/in_1')
// (12, 1, 'sp4_h_r_4')
// (12, 1, 'sp4_v_b_4')
// (12, 3, 'local_g0_6')
// (12, 3, 'lutff_6/in_2')
// (12, 3, 'sp4_h_r_14')
// (13, 1, 'local_g1_1')
// (13, 1, 'lutff_7/in_1')
// (13, 1, 'sp4_h_r_17')
// (13, 3, 'sp4_h_r_27')
// (14, 1, 'sp4_h_r_28')
// (14, 3, 'sp4_h_r_38')
// (15, 1, 'sp4_h_r_41')
// (15, 2, 'neigh_op_tnr_1')
// (15, 2, 'sp4_r_v_b_47')
// (15, 3, 'neigh_op_rgt_1')
// (15, 3, 'sp4_h_l_38')
// (15, 3, 'sp4_h_r_7')
// (15, 3, 'sp4_r_v_b_34')
// (15, 4, 'neigh_op_bnr_1')
// (15, 4, 'sp4_r_v_b_23')
// (15, 5, 'sp4_r_v_b_10')
// (16, 1, 'sp4_h_l_41')
// (16, 1, 'sp4_v_t_47')
// (16, 2, 'neigh_op_top_1')
// (16, 2, 'sp4_v_b_47')
// (16, 3, 'lutff_1/out')
// (16, 3, 'sp4_h_r_18')
// (16, 3, 'sp4_v_b_34')
// (16, 4, 'neigh_op_bot_1')
// (16, 4, 'sp4_v_b_23')
// (16, 5, 'sp4_v_b_10')
// (17, 2, 'neigh_op_tnl_1')
// (17, 3, 'neigh_op_lft_1')
// (17, 3, 'sp4_h_r_31')
// (17, 4, 'neigh_op_bnl_1')
// (18, 3, 'sp4_h_r_42')
// (19, 3, 'sp4_h_l_42')

wire n1530;
// (11, 1, 'local_g2_2')
// (11, 1, 'lutff_4/in_2')
// (11, 1, 'neigh_op_tnr_2')
// (11, 2, 'neigh_op_rgt_2')
// (11, 3, 'neigh_op_bnr_2')
// (12, 1, 'local_g1_2')
// (12, 1, 'lutff_4/in_1')
// (12, 1, 'neigh_op_top_2')
// (12, 2, 'lutff_2/out')
// (12, 3, 'local_g1_2')
// (12, 3, 'lutff_3/in_2')
// (12, 3, 'neigh_op_bot_2')
// (13, 1, 'local_g2_2')
// (13, 1, 'lutff_4/in_2')
// (13, 1, 'neigh_op_tnl_2')
// (13, 2, 'neigh_op_lft_2')
// (13, 3, 'neigh_op_bnl_2')

wire n1531;
// (11, 1, 'local_g2_4')
// (11, 1, 'lutff_0/in_2')
// (11, 1, 'neigh_op_tnr_4')
// (11, 2, 'neigh_op_rgt_4')
// (11, 3, 'neigh_op_bnr_4')
// (12, 1, 'local_g1_4')
// (12, 1, 'lutff_0/in_1')
// (12, 1, 'neigh_op_top_4')
// (12, 2, 'lutff_4/out')
// (12, 3, 'neigh_op_bot_4')
// (13, 1, 'local_g2_4')
// (13, 1, 'lutff_0/in_2')
// (13, 1, 'neigh_op_tnl_4')
// (13, 2, 'neigh_op_lft_4')
// (13, 3, 'neigh_op_bnl_4')

wire n1532;
// (11, 1, 'local_g2_5')
// (11, 1, 'lutff_5/in_2')
// (11, 1, 'sp4_r_v_b_13')
// (11, 2, 'sp4_r_v_b_0')
// (12, 0, 'span4_vert_13')
// (12, 1, 'local_g3_1')
// (12, 1, 'lutff_5/in_1')
// (12, 1, 'neigh_op_tnr_1')
// (12, 1, 'sp4_v_b_13')
// (12, 2, 'neigh_op_rgt_1')
// (12, 2, 'sp4_h_r_7')
// (12, 2, 'sp4_v_b_0')
// (12, 3, 'local_g1_1')
// (12, 3, 'lutff_4/in_2')
// (12, 3, 'neigh_op_bnr_1')
// (13, 1, 'local_g0_1')
// (13, 1, 'lutff_5/in_2')
// (13, 1, 'neigh_op_top_1')
// (13, 2, 'lutff_1/out')
// (13, 2, 'sp4_h_r_18')
// (13, 3, 'neigh_op_bot_1')
// (14, 1, 'neigh_op_tnl_1')
// (14, 2, 'neigh_op_lft_1')
// (14, 2, 'sp4_h_r_31')
// (14, 3, 'neigh_op_bnl_1')
// (15, 2, 'sp4_h_r_42')
// (16, 2, 'sp4_h_l_42')

wire n1533;
// (11, 1, 'local_g2_6')
// (11, 1, 'lutff_2/in_2')
// (11, 1, 'neigh_op_tnr_6')
// (11, 2, 'neigh_op_rgt_6')
// (11, 3, 'neigh_op_bnr_6')
// (12, 1, 'local_g1_6')
// (12, 1, 'lutff_2/in_1')
// (12, 1, 'neigh_op_top_6')
// (12, 2, 'lutff_6/out')
// (12, 3, 'local_g1_6')
// (12, 3, 'lutff_1/in_2')
// (12, 3, 'neigh_op_bot_6')
// (13, 1, 'local_g2_6')
// (13, 1, 'lutff_2/in_2')
// (13, 1, 'neigh_op_tnl_6')
// (13, 2, 'neigh_op_lft_6')
// (13, 3, 'neigh_op_bnl_6')

wire n1534;
// (11, 1, 'local_g3_6')
// (11, 1, 'lutff_6/in_1')
// (11, 1, 'sp4_r_v_b_46')
// (11, 2, 'sp4_r_v_b_35')
// (11, 3, 'sp4_r_v_b_22')
// (11, 4, 'sp4_r_v_b_11')
// (12, 0, 'span4_vert_46')
// (12, 1, 'local_g0_3')
// (12, 1, 'lutff_6/in_1')
// (12, 1, 'sp4_r_v_b_32')
// (12, 1, 'sp4_v_b_46')
// (12, 2, 'sp4_r_v_b_21')
// (12, 2, 'sp4_v_b_35')
// (12, 3, 'local_g2_0')
// (12, 3, 'lutff_5/in_1')
// (12, 3, 'sp4_r_v_b_8')
// (12, 3, 'sp4_v_b_22')
// (12, 4, 'sp4_h_r_11')
// (12, 4, 'sp4_v_b_11')
// (13, 0, 'span4_vert_32')
// (13, 1, 'local_g3_0')
// (13, 1, 'lutff_6/in_1')
// (13, 1, 'sp4_v_b_32')
// (13, 2, 'sp4_v_b_21')
// (13, 3, 'sp4_h_r_3')
// (13, 3, 'sp4_v_b_8')
// (13, 4, 'sp4_h_r_22')
// (14, 3, 'sp4_h_r_14')
// (14, 4, 'sp4_h_r_35')
// (15, 1, 'sp4_r_v_b_46')
// (15, 2, 'neigh_op_tnr_3')
// (15, 2, 'sp4_r_v_b_35')
// (15, 3, 'neigh_op_rgt_3')
// (15, 3, 'sp4_h_r_27')
// (15, 3, 'sp4_r_v_b_22')
// (15, 4, 'neigh_op_bnr_3')
// (15, 4, 'sp4_h_r_46')
// (15, 4, 'sp4_r_v_b_11')
// (16, 0, 'span4_vert_46')
// (16, 1, 'sp4_v_b_46')
// (16, 2, 'neigh_op_top_3')
// (16, 2, 'sp4_v_b_35')
// (16, 3, 'lutff_3/out')
// (16, 3, 'sp4_h_r_38')
// (16, 3, 'sp4_v_b_22')
// (16, 4, 'neigh_op_bot_3')
// (16, 4, 'sp4_h_l_46')
// (16, 4, 'sp4_v_b_11')
// (17, 2, 'neigh_op_tnl_3')
// (17, 3, 'neigh_op_lft_3')
// (17, 3, 'sp4_h_l_38')
// (17, 4, 'neigh_op_bnl_3')

wire n1535;
// (11, 1, 'local_g3_7')
// (11, 1, 'lutff_3/in_1')
// (11, 1, 'neigh_op_tnr_7')
// (11, 2, 'neigh_op_rgt_7')
// (11, 3, 'neigh_op_bnr_7')
// (12, 1, 'local_g0_7')
// (12, 1, 'lutff_3/in_2')
// (12, 1, 'neigh_op_top_7')
// (12, 2, 'lutff_7/out')
// (12, 3, 'local_g0_7')
// (12, 3, 'lutff_2/in_1')
// (12, 3, 'neigh_op_bot_7')
// (13, 1, 'local_g2_7')
// (13, 1, 'lutff_3/in_2')
// (13, 1, 'neigh_op_tnl_7')
// (13, 2, 'neigh_op_lft_7')
// (13, 3, 'neigh_op_bnl_7')

wire n1536;
// (11, 1, 'lutff_7/cout')
// (11, 2, 'carry_in')
// (11, 2, 'carry_in_mux')
// (11, 2, 'lutff_0/in_3')

wire n1537;
// (11, 1, 'neigh_op_tnr_0')
// (11, 2, 'neigh_op_rgt_0')
// (11, 3, 'neigh_op_bnr_0')
// (12, 1, 'neigh_op_top_0')
// (12, 2, 'local_g1_0')
// (12, 2, 'lutff_0/out')
// (12, 2, 'lutff_3/in_2')
// (12, 3, 'neigh_op_bot_0')
// (13, 1, 'neigh_op_tnl_0')
// (13, 2, 'neigh_op_lft_0')
// (13, 3, 'neigh_op_bnl_0')

wire n1538;
// (11, 1, 'neigh_op_tnr_3')
// (11, 2, 'neigh_op_rgt_3')
// (11, 2, 'sp4_r_v_b_38')
// (11, 3, 'neigh_op_bnr_3')
// (11, 3, 'sp4_r_v_b_27')
// (11, 4, 'sp4_r_v_b_14')
// (11, 5, 'sp4_r_v_b_3')
// (12, 1, 'neigh_op_top_3')
// (12, 1, 'sp4_v_t_38')
// (12, 2, 'lutff_3/out')
// (12, 2, 'sp4_v_b_38')
// (12, 3, 'neigh_op_bot_3')
// (12, 3, 'sp4_v_b_27')
// (12, 4, 'local_g0_6')
// (12, 4, 'lutff_6/in_2')
// (12, 4, 'sp4_v_b_14')
// (12, 5, 'sp4_v_b_3')
// (13, 1, 'neigh_op_tnl_3')
// (13, 2, 'neigh_op_lft_3')
// (13, 3, 'neigh_op_bnl_3')

wire n1539;
// (11, 1, 'sp4_r_v_b_41')
// (11, 2, 'local_g1_4')
// (11, 2, 'lutff_0/in_1')
// (11, 2, 'sp4_r_v_b_28')
// (11, 3, 'neigh_op_tnr_2')
// (11, 3, 'sp4_r_v_b_17')
// (11, 4, 'local_g2_2')
// (11, 4, 'lutff_7/in_1')
// (11, 4, 'neigh_op_rgt_2')
// (11, 4, 'sp4_r_v_b_4')
// (11, 5, 'local_g0_2')
// (11, 5, 'lutff_0/in_0')
// (11, 5, 'lutff_4/in_2')
// (11, 5, 'lutff_5/in_3')
// (11, 5, 'neigh_op_bnr_2')
// (12, 0, 'span4_vert_41')
// (12, 1, 'sp4_v_b_41')
// (12, 2, 'local_g2_4')
// (12, 2, 'lutff_3/in_3')
// (12, 2, 'sp4_v_b_28')
// (12, 3, 'local_g0_2')
// (12, 3, 'lutff_7/in_1')
// (12, 3, 'neigh_op_top_2')
// (12, 3, 'sp4_v_b_17')
// (12, 4, 'local_g3_2')
// (12, 4, 'lutff_2/out')
// (12, 4, 'lutff_3/in_0')
// (12, 4, 'sp4_v_b_4')
// (12, 5, 'neigh_op_bot_2')
// (13, 3, 'neigh_op_tnl_2')
// (13, 4, 'neigh_op_lft_2')
// (13, 5, 'neigh_op_bnl_2')

wire n1540;
// (11, 2, 'neigh_op_tnr_7')
// (11, 3, 'neigh_op_rgt_7')
// (11, 4, 'neigh_op_bnr_7')
// (12, 2, 'neigh_op_top_7')
// (12, 3, 'lutff_7/out')
// (12, 4, 'local_g1_7')
// (12, 4, 'lutff_3/in_3')
// (12, 4, 'neigh_op_bot_7')
// (13, 2, 'neigh_op_tnl_7')
// (13, 3, 'neigh_op_lft_7')
// (13, 4, 'neigh_op_bnl_7')

reg n1541 = 0;
// (11, 2, 'sp4_h_r_4')
// (11, 3, 'sp4_r_v_b_37')
// (11, 3, 'sp4_r_v_b_42')
// (11, 4, 'local_g1_0')
// (11, 4, 'lutff_3/in_2')
// (11, 4, 'sp4_r_v_b_24')
// (11, 4, 'sp4_r_v_b_31')
// (11, 5, 'local_g3_2')
// (11, 5, 'lutff_1/in_0')
// (11, 5, 'lutff_4/in_3')
// (11, 5, 'sp4_r_v_b_13')
// (11, 5, 'sp4_r_v_b_18')
// (11, 6, 'local_g1_0')
// (11, 6, 'lutff_2/in_1')
// (11, 6, 'sp4_r_v_b_0')
// (11, 6, 'sp4_r_v_b_7')
// (12, 2, 'local_g1_1')
// (12, 2, 'lutff_4/in_2')
// (12, 2, 'sp4_h_r_17')
// (12, 2, 'sp4_v_t_37')
// (12, 2, 'sp4_v_t_42')
// (12, 3, 'sp4_v_b_37')
// (12, 3, 'sp4_v_b_42')
// (12, 4, 'local_g2_0')
// (12, 4, 'lutff_7/in_3')
// (12, 4, 'sp4_v_b_24')
// (12, 4, 'sp4_v_b_31')
// (12, 5, 'sp4_v_b_13')
// (12, 5, 'sp4_v_b_18')
// (12, 6, 'sp4_h_r_7')
// (12, 6, 'sp4_v_b_0')
// (12, 6, 'sp4_v_b_7')
// (13, 2, 'sp4_h_r_28')
// (13, 6, 'sp4_h_r_18')
// (14, 2, 'sp4_h_r_41')
// (14, 3, 'sp4_r_v_b_47')
// (14, 4, 'sp4_r_v_b_34')
// (14, 5, 'local_g2_5')
// (14, 5, 'lutff_2/in_3')
// (14, 5, 'lutff_5/in_0')
// (14, 5, 'neigh_op_tnr_5')
// (14, 5, 'sp4_r_v_b_23')
// (14, 6, 'neigh_op_rgt_5')
// (14, 6, 'sp4_h_r_31')
// (14, 6, 'sp4_r_v_b_10')
// (14, 6, 'sp4_r_v_b_42')
// (14, 7, 'neigh_op_bnr_5')
// (14, 7, 'sp4_r_v_b_31')
// (14, 8, 'sp4_r_v_b_18')
// (14, 9, 'sp4_r_v_b_7')
// (14, 10, 'sp4_r_v_b_42')
// (14, 11, 'sp4_r_v_b_31')
// (14, 12, 'sp4_r_v_b_18')
// (14, 13, 'sp4_r_v_b_7')
// (14, 14, 'sp4_r_v_b_42')
// (14, 15, 'local_g1_7')
// (14, 15, 'lutff_0/in_0')
// (14, 15, 'lutff_1/in_3')
// (14, 15, 'sp4_r_v_b_31')
// (14, 16, 'sp4_r_v_b_18')
// (14, 17, 'sp4_r_v_b_7')
// (15, 2, 'sp4_h_l_41')
// (15, 2, 'sp4_v_t_47')
// (15, 3, 'local_g2_7')
// (15, 3, 'lutff_3/in_2')
// (15, 3, 'sp4_v_b_47')
// (15, 4, 'sp4_v_b_34')
// (15, 5, 'local_g1_5')
// (15, 5, 'lutff_5/in_3')
// (15, 5, 'lutff_7/in_3')
// (15, 5, 'neigh_op_top_5')
// (15, 5, 'sp4_v_b_23')
// (15, 5, 'sp4_v_t_42')
// (15, 6, 'local_g2_5')
// (15, 6, 'lutff_5/in_2')
// (15, 6, 'lutff_5/out')
// (15, 6, 'sp4_h_r_42')
// (15, 6, 'sp4_v_b_10')
// (15, 6, 'sp4_v_b_42')
// (15, 7, 'neigh_op_bot_5')
// (15, 7, 'sp4_v_b_31')
// (15, 8, 'sp4_v_b_18')
// (15, 9, 'sp4_v_b_7')
// (15, 9, 'sp4_v_t_42')
// (15, 10, 'sp4_v_b_42')
// (15, 11, 'sp4_v_b_31')
// (15, 12, 'sp4_v_b_18')
// (15, 13, 'sp4_v_b_7')
// (15, 13, 'sp4_v_t_42')
// (15, 14, 'sp4_v_b_42')
// (15, 15, 'sp4_v_b_31')
// (15, 16, 'sp4_v_b_18')
// (15, 17, 'sp4_v_b_7')
// (16, 5, 'neigh_op_tnl_5')
// (16, 6, 'neigh_op_lft_5')
// (16, 6, 'sp4_h_l_42')
// (16, 6, 'sp4_h_r_7')
// (16, 7, 'neigh_op_bnl_5')
// (17, 6, 'local_g0_2')
// (17, 6, 'lutff_0/in_2')
// (17, 6, 'sp4_h_r_18')
// (18, 6, 'sp4_h_r_31')
// (19, 6, 'sp4_h_r_42')
// (20, 6, 'sp4_h_l_42')

reg n1542 = 0;
// (11, 2, 'sp4_r_v_b_40')
// (11, 3, 'sp4_r_v_b_29')
// (11, 4, 'sp4_r_v_b_16')
// (11, 5, 'sp4_r_v_b_5')
// (12, 1, 'sp4_v_t_40')
// (12, 2, 'sp4_v_b_40')
// (12, 3, 'sp4_v_b_29')
// (12, 4, 'local_g1_0')
// (12, 4, 'lutff_4/in_1')
// (12, 4, 'sp4_v_b_16')
// (12, 5, 'sp4_h_r_5')
// (12, 5, 'sp4_v_b_5')
// (13, 5, 'sp4_h_r_16')
// (14, 4, 'neigh_op_tnr_4')
// (14, 5, 'neigh_op_rgt_4')
// (14, 5, 'sp4_h_r_29')
// (14, 6, 'local_g1_4')
// (14, 6, 'lutff_3/in_0')
// (14, 6, 'neigh_op_bnr_4')
// (15, 4, 'neigh_op_top_4')
// (15, 4, 'sp4_r_v_b_36')
// (15, 5, 'lutff_4/out')
// (15, 5, 'sp4_h_r_40')
// (15, 5, 'sp4_r_v_b_25')
// (15, 6, 'neigh_op_bot_4')
// (15, 6, 'sp4_r_v_b_12')
// (15, 7, 'sp4_r_v_b_1')
// (16, 3, 'sp4_v_t_36')
// (16, 4, 'neigh_op_tnl_4')
// (16, 4, 'sp4_v_b_36')
// (16, 5, 'local_g1_4')
// (16, 5, 'lutff_6/in_1')
// (16, 5, 'neigh_op_lft_4')
// (16, 5, 'sp4_h_l_40')
// (16, 5, 'sp4_v_b_25')
// (16, 6, 'local_g2_4')
// (16, 6, 'lutff_0/in_0')
// (16, 6, 'neigh_op_bnl_4')
// (16, 6, 'sp4_v_b_12')
// (16, 7, 'local_g1_1')
// (16, 7, 'lutff_5/in_3')
// (16, 7, 'sp4_v_b_1')

wire n1543;
// (11, 3, 'neigh_op_tnr_1')
// (11, 4, 'neigh_op_rgt_1')
// (11, 4, 'sp4_h_r_7')
// (11, 5, 'neigh_op_bnr_1')
// (12, 3, 'neigh_op_top_1')
// (12, 3, 'sp4_r_v_b_46')
// (12, 4, 'lutff_1/out')
// (12, 4, 'sp4_h_r_18')
// (12, 4, 'sp4_r_v_b_35')
// (12, 5, 'neigh_op_bot_1')
// (12, 5, 'sp4_r_v_b_22')
// (12, 6, 'sp4_r_v_b_11')
// (13, 2, 'sp4_h_r_4')
// (13, 2, 'sp4_v_t_46')
// (13, 3, 'local_g2_1')
// (13, 3, 'local_g3_1')
// (13, 3, 'lutff_0/in_3')
// (13, 3, 'lutff_4/in_2')
// (13, 3, 'lutff_5/in_2')
// (13, 3, 'neigh_op_tnl_1')
// (13, 3, 'sp4_v_b_46')
// (13, 4, 'local_g1_1')
// (13, 4, 'lutff_0/in_2')
// (13, 4, 'neigh_op_lft_1')
// (13, 4, 'sp4_h_r_31')
// (13, 4, 'sp4_v_b_35')
// (13, 5, 'neigh_op_bnl_1')
// (13, 5, 'sp4_v_b_22')
// (13, 6, 'sp4_v_b_11')
// (14, 1, 'sp4_r_v_b_36')
// (14, 1, 'sp4_r_v_b_42')
// (14, 2, 'sp4_h_r_17')
// (14, 2, 'sp4_r_v_b_25')
// (14, 2, 'sp4_r_v_b_31')
// (14, 3, 'local_g2_4')
// (14, 3, 'lutff_0/in_0')
// (14, 3, 'sp4_r_v_b_12')
// (14, 3, 'sp4_r_v_b_18')
// (14, 4, 'local_g2_2')
// (14, 4, 'lutff_7/in_3')
// (14, 4, 'sp4_h_r_42')
// (14, 4, 'sp4_r_v_b_1')
// (14, 4, 'sp4_r_v_b_7')
// (15, 0, 'span4_vert_36')
// (15, 0, 'span4_vert_42')
// (15, 1, 'sp4_v_b_36')
// (15, 1, 'sp4_v_b_42')
// (15, 2, 'local_g3_4')
// (15, 2, 'lutff_3/in_2')
// (15, 2, 'lutff_6/in_1')
// (15, 2, 'sp4_h_r_28')
// (15, 2, 'sp4_v_b_25')
// (15, 2, 'sp4_v_b_31')
// (15, 3, 'local_g1_2')
// (15, 3, 'lutff_5/in_2')
// (15, 3, 'sp4_v_b_12')
// (15, 3, 'sp4_v_b_18')
// (15, 4, 'local_g0_3')
// (15, 4, 'lutff_5/in_0')
// (15, 4, 'sp4_h_l_42')
// (15, 4, 'sp4_h_r_3')
// (15, 4, 'sp4_v_b_1')
// (15, 4, 'sp4_v_b_7')
// (16, 2, 'sp4_h_r_41')
// (16, 4, 'sp4_h_r_14')
// (17, 2, 'sp4_h_l_41')
// (17, 4, 'sp4_h_r_27')
// (18, 4, 'sp4_h_r_38')
// (19, 4, 'sp4_h_l_38')

wire n1544;
// (11, 3, 'neigh_op_tnr_3')
// (11, 4, 'neigh_op_rgt_3')
// (11, 5, 'neigh_op_bnr_3')
// (12, 3, 'neigh_op_top_3')
// (12, 4, 'local_g1_3')
// (12, 4, 'lutff_3/out')
// (12, 4, 'lutff_6/in_0')
// (12, 5, 'neigh_op_bot_3')
// (13, 3, 'neigh_op_tnl_3')
// (13, 4, 'neigh_op_lft_3')
// (13, 5, 'neigh_op_bnl_3')

wire n1545;
// (11, 3, 'neigh_op_tnr_4')
// (11, 4, 'neigh_op_rgt_4')
// (11, 5, 'neigh_op_bnr_4')
// (12, 3, 'neigh_op_top_4')
// (12, 4, 'lutff_4/out')
// (12, 5, 'local_g1_4')
// (12, 5, 'lutff_2/in_3')
// (12, 5, 'neigh_op_bot_4')
// (13, 3, 'neigh_op_tnl_4')
// (13, 4, 'neigh_op_lft_4')
// (13, 5, 'neigh_op_bnl_4')

wire n1546;
// (11, 3, 'neigh_op_tnr_5')
// (11, 4, 'neigh_op_rgt_5')
// (11, 5, 'neigh_op_bnr_5')
// (12, 3, 'neigh_op_top_5')
// (12, 4, 'local_g1_5')
// (12, 4, 'lutff_4/in_0')
// (12, 4, 'lutff_5/out')
// (12, 5, 'neigh_op_bot_5')
// (13, 3, 'neigh_op_tnl_5')
// (13, 4, 'neigh_op_lft_5')
// (13, 5, 'neigh_op_bnl_5')

wire n1547;
// (11, 3, 'sp4_h_r_6')
// (12, 3, 'sp4_h_r_19')
// (13, 3, 'sp4_h_r_30')
// (14, 2, 'neigh_op_tnr_5')
// (14, 3, 'neigh_op_rgt_5')
// (14, 3, 'sp4_h_r_43')
// (14, 4, 'neigh_op_bnr_5')
// (14, 4, 'sp4_r_v_b_43')
// (14, 5, 'sp4_r_v_b_30')
// (14, 6, 'sp4_r_v_b_19')
// (14, 7, 'sp4_r_v_b_6')
// (15, 2, 'neigh_op_top_5')
// (15, 3, 'local_g0_2')
// (15, 3, 'lutff_5/out')
// (15, 3, 'lutff_global/cen')
// (15, 3, 'sp4_h_l_43')
// (15, 3, 'sp4_h_r_10')
// (15, 3, 'sp4_v_t_43')
// (15, 4, 'local_g3_3')
// (15, 4, 'lutff_global/cen')
// (15, 4, 'neigh_op_bot_5')
// (15, 4, 'sp4_v_b_43')
// (15, 5, 'sp4_v_b_30')
// (15, 6, 'sp4_v_b_19')
// (15, 7, 'sp4_v_b_6')
// (16, 2, 'neigh_op_tnl_5')
// (16, 3, 'neigh_op_lft_5')
// (16, 3, 'sp4_h_r_23')
// (16, 4, 'neigh_op_bnl_5')
// (17, 3, 'sp4_h_r_34')
// (18, 3, 'sp4_h_r_47')
// (19, 3, 'sp4_h_l_47')

reg n1548 = 0;
// (11, 3, 'sp4_r_v_b_45')
// (11, 4, 'sp4_r_v_b_32')
// (11, 5, 'sp4_r_v_b_21')
// (11, 6, 'sp4_r_v_b_8')
// (11, 7, 'sp4_r_v_b_37')
// (11, 8, 'sp4_r_v_b_24')
// (11, 9, 'local_g2_0')
// (11, 9, 'lutff_1/in_1')
// (11, 9, 'neigh_op_tnr_0')
// (11, 9, 'sp4_r_v_b_13')
// (11, 10, 'neigh_op_rgt_0')
// (11, 10, 'sp4_r_v_b_0')
// (11, 11, 'neigh_op_bnr_0')
// (12, 0, 'span12_vert_19')
// (12, 1, 'sp12_v_b_19')
// (12, 2, 'sp12_v_b_16')
// (12, 2, 'sp4_v_t_45')
// (12, 3, 'sp12_v_b_15')
// (12, 3, 'sp4_v_b_45')
// (12, 4, 'sp12_v_b_12')
// (12, 4, 'sp4_v_b_32')
// (12, 5, 'local_g1_5')
// (12, 5, 'lutff_2/in_2')
// (12, 5, 'sp12_v_b_11')
// (12, 5, 'sp4_v_b_21')
// (12, 6, 'local_g2_0')
// (12, 6, 'lutff_2/in_0')
// (12, 6, 'sp12_v_b_8')
// (12, 6, 'sp4_v_b_8')
// (12, 6, 'sp4_v_t_37')
// (12, 7, 'sp12_v_b_7')
// (12, 7, 'sp4_v_b_37')
// (12, 8, 'sp12_v_b_4')
// (12, 8, 'sp4_v_b_24')
// (12, 9, 'local_g1_0')
// (12, 9, 'lutff_3/in_2')
// (12, 9, 'neigh_op_top_0')
// (12, 9, 'sp12_v_b_3')
// (12, 9, 'sp4_v_b_13')
// (12, 10, 'lutff_0/out')
// (12, 10, 'sp12_v_b_0')
// (12, 10, 'sp4_v_b_0')
// (12, 11, 'neigh_op_bot_0')
// (13, 9, 'neigh_op_tnl_0')
// (13, 10, 'neigh_op_lft_0')
// (13, 11, 'neigh_op_bnl_0')

wire n1549;
// (11, 3, 'sp4_r_v_b_47')
// (11, 4, 'local_g0_1')
// (11, 4, 'lutff_5/in_2')
// (11, 4, 'sp4_r_v_b_34')
// (11, 5, 'sp4_r_v_b_23')
// (11, 6, 'sp4_r_v_b_10')
// (12, 2, 'sp4_h_r_10')
// (12, 2, 'sp4_v_t_47')
// (12, 3, 'sp4_v_b_47')
// (12, 4, 'sp4_v_b_34')
// (12, 5, 'sp4_v_b_23')
// (12, 6, 'sp4_v_b_10')
// (13, 1, 'neigh_op_tnr_1')
// (13, 2, 'neigh_op_rgt_1')
// (13, 2, 'sp4_h_r_23')
// (13, 3, 'neigh_op_bnr_1')
// (14, 1, 'neigh_op_top_1')
// (14, 2, 'lutff_1/out')
// (14, 2, 'sp4_h_r_34')
// (14, 3, 'neigh_op_bot_1')
// (15, 1, 'neigh_op_tnl_1')
// (15, 2, 'local_g1_1')
// (15, 2, 'lutff_6/in_2')
// (15, 2, 'neigh_op_lft_1')
// (15, 2, 'sp4_h_r_47')
// (15, 3, 'neigh_op_bnl_1')
// (16, 2, 'sp4_h_l_47')

wire n1550;
// (11, 4, 'local_g0_2')
// (11, 4, 'lutff_1/in_1')
// (11, 4, 'sp4_h_r_2')
// (12, 4, 'sp4_h_r_15')
// (13, 1, 'neigh_op_tnr_0')
// (13, 2, 'local_g2_0')
// (13, 2, 'lutff_4/in_2')
// (13, 2, 'lutff_5/in_3')
// (13, 2, 'lutff_6/in_0')
// (13, 2, 'neigh_op_rgt_0')
// (13, 3, 'neigh_op_bnr_0')
// (13, 4, 'sp4_h_r_26')
// (14, 1, 'neigh_op_top_0')
// (14, 1, 'sp4_r_v_b_44')
// (14, 2, 'local_g0_0')
// (14, 2, 'lutff_0/out')
// (14, 2, 'lutff_1/in_1')
// (14, 2, 'lutff_5/in_1')
// (14, 2, 'lutff_6/in_2')
// (14, 2, 'sp4_r_v_b_33')
// (14, 3, 'neigh_op_bot_0')
// (14, 3, 'sp4_r_v_b_20')
// (14, 4, 'sp4_h_r_39')
// (14, 4, 'sp4_r_v_b_9')
// (15, 0, 'span4_vert_44')
// (15, 1, 'neigh_op_tnl_0')
// (15, 1, 'sp4_v_b_44')
// (15, 2, 'neigh_op_lft_0')
// (15, 2, 'sp4_v_b_33')
// (15, 3, 'neigh_op_bnl_0')
// (15, 3, 'sp4_v_b_20')
// (15, 4, 'sp4_h_l_39')
// (15, 4, 'sp4_v_b_9')

wire n1551;
// (11, 4, 'neigh_op_tnr_6')
// (11, 5, 'neigh_op_rgt_6')
// (11, 6, 'neigh_op_bnr_6')
// (12, 4, 'neigh_op_top_6')
// (12, 5, 'local_g0_6')
// (12, 5, 'lutff_2/in_0')
// (12, 5, 'lutff_6/out')
// (12, 6, 'neigh_op_bot_6')
// (13, 4, 'neigh_op_tnl_6')
// (13, 5, 'neigh_op_lft_6')
// (13, 6, 'neigh_op_bnl_6')

wire n1552;
// (11, 4, 'neigh_op_tnr_7')
// (11, 5, 'neigh_op_rgt_7')
// (11, 6, 'neigh_op_bnr_7')
// (12, 3, 'sp4_r_v_b_39')
// (12, 4, 'neigh_op_top_7')
// (12, 4, 'sp4_r_v_b_26')
// (12, 5, 'lutff_7/out')
// (12, 5, 'sp4_r_v_b_15')
// (12, 6, 'neigh_op_bot_7')
// (12, 6, 'sp4_r_v_b_2')
// (13, 2, 'sp4_h_r_2')
// (13, 2, 'sp4_h_r_7')
// (13, 2, 'sp4_v_t_39')
// (13, 3, 'sp4_v_b_39')
// (13, 4, 'neigh_op_tnl_7')
// (13, 4, 'sp4_v_b_26')
// (13, 5, 'neigh_op_lft_7')
// (13, 5, 'sp4_v_b_15')
// (13, 6, 'neigh_op_bnl_7')
// (13, 6, 'sp4_v_b_2')
// (14, 2, 'sp4_h_r_15')
// (14, 2, 'sp4_h_r_18')
// (15, 2, 'local_g2_2')
// (15, 2, 'lutff_global/cen')
// (15, 2, 'sp4_h_r_26')
// (15, 2, 'sp4_h_r_31')
// (16, 2, 'local_g2_2')
// (16, 2, 'lutff_global/cen')
// (16, 2, 'sp4_h_r_39')
// (16, 2, 'sp4_h_r_42')
// (17, 2, 'sp4_h_l_39')
// (17, 2, 'sp4_h_l_42')

reg n1553 = 0;
// (11, 4, 'sp4_r_v_b_36')
// (11, 5, 'sp4_r_v_b_25')
// (11, 6, 'sp4_r_v_b_12')
// (11, 7, 'sp4_r_v_b_1')
// (11, 8, 'sp4_r_v_b_36')
// (11, 9, 'sp4_r_v_b_25')
// (11, 10, 'sp4_r_v_b_12')
// (11, 11, 'sp4_r_v_b_1')
// (11, 12, 'sp4_r_v_b_47')
// (11, 13, 'sp4_r_v_b_34')
// (11, 14, 'sp4_r_v_b_23')
// (11, 15, 'sp4_r_v_b_10')
// (11, 16, 'sp4_r_v_b_39')
// (11, 17, 'sp4_r_v_b_26')
// (11, 18, 'neigh_op_tnr_1')
// (11, 18, 'sp4_r_v_b_15')
// (11, 19, 'neigh_op_rgt_1')
// (11, 19, 'sp4_r_v_b_2')
// (11, 20, 'neigh_op_bnr_1')
// (12, 3, 'sp4_h_r_6')
// (12, 3, 'sp4_v_t_36')
// (12, 4, 'sp4_v_b_36')
// (12, 5, 'sp4_v_b_25')
// (12, 6, 'sp4_v_b_12')
// (12, 7, 'sp4_v_b_1')
// (12, 7, 'sp4_v_t_36')
// (12, 8, 'sp4_v_b_36')
// (12, 9, 'sp4_v_b_25')
// (12, 10, 'sp4_v_b_12')
// (12, 11, 'sp4_v_b_1')
// (12, 11, 'sp4_v_t_47')
// (12, 12, 'sp4_v_b_47')
// (12, 13, 'sp4_v_b_34')
// (12, 14, 'sp4_v_b_23')
// (12, 15, 'sp4_v_b_10')
// (12, 15, 'sp4_v_t_39')
// (12, 16, 'sp4_v_b_39')
// (12, 17, 'sp4_v_b_26')
// (12, 18, 'neigh_op_top_1')
// (12, 18, 'sp4_v_b_15')
// (12, 19, 'lutff_1/out')
// (12, 19, 'sp4_v_b_2')
// (12, 20, 'neigh_op_bot_1')
// (13, 3, 'local_g1_3')
// (13, 3, 'lutff_1/in_3')
// (13, 3, 'sp4_h_r_19')
// (13, 18, 'local_g2_1')
// (13, 18, 'lutff_5/in_2')
// (13, 18, 'neigh_op_tnl_1')
// (13, 19, 'local_g0_1')
// (13, 19, 'lutff_2/in_1')
// (13, 19, 'neigh_op_lft_1')
// (13, 20, 'local_g2_1')
// (13, 20, 'lutff_2/in_1')
// (13, 20, 'neigh_op_bnl_1')
// (14, 3, 'sp4_h_r_30')
// (15, 3, 'sp4_h_r_43')
// (16, 3, 'sp4_h_l_43')

reg n1554 = 0;
// (11, 4, 'sp4_r_v_b_41')
// (11, 5, 'sp4_r_v_b_28')
// (11, 6, 'sp4_r_v_b_17')
// (11, 7, 'sp4_r_v_b_4')
// (12, 3, 'sp4_h_r_4')
// (12, 3, 'sp4_v_t_41')
// (12, 4, 'sp4_v_b_41')
// (12, 5, 'sp4_v_b_28')
// (12, 6, 'local_g1_1')
// (12, 6, 'lutff_6/in_2')
// (12, 6, 'sp4_v_b_17')
// (12, 7, 'sp4_v_b_4')
// (13, 2, 'neigh_op_tnr_6')
// (13, 3, 'local_g2_6')
// (13, 3, 'lutff_7/in_1')
// (13, 3, 'neigh_op_rgt_6')
// (13, 3, 'sp4_h_r_17')
// (13, 3, 'sp4_r_v_b_44')
// (13, 4, 'neigh_op_bnr_6')
// (13, 4, 'sp4_r_v_b_33')
// (13, 5, 'sp4_r_v_b_20')
// (13, 6, 'local_g2_1')
// (13, 6, 'lutff_0/in_3')
// (13, 6, 'sp4_r_v_b_9')
// (14, 2, 'neigh_op_top_6')
// (14, 2, 'sp4_v_t_44')
// (14, 3, 'lutff_6/out')
// (14, 3, 'sp4_h_r_28')
// (14, 3, 'sp4_v_b_44')
// (14, 4, 'neigh_op_bot_6')
// (14, 4, 'sp4_v_b_33')
// (14, 5, 'sp4_v_b_20')
// (14, 6, 'sp4_v_b_9')
// (15, 2, 'neigh_op_tnl_6')
// (15, 3, 'neigh_op_lft_6')
// (15, 3, 'sp4_h_r_41')
// (15, 4, 'neigh_op_bnl_6')
// (16, 3, 'sp4_h_l_41')

reg n1555 = 0;
// (11, 4, 'sp4_r_v_b_46')
// (11, 5, 'sp4_r_v_b_35')
// (11, 6, 'sp4_r_v_b_22')
// (11, 7, 'sp4_r_v_b_11')
// (12, 3, 'sp4_h_r_5')
// (12, 3, 'sp4_v_t_46')
// (12, 4, 'sp4_v_b_46')
// (12, 5, 'sp4_v_b_35')
// (12, 6, 'local_g1_6')
// (12, 6, 'lutff_4/in_3')
// (12, 6, 'sp4_v_b_22')
// (12, 7, 'sp4_v_b_11')
// (13, 3, 'sp4_h_r_16')
// (14, 3, 'sp4_h_r_29')
// (15, 1, 'sp4_r_v_b_24')
// (15, 1, 'sp4_r_v_b_40')
// (15, 2, 'local_g2_0')
// (15, 2, 'lutff_5/in_3')
// (15, 2, 'neigh_op_tnr_0')
// (15, 2, 'sp4_r_v_b_13')
// (15, 2, 'sp4_r_v_b_29')
// (15, 3, 'neigh_op_rgt_0')
// (15, 3, 'sp4_h_r_40')
// (15, 3, 'sp4_r_v_b_0')
// (15, 3, 'sp4_r_v_b_16')
// (15, 4, 'neigh_op_bnr_0')
// (15, 4, 'sp4_r_v_b_5')
// (15, 5, 'sp4_r_v_b_45')
// (15, 6, 'sp4_r_v_b_32')
// (15, 7, 'sp4_r_v_b_21')
// (15, 8, 'local_g2_0')
// (15, 8, 'lutff_3/in_3')
// (15, 8, 'sp4_r_v_b_8')
// (16, 0, 'span4_vert_24')
// (16, 0, 'span4_vert_40')
// (16, 1, 'sp4_v_b_24')
// (16, 1, 'sp4_v_b_40')
// (16, 2, 'neigh_op_top_0')
// (16, 2, 'sp4_v_b_13')
// (16, 2, 'sp4_v_b_29')
// (16, 3, 'lutff_0/out')
// (16, 3, 'sp4_h_l_40')
// (16, 3, 'sp4_v_b_0')
// (16, 3, 'sp4_v_b_16')
// (16, 4, 'neigh_op_bot_0')
// (16, 4, 'sp4_v_b_5')
// (16, 4, 'sp4_v_t_45')
// (16, 5, 'sp4_v_b_45')
// (16, 6, 'sp4_v_b_32')
// (16, 7, 'sp4_v_b_21')
// (16, 8, 'sp4_v_b_8')
// (17, 2, 'neigh_op_tnl_0')
// (17, 3, 'neigh_op_lft_0')
// (17, 4, 'neigh_op_bnl_0')

reg n1556 = 0;
// (11, 4, 'sp4_r_v_b_47')
// (11, 5, 'sp4_r_v_b_34')
// (11, 6, 'sp4_r_v_b_23')
// (11, 7, 'sp4_r_v_b_10')
// (11, 8, 'sp4_r_v_b_47')
// (11, 9, 'sp4_r_v_b_34')
// (11, 10, 'sp4_r_v_b_23')
// (11, 11, 'sp4_r_v_b_10')
// (12, 3, 'sp4_v_t_47')
// (12, 4, 'sp4_v_b_47')
// (12, 5, 'sp4_v_b_34')
// (12, 6, 'local_g0_7')
// (12, 6, 'lutff_4/in_1')
// (12, 6, 'sp4_v_b_23')
// (12, 7, 'sp4_v_b_10')
// (12, 7, 'sp4_v_t_47')
// (12, 8, 'sp4_v_b_47')
// (12, 9, 'sp4_v_b_34')
// (12, 10, 'sp4_v_b_23')
// (12, 11, 'sp4_h_r_10')
// (12, 11, 'sp4_v_b_10')
// (13, 9, 'sp4_r_v_b_42')
// (13, 10, 'local_g2_1')
// (13, 10, 'lutff_1/in_2')
// (13, 10, 'neigh_op_tnr_1')
// (13, 10, 'sp4_r_v_b_31')
// (13, 11, 'neigh_op_rgt_1')
// (13, 11, 'sp4_h_r_23')
// (13, 11, 'sp4_r_v_b_18')
// (13, 12, 'neigh_op_bnr_1')
// (13, 12, 'sp4_r_v_b_7')
// (13, 13, 'sp4_r_v_b_42')
// (13, 14, 'sp4_r_v_b_31')
// (13, 15, 'sp4_r_v_b_18')
// (13, 16, 'sp4_r_v_b_7')
// (14, 8, 'local_g1_0')
// (14, 8, 'lutff_7/in_2')
// (14, 8, 'sp4_h_r_0')
// (14, 8, 'sp4_v_t_42')
// (14, 9, 'sp4_v_b_42')
// (14, 10, 'neigh_op_top_1')
// (14, 10, 'sp4_v_b_31')
// (14, 11, 'lutff_1/out')
// (14, 11, 'sp4_h_r_34')
// (14, 11, 'sp4_v_b_18')
// (14, 12, 'neigh_op_bot_1')
// (14, 12, 'sp4_v_b_7')
// (14, 12, 'sp4_v_t_42')
// (14, 13, 'sp4_v_b_42')
// (14, 14, 'local_g3_7')
// (14, 14, 'lutff_0/in_0')
// (14, 14, 'sp4_v_b_31')
// (14, 15, 'sp4_v_b_18')
// (14, 16, 'sp4_v_b_7')
// (15, 8, 'sp4_h_r_13')
// (15, 10, 'neigh_op_tnl_1')
// (15, 11, 'neigh_op_lft_1')
// (15, 11, 'sp4_h_r_47')
// (15, 12, 'neigh_op_bnl_1')
// (16, 8, 'sp4_h_r_24')
// (16, 11, 'sp4_h_l_47')
// (17, 8, 'sp4_h_r_37')
// (18, 8, 'sp4_h_l_37')

wire n1557;
// (11, 5, 'neigh_op_tnr_1')
// (11, 6, 'neigh_op_rgt_1')
// (11, 7, 'local_g0_1')
// (11, 7, 'lutff_7/in_0')
// (11, 7, 'neigh_op_bnr_1')
// (12, 5, 'neigh_op_top_1')
// (12, 6, 'lutff_1/out')
// (12, 7, 'neigh_op_bot_1')
// (13, 5, 'neigh_op_tnl_1')
// (13, 6, 'neigh_op_lft_1')
// (13, 7, 'neigh_op_bnl_1')

wire n1558;
// (11, 5, 'neigh_op_tnr_2')
// (11, 6, 'neigh_op_rgt_2')
// (11, 7, 'neigh_op_bnr_2')
// (12, 5, 'neigh_op_top_2')
// (12, 6, 'local_g3_2')
// (12, 6, 'lutff_2/out')
// (12, 6, 'lutff_6/in_3')
// (12, 7, 'neigh_op_bot_2')
// (13, 5, 'neigh_op_tnl_2')
// (13, 6, 'neigh_op_lft_2')
// (13, 7, 'neigh_op_bnl_2')

wire n1559;
// (11, 5, 'neigh_op_tnr_3')
// (11, 6, 'neigh_op_rgt_3')
// (11, 7, 'neigh_op_bnr_3')
// (12, 5, 'neigh_op_top_3')
// (12, 6, 'local_g0_3')
// (12, 6, 'lutff_0/in_3')
// (12, 6, 'lutff_3/out')
// (12, 7, 'neigh_op_bot_3')
// (13, 5, 'neigh_op_tnl_3')
// (13, 6, 'neigh_op_lft_3')
// (13, 7, 'neigh_op_bnl_3')

wire n1560;
// (11, 5, 'neigh_op_tnr_4')
// (11, 6, 'neigh_op_rgt_4')
// (11, 7, 'neigh_op_bnr_4')
// (12, 5, 'neigh_op_top_4')
// (12, 5, 'sp4_r_v_b_36')
// (12, 6, 'lutff_4/out')
// (12, 6, 'sp4_r_v_b_25')
// (12, 7, 'neigh_op_bot_4')
// (12, 7, 'sp4_r_v_b_12')
// (12, 8, 'sp4_r_v_b_1')
// (13, 4, 'sp4_v_t_36')
// (13, 5, 'neigh_op_tnl_4')
// (13, 5, 'sp4_v_b_36')
// (13, 6, 'neigh_op_lft_4')
// (13, 6, 'sp4_v_b_25')
// (13, 7, 'neigh_op_bnl_4')
// (13, 7, 'sp4_v_b_12')
// (13, 8, 'local_g1_1')
// (13, 8, 'lutff_2/in_2')
// (13, 8, 'sp4_v_b_1')

wire n1561;
// (11, 5, 'neigh_op_tnr_5')
// (11, 6, 'neigh_op_rgt_5')
// (11, 7, 'neigh_op_bnr_5')
// (12, 5, 'neigh_op_top_5')
// (12, 6, 'lutff_5/out')
// (12, 7, 'neigh_op_bot_5')
// (13, 5, 'neigh_op_tnl_5')
// (13, 6, 'local_g0_5')
// (13, 6, 'lutff_4/in_3')
// (13, 6, 'neigh_op_lft_5')
// (13, 7, 'neigh_op_bnl_5')

wire n1562;
// (11, 5, 'neigh_op_tnr_6')
// (11, 5, 'sp4_r_v_b_41')
// (11, 6, 'neigh_op_rgt_6')
// (11, 6, 'sp4_r_v_b_28')
// (11, 7, 'neigh_op_bnr_6')
// (11, 7, 'sp4_r_v_b_17')
// (11, 8, 'sp4_r_v_b_4')
// (12, 4, 'sp4_v_t_41')
// (12, 5, 'neigh_op_top_6')
// (12, 5, 'sp4_v_b_41')
// (12, 6, 'lutff_6/out')
// (12, 6, 'sp4_v_b_28')
// (12, 7, 'local_g0_1')
// (12, 7, 'lutff_0/in_1')
// (12, 7, 'neigh_op_bot_6')
// (12, 7, 'sp4_v_b_17')
// (12, 8, 'sp4_v_b_4')
// (13, 5, 'neigh_op_tnl_6')
// (13, 6, 'neigh_op_lft_6')
// (13, 7, 'neigh_op_bnl_6')

wire n1563;
// (11, 5, 'sp4_r_v_b_38')
// (11, 6, 'local_g1_3')
// (11, 6, 'lutff_4/in_2')
// (11, 6, 'sp4_r_v_b_27')
// (11, 7, 'sp4_r_v_b_14')
// (11, 8, 'sp4_r_v_b_3')
// (11, 9, 'sp4_r_v_b_41')
// (11, 10, 'sp4_r_v_b_28')
// (11, 11, 'local_g3_1')
// (11, 11, 'lutff_7/in_3')
// (11, 11, 'sp4_r_v_b_17')
// (11, 12, 'sp4_r_v_b_4')
// (11, 13, 'sp4_r_v_b_37')
// (11, 14, 'local_g0_0')
// (11, 14, 'lutff_5/in_1')
// (11, 14, 'sp4_r_v_b_24')
// (11, 15, 'sp4_r_v_b_13')
// (11, 16, 'sp4_r_v_b_0')
// (12, 2, 'sp4_r_v_b_47')
// (12, 3, 'sp4_r_v_b_34')
// (12, 4, 'local_g3_7')
// (12, 4, 'lutff_2/in_0')
// (12, 4, 'sp4_r_v_b_23')
// (12, 4, 'sp4_v_t_38')
// (12, 5, 'sp4_r_v_b_10')
// (12, 5, 'sp4_v_b_38')
// (12, 6, 'sp4_v_b_27')
// (12, 7, 'sp4_v_b_14')
// (12, 8, 'sp4_h_r_10')
// (12, 8, 'sp4_v_b_3')
// (12, 8, 'sp4_v_t_41')
// (12, 9, 'sp4_v_b_41')
// (12, 10, 'local_g3_4')
// (12, 10, 'lutff_1/in_2')
// (12, 10, 'sp4_v_b_28')
// (12, 11, 'sp4_v_b_17')
// (12, 12, 'sp4_v_b_4')
// (12, 12, 'sp4_v_t_37')
// (12, 13, 'sp4_v_b_37')
// (12, 14, 'sp4_v_b_24')
// (12, 15, 'sp4_v_b_13')
// (12, 16, 'sp4_v_b_0')
// (13, 1, 'sp4_v_t_47')
// (13, 2, 'sp4_v_b_47')
// (13, 3, 'sp4_v_b_34')
// (13, 4, 'sp4_v_b_23')
// (13, 5, 'sp4_h_r_5')
// (13, 5, 'sp4_v_b_10')
// (13, 8, 'sp4_h_r_23')
// (13, 15, 'sp4_h_r_5')
// (14, 5, 'sp4_h_r_16')
// (14, 8, 'sp4_h_r_34')
// (14, 15, 'local_g1_0')
// (14, 15, 'lutff_3/in_2')
// (14, 15, 'sp4_h_r_16')
// (15, 4, 'neigh_op_tnr_4')
// (15, 5, 'neigh_op_rgt_4')
// (15, 5, 'sp4_h_r_29')
// (15, 5, 'sp4_r_v_b_40')
// (15, 6, 'neigh_op_bnr_4')
// (15, 6, 'sp4_r_v_b_29')
// (15, 7, 'sp4_r_v_b_16')
// (15, 8, 'sp4_h_r_47')
// (15, 8, 'sp4_r_v_b_5')
// (15, 15, 'sp4_h_r_29')
// (16, 4, 'neigh_op_top_4')
// (16, 4, 'sp4_r_v_b_36')
// (16, 4, 'sp4_v_t_40')
// (16, 5, 'lutff_4/out')
// (16, 5, 'sp4_h_r_40')
// (16, 5, 'sp4_r_v_b_25')
// (16, 5, 'sp4_v_b_40')
// (16, 6, 'neigh_op_bot_4')
// (16, 6, 'sp4_r_v_b_12')
// (16, 6, 'sp4_v_b_29')
// (16, 7, 'sp4_r_v_b_1')
// (16, 7, 'sp4_v_b_16')
// (16, 8, 'sp4_h_l_47')
// (16, 8, 'sp4_r_v_b_41')
// (16, 8, 'sp4_v_b_5')
// (16, 9, 'sp4_r_v_b_28')
// (16, 10, 'sp4_r_v_b_17')
// (16, 11, 'sp4_r_v_b_4')
// (16, 12, 'sp4_r_v_b_37')
// (16, 13, 'sp4_r_v_b_24')
// (16, 14, 'sp4_r_v_b_13')
// (16, 15, 'sp4_h_r_40')
// (16, 15, 'sp4_r_v_b_0')
// (17, 3, 'sp4_v_t_36')
// (17, 4, 'neigh_op_tnl_4')
// (17, 4, 'sp4_v_b_36')
// (17, 5, 'neigh_op_lft_4')
// (17, 5, 'sp4_h_l_40')
// (17, 5, 'sp4_v_b_25')
// (17, 6, 'neigh_op_bnl_4')
// (17, 6, 'sp4_v_b_12')
// (17, 7, 'sp4_v_b_1')
// (17, 7, 'sp4_v_t_41')
// (17, 8, 'sp4_v_b_41')
// (17, 9, 'sp4_v_b_28')
// (17, 10, 'sp4_v_b_17')
// (17, 11, 'sp4_v_b_4')
// (17, 11, 'sp4_v_t_37')
// (17, 12, 'sp4_v_b_37')
// (17, 13, 'sp4_v_b_24')
// (17, 14, 'sp4_v_b_13')
// (17, 15, 'sp4_h_l_40')
// (17, 15, 'sp4_v_b_0')

wire n1564;
// (11, 5, 'sp4_r_v_b_46')
// (11, 6, 'local_g2_3')
// (11, 6, 'lutff_0/in_3')
// (11, 6, 'sp4_r_v_b_35')
// (11, 7, 'local_g3_6')
// (11, 7, 'lutff_1/in_0')
// (11, 7, 'sp4_r_v_b_22')
// (11, 8, 'sp4_r_v_b_11')
// (11, 9, 'sp4_r_v_b_46')
// (11, 10, 'neigh_op_tnr_3')
// (11, 10, 'sp4_r_v_b_35')
// (11, 11, 'local_g2_3')
// (11, 11, 'lutff_6/in_3')
// (11, 11, 'lutff_7/in_0')
// (11, 11, 'neigh_op_rgt_3')
// (11, 11, 'sp4_r_v_b_22')
// (11, 12, 'neigh_op_bnr_3')
// (11, 12, 'sp4_r_v_b_11')
// (12, 4, 'sp4_v_t_46')
// (12, 5, 'local_g3_6')
// (12, 5, 'lutff_7/in_2')
// (12, 5, 'sp4_v_b_46')
// (12, 6, 'local_g2_3')
// (12, 6, 'lutff_7/in_2')
// (12, 6, 'sp4_v_b_35')
// (12, 7, 'sp4_v_b_22')
// (12, 8, 'sp4_v_b_11')
// (12, 8, 'sp4_v_t_46')
// (12, 9, 'sp4_v_b_46')
// (12, 10, 'neigh_op_top_3')
// (12, 10, 'sp4_v_b_35')
// (12, 11, 'lutff_3/out')
// (12, 11, 'sp4_v_b_22')
// (12, 12, 'neigh_op_bot_3')
// (12, 12, 'sp4_v_b_11')
// (13, 10, 'neigh_op_tnl_3')
// (13, 11, 'neigh_op_lft_3')
// (13, 12, 'neigh_op_bnl_3')

wire n1565;
// (11, 5, 'sp4_r_v_b_47')
// (11, 6, 'sp4_r_v_b_34')
// (11, 7, 'local_g3_7')
// (11, 7, 'lutff_2/in_2')
// (11, 7, 'sp4_r_v_b_23')
// (11, 8, 'sp4_r_v_b_10')
// (12, 4, 'sp4_h_r_4')
// (12, 4, 'sp4_v_t_47')
// (12, 5, 'sp4_v_b_47')
// (12, 6, 'sp4_v_b_34')
// (12, 7, 'sp4_v_b_23')
// (12, 8, 'sp4_v_b_10')
// (13, 3, 'neigh_op_tnr_6')
// (13, 4, 'neigh_op_rgt_6')
// (13, 4, 'sp4_h_r_17')
// (13, 5, 'neigh_op_bnr_6')
// (14, 3, 'neigh_op_top_6')
// (14, 4, 'lutff_6/out')
// (14, 4, 'sp4_h_r_28')
// (14, 5, 'neigh_op_bot_6')
// (15, 3, 'neigh_op_tnl_6')
// (15, 4, 'neigh_op_lft_6')
// (15, 4, 'sp4_h_r_41')
// (15, 5, 'neigh_op_bnl_6')
// (16, 4, 'sp4_h_l_41')

wire n1566;
// (11, 6, 'local_g3_1')
// (11, 6, 'lutff_1/in_3')
// (11, 6, 'sp4_r_v_b_41')
// (11, 7, 'sp4_r_v_b_28')
// (11, 8, 'sp4_r_v_b_17')
// (11, 9, 'sp4_r_v_b_4')
// (11, 10, 'neigh_op_tnr_0')
// (11, 10, 'sp4_r_v_b_45')
// (11, 11, 'neigh_op_rgt_0')
// (11, 11, 'sp4_r_v_b_32')
// (11, 12, 'neigh_op_bnr_0')
// (11, 12, 'sp4_r_v_b_21')
// (11, 13, 'sp4_r_v_b_8')
// (12, 5, 'sp4_v_t_41')
// (12, 6, 'sp4_v_b_41')
// (12, 7, 'sp4_v_b_28')
// (12, 8, 'sp4_v_b_17')
// (12, 9, 'sp4_v_b_4')
// (12, 9, 'sp4_v_t_45')
// (12, 10, 'neigh_op_top_0')
// (12, 10, 'sp4_v_b_45')
// (12, 11, 'lutff_0/out')
// (12, 11, 'sp4_v_b_32')
// (12, 12, 'neigh_op_bot_0')
// (12, 12, 'sp4_v_b_21')
// (12, 13, 'sp4_v_b_8')
// (13, 10, 'neigh_op_tnl_0')
// (13, 11, 'neigh_op_lft_0')
// (13, 12, 'neigh_op_bnl_0')

wire n1567;
// (11, 6, 'neigh_op_tnr_0')
// (11, 7, 'neigh_op_rgt_0')
// (11, 8, 'neigh_op_bnr_0')
// (12, 6, 'neigh_op_top_0')
// (12, 7, 'lutff_0/out')
// (12, 8, 'neigh_op_bot_0')
// (13, 6, 'neigh_op_tnl_0')
// (13, 7, 'neigh_op_lft_0')
// (13, 8, 'local_g3_0')
// (13, 8, 'lutff_2/in_3')
// (13, 8, 'neigh_op_bnl_0')

wire n1568;
// (11, 6, 'neigh_op_tnr_1')
// (11, 7, 'neigh_op_rgt_1')
// (11, 8, 'neigh_op_bnr_1')
// (12, 6, 'neigh_op_top_1')
// (12, 7, 'lutff_1/out')
// (12, 8, 'neigh_op_bot_1')
// (13, 6, 'neigh_op_tnl_1')
// (13, 7, 'local_g0_1')
// (13, 7, 'lutff_3/in_0')
// (13, 7, 'neigh_op_lft_1')
// (13, 8, 'neigh_op_bnl_1')

wire n1569;
// (11, 6, 'neigh_op_tnr_2')
// (11, 7, 'neigh_op_rgt_2')
// (11, 8, 'neigh_op_bnr_2')
// (12, 6, 'neigh_op_top_2')
// (12, 7, 'lutff_2/out')
// (12, 8, 'local_g1_2')
// (12, 8, 'lutff_1/in_2')
// (12, 8, 'neigh_op_bot_2')
// (13, 6, 'neigh_op_tnl_2')
// (13, 7, 'neigh_op_lft_2')
// (13, 8, 'neigh_op_bnl_2')

reg n1570 = 0;
// (11, 6, 'neigh_op_tnr_3')
// (11, 7, 'neigh_op_rgt_3')
// (11, 8, 'neigh_op_bnr_3')
// (12, 6, 'local_g1_3')
// (12, 6, 'lutff_1/in_1')
// (12, 6, 'lutff_5/in_3')
// (12, 6, 'neigh_op_top_3')
// (12, 7, 'local_g0_3')
// (12, 7, 'lutff_3/out')
// (12, 7, 'lutff_4/in_1')
// (12, 8, 'neigh_op_bot_3')
// (13, 6, 'neigh_op_tnl_3')
// (13, 7, 'neigh_op_lft_3')
// (13, 8, 'neigh_op_bnl_3')

wire n1571;
// (11, 6, 'neigh_op_tnr_4')
// (11, 7, 'neigh_op_rgt_4')
// (11, 8, 'neigh_op_bnr_4')
// (12, 6, 'neigh_op_top_4')
// (12, 7, 'lutff_4/out')
// (12, 8, 'local_g1_4')
// (12, 8, 'lutff_7/in_2')
// (12, 8, 'neigh_op_bot_4')
// (13, 6, 'neigh_op_tnl_4')
// (13, 7, 'neigh_op_lft_4')
// (13, 8, 'neigh_op_bnl_4')

wire n1572;
// (11, 6, 'neigh_op_tnr_5')
// (11, 7, 'neigh_op_rgt_5')
// (11, 8, 'neigh_op_bnr_5')
// (12, 6, 'neigh_op_top_5')
// (12, 7, 'local_g3_5')
// (12, 7, 'lutff_4/in_0')
// (12, 7, 'lutff_5/out')
// (12, 8, 'neigh_op_bot_5')
// (13, 6, 'neigh_op_tnl_5')
// (13, 7, 'neigh_op_lft_5')
// (13, 8, 'neigh_op_bnl_5')

reg n1573 = 0;
// (11, 6, 'neigh_op_tnr_6')
// (11, 7, 'neigh_op_rgt_6')
// (11, 7, 'sp4_h_r_1')
// (11, 8, 'neigh_op_bnr_6')
// (12, 6, 'neigh_op_top_6')
// (12, 7, 'local_g2_6')
// (12, 7, 'lutff_6/out')
// (12, 7, 'lutff_7/in_3')
// (12, 7, 'sp4_h_r_12')
// (12, 8, 'neigh_op_bot_6')
// (13, 6, 'neigh_op_tnl_6')
// (13, 7, 'neigh_op_lft_6')
// (13, 7, 'sp4_h_r_25')
// (13, 8, 'neigh_op_bnl_6')
// (14, 7, 'local_g3_4')
// (14, 7, 'lutff_3/in_0')
// (14, 7, 'sp4_h_r_36')
// (15, 7, 'local_g1_4')
// (15, 7, 'lutff_2/in_1')
// (15, 7, 'sp4_h_l_36')
// (15, 7, 'sp4_h_r_4')
// (16, 7, 'sp4_h_r_17')
// (17, 7, 'sp4_h_r_28')
// (18, 7, 'sp4_h_r_41')
// (19, 7, 'sp4_h_l_41')

wire n1574;
// (11, 6, 'sp4_r_v_b_40')
// (11, 7, 'local_g0_5')
// (11, 7, 'lutff_0/in_1')
// (11, 7, 'sp4_r_v_b_29')
// (11, 8, 'sp4_r_v_b_16')
// (11, 9, 'sp4_r_v_b_5')
// (12, 4, 'neigh_op_tnr_3')
// (12, 5, 'neigh_op_rgt_3')
// (12, 5, 'sp4_h_r_11')
// (12, 5, 'sp4_v_t_40')
// (12, 6, 'neigh_op_bnr_3')
// (12, 6, 'sp4_v_b_40')
// (12, 7, 'sp4_v_b_29')
// (12, 8, 'sp4_v_b_16')
// (12, 9, 'sp4_v_b_5')
// (13, 4, 'neigh_op_top_3')
// (13, 5, 'lutff_3/out')
// (13, 5, 'sp4_h_r_22')
// (13, 6, 'neigh_op_bot_3')
// (14, 4, 'neigh_op_tnl_3')
// (14, 5, 'neigh_op_lft_3')
// (14, 5, 'sp4_h_r_35')
// (14, 6, 'neigh_op_bnl_3')
// (15, 5, 'sp4_h_r_46')
// (16, 5, 'sp4_h_l_46')

reg n1575 = 0;
// (11, 7, 'local_g2_4')
// (11, 7, 'lutff_3/in_3')
// (11, 7, 'neigh_op_tnr_4')
// (11, 8, 'local_g3_4')
// (11, 8, 'lutff_4/in_3')
// (11, 8, 'neigh_op_rgt_4')
// (11, 9, 'neigh_op_bnr_4')
// (12, 7, 'neigh_op_top_4')
// (12, 8, 'local_g2_4')
// (12, 8, 'lutff_3/in_1')
// (12, 8, 'lutff_4/out')
// (12, 8, 'lutff_7/in_3')
// (12, 9, 'neigh_op_bot_4')
// (13, 7, 'neigh_op_tnl_4')
// (13, 8, 'neigh_op_lft_4')
// (13, 9, 'neigh_op_bnl_4')

reg n1576 = 0;
// (11, 7, 'local_g2_6')
// (11, 7, 'lutff_4/in_2')
// (11, 7, 'lutff_7/in_3')
// (11, 7, 'neigh_op_tnr_6')
// (11, 8, 'neigh_op_rgt_6')
// (11, 9, 'neigh_op_bnr_6')
// (12, 7, 'local_g1_6')
// (12, 7, 'lutff_2/in_1')
// (12, 7, 'lutff_5/in_0')
// (12, 7, 'neigh_op_top_6')
// (12, 8, 'lutff_6/out')
// (12, 9, 'neigh_op_bot_6')
// (13, 7, 'neigh_op_tnl_6')
// (13, 8, 'neigh_op_lft_6')
// (13, 9, 'neigh_op_bnl_6')

reg n1577 = 0;
// (11, 7, 'local_g3_1')
// (11, 7, 'lutff_0/in_0')
// (11, 7, 'sp4_r_v_b_41')
// (11, 8, 'local_g1_4')
// (11, 8, 'lutff_7/in_2')
// (11, 8, 'sp4_r_v_b_28')
// (11, 9, 'neigh_op_tnr_2')
// (11, 9, 'sp4_r_v_b_17')
// (11, 10, 'neigh_op_rgt_2')
// (11, 10, 'sp4_r_v_b_4')
// (11, 11, 'neigh_op_bnr_2')
// (12, 6, 'sp4_v_t_41')
// (12, 7, 'sp4_v_b_41')
// (12, 8, 'sp4_v_b_28')
// (12, 9, 'local_g0_2')
// (12, 9, 'lutff_0/in_0')
// (12, 9, 'lutff_7/in_1')
// (12, 9, 'neigh_op_top_2')
// (12, 9, 'sp4_v_b_17')
// (12, 10, 'lutff_2/out')
// (12, 10, 'sp4_v_b_4')
// (12, 11, 'neigh_op_bot_2')
// (13, 9, 'neigh_op_tnl_2')
// (13, 10, 'neigh_op_lft_2')
// (13, 11, 'neigh_op_bnl_2')

wire n1578;
// (11, 7, 'neigh_op_tnr_1')
// (11, 8, 'neigh_op_rgt_1')
// (11, 9, 'neigh_op_bnr_1')
// (12, 7, 'neigh_op_top_1')
// (12, 8, 'lutff_1/out')
// (12, 9, 'local_g0_1')
// (12, 9, 'lutff_1/in_2')
// (12, 9, 'neigh_op_bot_1')
// (13, 7, 'neigh_op_tnl_1')
// (13, 8, 'neigh_op_lft_1')
// (13, 9, 'neigh_op_bnl_1')

reg n1579 = 0;
// (11, 7, 'neigh_op_tnr_2')
// (11, 8, 'local_g3_2')
// (11, 8, 'lutff_2/in_1')
// (11, 8, 'neigh_op_rgt_2')
// (11, 9, 'neigh_op_bnr_2')
// (12, 7, 'neigh_op_top_2')
// (12, 8, 'lutff_2/out')
// (12, 9, 'neigh_op_bot_2')
// (13, 7, 'local_g2_2')
// (13, 7, 'lutff_1/in_1')
// (13, 7, 'neigh_op_tnl_2')
// (13, 8, 'local_g1_2')
// (13, 8, 'lutff_4/in_1')
// (13, 8, 'lutff_7/in_0')
// (13, 8, 'neigh_op_lft_2')
// (13, 9, 'neigh_op_bnl_2')

wire n1580;
// (11, 7, 'neigh_op_tnr_3')
// (11, 8, 'neigh_op_rgt_3')
// (11, 9, 'neigh_op_bnr_3')
// (12, 7, 'neigh_op_top_3')
// (12, 8, 'lutff_3/out')
// (12, 9, 'local_g1_3')
// (12, 9, 'lutff_1/in_1')
// (12, 9, 'neigh_op_bot_3')
// (13, 7, 'neigh_op_tnl_3')
// (13, 8, 'neigh_op_lft_3')
// (13, 9, 'neigh_op_bnl_3')

wire n1581;
// (11, 7, 'neigh_op_tnr_5')
// (11, 8, 'neigh_op_rgt_5')
// (11, 9, 'neigh_op_bnr_5')
// (12, 7, 'local_g0_5')
// (12, 7, 'lutff_0/in_3')
// (12, 7, 'neigh_op_top_5')
// (12, 8, 'lutff_5/out')
// (12, 9, 'neigh_op_bot_5')
// (13, 7, 'neigh_op_tnl_5')
// (13, 8, 'neigh_op_lft_5')
// (13, 9, 'neigh_op_bnl_5')

wire n1582;
// (11, 7, 'neigh_op_tnr_7')
// (11, 8, 'neigh_op_rgt_7')
// (11, 9, 'neigh_op_bnr_7')
// (12, 7, 'neigh_op_top_7')
// (12, 8, 'lutff_7/out')
// (12, 9, 'neigh_op_bot_7')
// (13, 7, 'neigh_op_tnl_7')
// (13, 8, 'local_g1_7')
// (13, 8, 'lutff_2/in_0')
// (13, 8, 'neigh_op_lft_7')
// (13, 9, 'neigh_op_bnl_7')

wire n1583;
// (11, 8, 'neigh_op_tnr_0')
// (11, 9, 'neigh_op_rgt_0')
// (11, 10, 'neigh_op_bnr_0')
// (12, 8, 'local_g1_0')
// (12, 8, 'lutff_5/in_0')
// (12, 8, 'neigh_op_top_0')
// (12, 9, 'lutff_0/out')
// (12, 10, 'neigh_op_bot_0')
// (13, 8, 'neigh_op_tnl_0')
// (13, 9, 'neigh_op_lft_0')
// (13, 10, 'neigh_op_bnl_0')

wire n1584;
// (11, 8, 'neigh_op_tnr_1')
// (11, 9, 'neigh_op_rgt_1')
// (11, 10, 'neigh_op_bnr_1')
// (12, 8, 'neigh_op_top_1')
// (12, 9, 'local_g3_1')
// (12, 9, 'lutff_1/out')
// (12, 9, 'lutff_2/in_0')
// (12, 10, 'neigh_op_bot_1')
// (13, 8, 'neigh_op_tnl_1')
// (13, 9, 'neigh_op_lft_1')
// (13, 10, 'neigh_op_bnl_1')

wire n1585;
// (11, 8, 'neigh_op_tnr_2')
// (11, 9, 'neigh_op_rgt_2')
// (11, 10, 'neigh_op_bnr_2')
// (12, 8, 'neigh_op_top_2')
// (12, 9, 'lutff_2/out')
// (12, 10, 'neigh_op_bot_2')
// (13, 8, 'neigh_op_tnl_2')
// (13, 9, 'local_g1_2')
// (13, 9, 'lutff_0/in_3')
// (13, 9, 'neigh_op_lft_2')
// (13, 10, 'neigh_op_bnl_2')

wire n1586;
// (11, 8, 'neigh_op_tnr_3')
// (11, 9, 'neigh_op_rgt_3')
// (11, 10, 'neigh_op_bnr_3')
// (12, 8, 'neigh_op_top_3')
// (12, 9, 'local_g3_3')
// (12, 9, 'lutff_1/in_3')
// (12, 9, 'lutff_3/out')
// (12, 10, 'neigh_op_bot_3')
// (13, 8, 'neigh_op_tnl_3')
// (13, 9, 'neigh_op_lft_3')
// (13, 10, 'neigh_op_bnl_3')

wire n1587;
// (11, 8, 'neigh_op_tnr_4')
// (11, 9, 'neigh_op_rgt_4')
// (11, 10, 'neigh_op_bnr_4')
// (12, 8, 'neigh_op_top_4')
// (12, 9, 'local_g3_4')
// (12, 9, 'lutff_1/in_0')
// (12, 9, 'lutff_4/out')
// (12, 10, 'neigh_op_bot_4')
// (13, 8, 'neigh_op_tnl_4')
// (13, 9, 'neigh_op_lft_4')
// (13, 10, 'neigh_op_bnl_4')

wire n1588;
// (11, 8, 'neigh_op_tnr_5')
// (11, 9, 'neigh_op_rgt_5')
// (11, 10, 'neigh_op_bnr_5')
// (12, 8, 'neigh_op_top_5')
// (12, 9, 'local_g3_5')
// (12, 9, 'lutff_4/in_0')
// (12, 9, 'lutff_5/out')
// (12, 10, 'neigh_op_bot_5')
// (13, 8, 'neigh_op_tnl_5')
// (13, 9, 'neigh_op_lft_5')
// (13, 10, 'neigh_op_bnl_5')

reg n1589 = 0;
// (11, 8, 'neigh_op_tnr_6')
// (11, 9, 'neigh_op_rgt_6')
// (11, 9, 'sp4_r_v_b_44')
// (11, 10, 'neigh_op_bnr_6')
// (11, 10, 'sp4_r_v_b_33')
// (11, 11, 'sp4_r_v_b_20')
// (11, 12, 'sp4_r_v_b_9')
// (11, 13, 'sp4_r_v_b_40')
// (11, 14, 'sp4_r_v_b_29')
// (11, 15, 'sp4_r_v_b_16')
// (11, 16, 'local_g1_5')
// (11, 16, 'lutff_5/in_1')
// (11, 16, 'sp4_r_v_b_5')
// (12, 8, 'neigh_op_top_6')
// (12, 8, 'sp4_v_t_44')
// (12, 9, 'lutff_6/out')
// (12, 9, 'sp4_v_b_44')
// (12, 10, 'neigh_op_bot_6')
// (12, 10, 'sp4_v_b_33')
// (12, 11, 'sp4_v_b_20')
// (12, 12, 'sp4_v_b_9')
// (12, 12, 'sp4_v_t_40')
// (12, 13, 'sp4_v_b_40')
// (12, 14, 'sp4_v_b_29')
// (12, 15, 'sp4_v_b_16')
// (12, 16, 'sp4_v_b_5')
// (13, 8, 'neigh_op_tnl_6')
// (13, 9, 'neigh_op_lft_6')
// (13, 10, 'neigh_op_bnl_6')

wire n1590;
// (11, 8, 'neigh_op_tnr_7')
// (11, 9, 'neigh_op_rgt_7')
// (11, 10, 'neigh_op_bnr_7')
// (12, 8, 'neigh_op_top_7')
// (12, 9, 'local_g2_7')
// (12, 9, 'lutff_2/in_3')
// (12, 9, 'lutff_7/out')
// (12, 10, 'neigh_op_bot_7')
// (13, 8, 'neigh_op_tnl_7')
// (13, 9, 'neigh_op_lft_7')
// (13, 10, 'neigh_op_bnl_7')

wire n1591;
// (11, 8, 'sp4_h_r_9')
// (12, 8, 'sp4_h_r_20')
// (13, 8, 'sp4_h_r_33')
// (14, 8, 'sp4_h_r_44')
// (14, 9, 'sp4_r_v_b_39')
// (14, 10, 'sp4_r_v_b_26')
// (14, 11, 'sp4_r_v_b_15')
// (14, 12, 'sp4_r_v_b_2')
// (15, 8, 'local_g0_2')
// (15, 8, 'lutff_global/cen')
// (15, 8, 'sp4_h_l_44')
// (15, 8, 'sp4_h_r_1')
// (15, 8, 'sp4_h_r_10')
// (15, 8, 'sp4_v_t_39')
// (15, 9, 'sp4_v_b_39')
// (15, 10, 'local_g2_2')
// (15, 10, 'lutff_global/cen')
// (15, 10, 'sp4_v_b_26')
// (15, 11, 'sp4_v_b_15')
// (15, 12, 'sp4_v_b_2')
// (16, 8, 'sp4_h_r_12')
// (16, 8, 'sp4_h_r_23')
// (17, 7, 'neigh_op_tnr_2')
// (17, 8, 'neigh_op_rgt_2')
// (17, 8, 'sp4_h_r_25')
// (17, 8, 'sp4_h_r_34')
// (17, 9, 'local_g0_2')
// (17, 9, 'lutff_global/cen')
// (17, 9, 'neigh_op_bnr_2')
// (18, 5, 'sp4_r_v_b_40')
// (18, 6, 'sp4_r_v_b_29')
// (18, 7, 'neigh_op_top_2')
// (18, 7, 'sp4_r_v_b_16')
// (18, 8, 'lutff_2/out')
// (18, 8, 'sp4_h_r_36')
// (18, 8, 'sp4_h_r_47')
// (18, 8, 'sp4_r_v_b_5')
// (18, 9, 'neigh_op_bot_2')
// (19, 4, 'sp4_v_t_40')
// (19, 5, 'sp4_v_b_40')
// (19, 6, 'sp4_v_b_29')
// (19, 7, 'neigh_op_tnl_2')
// (19, 7, 'sp4_v_b_16')
// (19, 8, 'neigh_op_lft_2')
// (19, 8, 'sp4_h_l_36')
// (19, 8, 'sp4_h_l_47')
// (19, 8, 'sp4_v_b_5')
// (19, 9, 'neigh_op_bnl_2')

reg n1592 = 0;
// (11, 8, 'sp4_r_v_b_39')
// (11, 9, 'sp4_r_v_b_26')
// (11, 10, 'neigh_op_tnr_1')
// (11, 10, 'sp4_r_v_b_15')
// (11, 11, 'neigh_op_rgt_1')
// (11, 11, 'sp4_r_v_b_2')
// (11, 12, 'neigh_op_bnr_1')
// (12, 7, 'local_g1_2')
// (12, 7, 'lutff_1/in_2')
// (12, 7, 'sp4_h_r_2')
// (12, 7, 'sp4_v_t_39')
// (12, 8, 'sp4_r_v_b_38')
// (12, 8, 'sp4_v_b_39')
// (12, 9, 'sp4_r_v_b_27')
// (12, 9, 'sp4_v_b_26')
// (12, 10, 'neigh_op_top_1')
// (12, 10, 'sp4_r_v_b_14')
// (12, 10, 'sp4_v_b_15')
// (12, 11, 'lutff_1/out')
// (12, 11, 'sp4_r_v_b_3')
// (12, 11, 'sp4_v_b_2')
// (12, 12, 'neigh_op_bot_1')
// (13, 7, 'sp4_h_r_15')
// (13, 7, 'sp4_v_t_38')
// (13, 8, 'local_g2_6')
// (13, 8, 'lutff_6/in_2')
// (13, 8, 'sp4_v_b_38')
// (13, 9, 'local_g3_3')
// (13, 9, 'lutff_2/in_0')
// (13, 9, 'sp4_v_b_27')
// (13, 10, 'neigh_op_tnl_1')
// (13, 10, 'sp4_v_b_14')
// (13, 11, 'neigh_op_lft_1')
// (13, 11, 'sp4_v_b_3')
// (13, 12, 'local_g2_1')
// (13, 12, 'lutff_1/in_0')
// (13, 12, 'neigh_op_bnl_1')
// (14, 7, 'sp4_h_r_26')
// (15, 7, 'sp4_h_r_39')
// (16, 7, 'sp4_h_l_39')

reg n1593 = 0;
// (11, 8, 'sp4_r_v_b_45')
// (11, 9, 'sp4_r_v_b_32')
// (11, 10, 'sp4_r_v_b_21')
// (11, 11, 'sp4_r_v_b_8')
// (12, 5, 'sp4_r_v_b_43')
// (12, 6, 'sp4_r_v_b_30')
// (12, 7, 'sp4_h_r_8')
// (12, 7, 'sp4_r_v_b_19')
// (12, 7, 'sp4_v_t_45')
// (12, 8, 'sp4_r_v_b_6')
// (12, 8, 'sp4_v_b_45')
// (12, 9, 'local_g2_6')
// (12, 9, 'lutff_3/in_1')
// (12, 9, 'sp4_r_v_b_38')
// (12, 9, 'sp4_v_b_32')
// (12, 10, 'neigh_op_tnr_7')
// (12, 10, 'sp4_r_v_b_27')
// (12, 10, 'sp4_v_b_21')
// (12, 11, 'neigh_op_rgt_7')
// (12, 11, 'sp4_h_r_3')
// (12, 11, 'sp4_r_v_b_14')
// (12, 11, 'sp4_v_b_8')
// (12, 12, 'neigh_op_bnr_7')
// (12, 12, 'sp4_r_v_b_3')
// (13, 4, 'sp4_v_t_43')
// (13, 5, 'sp4_v_b_43')
// (13, 6, 'sp4_v_b_30')
// (13, 7, 'local_g0_3')
// (13, 7, 'lutff_2/in_1')
// (13, 7, 'sp4_h_r_21')
// (13, 7, 'sp4_v_b_19')
// (13, 8, 'sp4_v_b_6')
// (13, 8, 'sp4_v_t_38')
// (13, 9, 'sp4_r_v_b_39')
// (13, 9, 'sp4_v_b_38')
// (13, 10, 'local_g1_7')
// (13, 10, 'lutff_6/in_0')
// (13, 10, 'neigh_op_top_7')
// (13, 10, 'sp4_r_v_b_26')
// (13, 10, 'sp4_v_b_27')
// (13, 11, 'lutff_7/out')
// (13, 11, 'sp4_h_r_14')
// (13, 11, 'sp4_r_v_b_15')
// (13, 11, 'sp4_v_b_14')
// (13, 12, 'neigh_op_bot_7')
// (13, 12, 'sp4_r_v_b_2')
// (13, 12, 'sp4_v_b_3')
// (14, 7, 'sp4_h_r_32')
// (14, 8, 'sp4_v_t_39')
// (14, 9, 'sp4_v_b_39')
// (14, 10, 'neigh_op_tnl_7')
// (14, 10, 'sp4_v_b_26')
// (14, 11, 'neigh_op_lft_7')
// (14, 11, 'sp4_h_r_27')
// (14, 11, 'sp4_v_b_15')
// (14, 12, 'local_g3_7')
// (14, 12, 'lutff_0/in_2')
// (14, 12, 'neigh_op_bnl_7')
// (14, 12, 'sp4_h_r_2')
// (14, 12, 'sp4_v_b_2')
// (15, 7, 'local_g3_5')
// (15, 7, 'lutff_6/in_2')
// (15, 7, 'sp4_h_r_45')
// (15, 11, 'sp4_h_r_38')
// (15, 12, 'local_g0_7')
// (15, 12, 'lutff_1/in_0')
// (15, 12, 'sp4_h_r_15')
// (16, 7, 'sp4_h_l_45')
// (16, 11, 'sp4_h_l_38')
// (16, 12, 'sp4_h_r_26')
// (17, 12, 'sp4_h_r_39')
// (18, 12, 'sp4_h_l_39')

wire n1594;
// (11, 9, 'sp4_h_r_1')
// (12, 9, 'sp4_h_r_12')
// (13, 9, 'local_g3_1')
// (13, 9, 'lutff_0/in_2')
// (13, 9, 'sp4_h_r_25')
// (14, 9, 'neigh_op_tnr_2')
// (14, 9, 'sp4_h_r_36')
// (14, 10, 'neigh_op_rgt_2')
// (14, 10, 'sp4_r_v_b_36')
// (14, 11, 'neigh_op_bnr_2')
// (14, 11, 'sp4_r_v_b_25')
// (14, 12, 'sp4_r_v_b_12')
// (14, 13, 'sp4_r_v_b_1')
// (15, 9, 'neigh_op_top_2')
// (15, 9, 'sp4_h_l_36')
// (15, 9, 'sp4_v_t_36')
// (15, 10, 'lutff_2/out')
// (15, 10, 'sp4_v_b_36')
// (15, 11, 'neigh_op_bot_2')
// (15, 11, 'sp4_v_b_25')
// (15, 12, 'sp4_v_b_12')
// (15, 13, 'sp4_v_b_1')
// (16, 9, 'neigh_op_tnl_2')
// (16, 10, 'neigh_op_lft_2')
// (16, 11, 'neigh_op_bnl_2')

reg n1595 = 0;
// (11, 9, 'sp4_h_r_10')
// (12, 9, 'sp4_h_r_23')
// (13, 3, 'local_g1_2')
// (13, 3, 'lutff_4/in_3')
// (13, 3, 'sp4_h_r_10')
// (13, 9, 'local_g3_2')
// (13, 9, 'lutff_3/in_2')
// (13, 9, 'sp4_h_r_34')
// (14, 2, 'neigh_op_tnr_1')
// (14, 2, 'sp4_r_v_b_47')
// (14, 3, 'neigh_op_rgt_1')
// (14, 3, 'sp4_h_r_23')
// (14, 3, 'sp4_r_v_b_34')
// (14, 4, 'neigh_op_bnr_1')
// (14, 4, 'sp4_r_v_b_23')
// (14, 4, 'sp4_r_v_b_45')
// (14, 5, 'sp4_r_v_b_10')
// (14, 5, 'sp4_r_v_b_32')
// (14, 6, 'sp4_r_v_b_21')
// (14, 6, 'sp4_r_v_b_47')
// (14, 7, 'sp4_r_v_b_34')
// (14, 7, 'sp4_r_v_b_8')
// (14, 8, 'sp4_r_v_b_23')
// (14, 9, 'local_g2_2')
// (14, 9, 'lutff_0/in_0')
// (14, 9, 'sp4_h_r_47')
// (14, 9, 'sp4_r_v_b_10')
// (15, 0, 'span12_vert_22')
// (15, 1, 'sp12_v_b_22')
// (15, 1, 'sp4_v_t_47')
// (15, 2, 'neigh_op_top_1')
// (15, 2, 'sp12_v_b_21')
// (15, 2, 'sp4_v_b_47')
// (15, 3, 'lutff_1/out')
// (15, 3, 'sp12_v_b_18')
// (15, 3, 'sp4_h_r_2')
// (15, 3, 'sp4_h_r_34')
// (15, 3, 'sp4_v_b_34')
// (15, 3, 'sp4_v_t_45')
// (15, 4, 'neigh_op_bot_1')
// (15, 4, 'sp12_v_b_17')
// (15, 4, 'sp4_v_b_23')
// (15, 4, 'sp4_v_b_45')
// (15, 5, 'sp12_v_b_14')
// (15, 5, 'sp4_v_b_10')
// (15, 5, 'sp4_v_b_32')
// (15, 5, 'sp4_v_t_47')
// (15, 6, 'sp12_v_b_13')
// (15, 6, 'sp4_v_b_21')
// (15, 6, 'sp4_v_b_47')
// (15, 7, 'local_g0_0')
// (15, 7, 'lutff_1/in_1')
// (15, 7, 'sp12_v_b_10')
// (15, 7, 'sp4_v_b_34')
// (15, 7, 'sp4_v_b_8')
// (15, 8, 'sp12_v_b_9')
// (15, 8, 'sp4_v_b_23')
// (15, 9, 'local_g3_6')
// (15, 9, 'lutff_2/in_3')
// (15, 9, 'sp12_v_b_6')
// (15, 9, 'sp4_h_l_47')
// (15, 9, 'sp4_v_b_10')
// (15, 10, 'sp12_v_b_5')
// (15, 11, 'sp12_v_b_2')
// (15, 12, 'sp12_v_b_1')
// (16, 2, 'neigh_op_tnl_1')
// (16, 3, 'neigh_op_lft_1')
// (16, 3, 'sp4_h_r_15')
// (16, 3, 'sp4_h_r_47')
// (16, 4, 'neigh_op_bnl_1')
// (17, 3, 'sp4_h_l_47')
// (17, 3, 'sp4_h_r_26')
// (18, 3, 'sp4_h_r_39')
// (19, 3, 'sp4_h_l_39')

reg n1596 = 0;
// (11, 9, 'sp4_h_r_11')
// (12, 9, 'sp4_h_r_22')
// (13, 8, 'neigh_op_tnr_7')
// (13, 9, 'neigh_op_rgt_7')
// (13, 9, 'sp4_h_r_35')
// (13, 10, 'neigh_op_bnr_7')
// (14, 7, 'sp4_r_v_b_39')
// (14, 8, 'neigh_op_top_7')
// (14, 8, 'sp4_r_v_b_26')
// (14, 9, 'lutff_7/out')
// (14, 9, 'sp4_h_r_46')
// (14, 9, 'sp4_r_v_b_15')
// (14, 10, 'neigh_op_bot_7')
// (14, 10, 'sp4_r_v_b_2')
// (15, 6, 'sp4_v_t_39')
// (15, 7, 'local_g3_7')
// (15, 7, 'lutff_2/in_2')
// (15, 7, 'sp4_v_b_39')
// (15, 8, 'neigh_op_tnl_7')
// (15, 8, 'sp4_v_b_26')
// (15, 9, 'local_g0_7')
// (15, 9, 'lutff_0/in_3')
// (15, 9, 'neigh_op_lft_7')
// (15, 9, 'sp4_h_l_46')
// (15, 9, 'sp4_h_r_2')
// (15, 9, 'sp4_v_b_15')
// (15, 10, 'neigh_op_bnl_7')
// (15, 10, 'sp4_v_b_2')
// (16, 9, 'sp4_h_r_15')
// (17, 9, 'sp4_h_r_26')
// (18, 9, 'local_g2_7')
// (18, 9, 'lutff_6/in_1')
// (18, 9, 'sp4_h_r_39')
// (19, 9, 'sp4_h_l_39')

reg n1597 = 0;
// (11, 9, 'sp4_h_r_5')
// (12, 9, 'sp4_h_r_16')
// (13, 8, 'neigh_op_tnr_4')
// (13, 9, 'neigh_op_rgt_4')
// (13, 9, 'sp4_h_r_29')
// (13, 10, 'neigh_op_bnr_4')
// (14, 8, 'neigh_op_top_4')
// (14, 9, 'lutff_4/out')
// (14, 9, 'sp4_h_r_40')
// (14, 10, 'neigh_op_bot_4')
// (15, 8, 'local_g3_4')
// (15, 8, 'lutff_0/in_1')
// (15, 8, 'lutff_6/in_1')
// (15, 8, 'neigh_op_tnl_4')
// (15, 9, 'neigh_op_lft_4')
// (15, 9, 'sp4_h_l_40')
// (15, 9, 'sp4_h_r_5')
// (15, 10, 'neigh_op_bnl_4')
// (16, 9, 'local_g0_0')
// (16, 9, 'lutff_3/in_1')
// (16, 9, 'sp4_h_r_16')
// (17, 9, 'sp4_h_r_29')
// (18, 9, 'sp4_h_r_40')
// (19, 9, 'sp4_h_l_40')

reg n1598 = 0;
// (11, 9, 'sp4_r_v_b_36')
// (11, 10, 'neigh_op_tnr_6')
// (11, 10, 'sp4_r_v_b_25')
// (11, 11, 'neigh_op_rgt_6')
// (11, 11, 'sp4_r_v_b_12')
// (11, 12, 'neigh_op_bnr_6')
// (11, 12, 'sp4_r_v_b_1')
// (12, 8, 'local_g0_6')
// (12, 8, 'lutff_7/in_1')
// (12, 8, 'sp4_h_r_6')
// (12, 8, 'sp4_v_t_36')
// (12, 9, 'sp4_r_v_b_37')
// (12, 9, 'sp4_v_b_36')
// (12, 10, 'neigh_op_top_6')
// (12, 10, 'sp4_r_v_b_24')
// (12, 10, 'sp4_v_b_25')
// (12, 11, 'lutff_6/out')
// (12, 11, 'sp4_r_v_b_13')
// (12, 11, 'sp4_r_v_b_45')
// (12, 11, 'sp4_v_b_12')
// (12, 12, 'neigh_op_bot_6')
// (12, 12, 'sp4_r_v_b_0')
// (12, 12, 'sp4_r_v_b_32')
// (12, 12, 'sp4_v_b_1')
// (12, 13, 'sp4_r_v_b_21')
// (12, 14, 'sp4_r_v_b_8')
// (13, 8, 'sp4_h_r_19')
// (13, 8, 'sp4_v_t_37')
// (13, 9, 'local_g3_5')
// (13, 9, 'lutff_1/in_1')
// (13, 9, 'sp4_v_b_37')
// (13, 10, 'neigh_op_tnl_6')
// (13, 10, 'sp4_v_b_24')
// (13, 10, 'sp4_v_t_45')
// (13, 11, 'local_g0_6')
// (13, 11, 'lutff_1/in_1')
// (13, 11, 'neigh_op_lft_6')
// (13, 11, 'sp4_v_b_13')
// (13, 11, 'sp4_v_b_45')
// (13, 12, 'neigh_op_bnl_6')
// (13, 12, 'sp4_v_b_0')
// (13, 12, 'sp4_v_b_32')
// (13, 13, 'sp4_v_b_21')
// (13, 14, 'local_g1_0')
// (13, 14, 'lutff_3/in_0')
// (13, 14, 'sp4_v_b_8')
// (14, 8, 'sp4_h_r_30')
// (15, 8, 'sp4_h_r_43')
// (16, 8, 'sp4_h_l_43')

reg n1599 = 0;
// (11, 9, 'sp4_r_v_b_47')
// (11, 10, 'local_g0_1')
// (11, 10, 'lutff_1/in_2')
// (11, 10, 'sp4_r_v_b_34')
// (11, 11, 'neigh_op_tnr_5')
// (11, 11, 'sp4_r_v_b_23')
// (11, 12, 'neigh_op_rgt_5')
// (11, 12, 'sp4_r_v_b_10')
// (11, 12, 'sp4_r_v_b_42')
// (11, 13, 'local_g0_5')
// (11, 13, 'lutff_5/in_2')
// (11, 13, 'neigh_op_bnr_5')
// (11, 13, 'sp4_r_v_b_31')
// (11, 13, 'sp4_r_v_b_41')
// (11, 14, 'local_g3_2')
// (11, 14, 'lutff_6/in_1')
// (11, 14, 'sp4_r_v_b_18')
// (11, 14, 'sp4_r_v_b_28')
// (11, 15, 'local_g3_1')
// (11, 15, 'lutff_5/in_3')
// (11, 15, 'lutff_7/in_3')
// (11, 15, 'sp4_r_v_b_17')
// (11, 15, 'sp4_r_v_b_7')
// (11, 16, 'sp4_r_v_b_4')
// (12, 8, 'sp4_v_t_47')
// (12, 9, 'sp4_v_b_47')
// (12, 10, 'sp4_v_b_34')
// (12, 11, 'neigh_op_top_5')
// (12, 11, 'sp4_v_b_23')
// (12, 11, 'sp4_v_t_42')
// (12, 12, 'lutff_5/out')
// (12, 12, 'sp4_h_r_10')
// (12, 12, 'sp4_v_b_10')
// (12, 12, 'sp4_v_b_42')
// (12, 12, 'sp4_v_t_41')
// (12, 13, 'neigh_op_bot_5')
// (12, 13, 'sp4_v_b_31')
// (12, 13, 'sp4_v_b_41')
// (12, 14, 'sp4_v_b_18')
// (12, 14, 'sp4_v_b_28')
// (12, 15, 'sp4_v_b_17')
// (12, 15, 'sp4_v_b_7')
// (12, 16, 'sp4_v_b_4')
// (13, 11, 'neigh_op_tnl_5')
// (13, 12, 'neigh_op_lft_5')
// (13, 12, 'sp4_h_r_23')
// (13, 13, 'neigh_op_bnl_5')
// (14, 12, 'sp4_h_r_34')
// (15, 12, 'sp4_h_r_47')
// (16, 12, 'sp4_h_l_47')

wire n1600;
// (11, 10, 'neigh_op_tnr_7')
// (11, 11, 'neigh_op_rgt_7')
// (11, 12, 'neigh_op_bnr_7')
// (12, 10, 'neigh_op_top_7')
// (12, 11, 'lutff_7/out')
// (12, 12, 'local_g1_7')
// (12, 12, 'lutff_2/in_2')
// (12, 12, 'neigh_op_bot_7')
// (13, 10, 'neigh_op_tnl_7')
// (13, 11, 'neigh_op_lft_7')
// (13, 12, 'neigh_op_bnl_7')

wire n1601;
// (11, 11, 'local_g3_3')
// (11, 11, 'lutff_4/in_0')
// (11, 11, 'neigh_op_tnr_3')
// (11, 12, 'neigh_op_rgt_3')
// (11, 13, 'neigh_op_bnr_3')
// (12, 11, 'neigh_op_top_3')
// (12, 12, 'lutff_3/out')
// (12, 13, 'neigh_op_bot_3')
// (13, 11, 'neigh_op_tnl_3')
// (13, 12, 'neigh_op_lft_3')
// (13, 13, 'neigh_op_bnl_3')

wire n1602;
// (11, 11, 'lutff_1/cout')
// (11, 11, 'lutff_2/in_3')

wire n1603;
// (11, 11, 'lutff_3/cout')
// (11, 11, 'lutff_4/in_3')

wire n1604;
// (11, 11, 'neigh_op_tnr_1')
// (11, 12, 'neigh_op_rgt_1')
// (11, 13, 'neigh_op_bnr_1')
// (12, 11, 'neigh_op_top_1')
// (12, 12, 'lutff_1/out')
// (12, 13, 'local_g0_1')
// (12, 13, 'lutff_0/in_1')
// (12, 13, 'neigh_op_bot_1')
// (13, 11, 'neigh_op_tnl_1')
// (13, 12, 'neigh_op_lft_1')
// (13, 13, 'neigh_op_bnl_1')

wire n1605;
// (11, 11, 'neigh_op_tnr_2')
// (11, 12, 'neigh_op_rgt_2')
// (11, 12, 'sp4_r_v_b_36')
// (11, 13, 'neigh_op_bnr_2')
// (11, 13, 'sp4_r_v_b_25')
// (11, 14, 'sp4_r_v_b_12')
// (11, 15, 'sp4_r_v_b_1')
// (12, 11, 'neigh_op_top_2')
// (12, 11, 'sp4_v_t_36')
// (12, 12, 'lutff_2/out')
// (12, 12, 'sp4_v_b_36')
// (12, 13, 'neigh_op_bot_2')
// (12, 13, 'sp4_v_b_25')
// (12, 14, 'local_g1_4')
// (12, 14, 'lutff_4/in_3')
// (12, 14, 'sp4_v_b_12')
// (12, 15, 'sp4_v_b_1')
// (13, 11, 'neigh_op_tnl_2')
// (13, 12, 'neigh_op_lft_2')
// (13, 13, 'neigh_op_bnl_2')

wire n1606;
// (11, 11, 'neigh_op_tnr_4')
// (11, 12, 'neigh_op_rgt_4')
// (11, 13, 'neigh_op_bnr_4')
// (12, 11, 'neigh_op_top_4')
// (12, 12, 'local_g3_4')
// (12, 12, 'lutff_1/in_2')
// (12, 12, 'lutff_4/out')
// (12, 13, 'neigh_op_bot_4')
// (13, 11, 'neigh_op_tnl_4')
// (13, 12, 'neigh_op_lft_4')
// (13, 13, 'neigh_op_bnl_4')

wire n1607;
// (11, 11, 'neigh_op_tnr_6')
// (11, 12, 'neigh_op_rgt_6')
// (11, 13, 'neigh_op_bnr_6')
// (12, 11, 'neigh_op_top_6')
// (12, 12, 'local_g1_6')
// (12, 12, 'lutff_0/in_1')
// (12, 12, 'lutff_6/out')
// (12, 13, 'local_g0_6')
// (12, 13, 'lutff_2/in_0')
// (12, 13, 'neigh_op_bot_6')
// (13, 11, 'neigh_op_tnl_6')
// (13, 12, 'neigh_op_lft_6')
// (13, 13, 'neigh_op_bnl_6')

reg n1608 = 0;
// (11, 11, 'sp4_h_r_6')
// (11, 15, 'sp4_h_r_0')
// (12, 11, 'local_g1_3')
// (12, 11, 'lutff_0/in_0')
// (12, 11, 'lutff_3/in_3')
// (12, 11, 'sp4_h_r_19')
// (12, 15, 'local_g1_5')
// (12, 15, 'lutff_3/in_1')
// (12, 15, 'lutff_5/in_1')
// (12, 15, 'sp4_h_r_13')
// (13, 11, 'sp4_h_r_30')
// (13, 15, 'sp4_h_r_24')
// (14, 11, 'sp4_h_r_43')
// (14, 12, 'sp4_r_v_b_37')
// (14, 12, 'sp4_r_v_b_38')
// (14, 13, 'sp4_r_v_b_24')
// (14, 13, 'sp4_r_v_b_27')
// (14, 14, 'sp4_r_v_b_13')
// (14, 14, 'sp4_r_v_b_14')
// (14, 15, 'local_g1_3')
// (14, 15, 'lutff_3/in_3')
// (14, 15, 'sp4_h_r_37')
// (14, 15, 'sp4_r_v_b_0')
// (14, 15, 'sp4_r_v_b_3')
// (15, 11, 'sp4_h_l_43')
// (15, 11, 'sp4_h_r_3')
// (15, 11, 'sp4_h_r_6')
// (15, 11, 'sp4_v_t_37')
// (15, 11, 'sp4_v_t_38')
// (15, 12, 'sp4_v_b_37')
// (15, 12, 'sp4_v_b_38')
// (15, 13, 'sp4_v_b_24')
// (15, 13, 'sp4_v_b_27')
// (15, 14, 'sp4_v_b_13')
// (15, 14, 'sp4_v_b_14')
// (15, 15, 'local_g1_0')
// (15, 15, 'lutff_7/in_0')
// (15, 15, 'sp4_h_l_37')
// (15, 15, 'sp4_v_b_0')
// (15, 15, 'sp4_v_b_3')
// (16, 11, 'sp4_h_r_14')
// (16, 11, 'sp4_h_r_19')
// (17, 11, 'sp4_h_r_27')
// (17, 11, 'sp4_h_r_30')
// (18, 11, 'sp4_h_r_38')
// (18, 11, 'sp4_h_r_43')
// (19, 11, 'sp4_h_l_38')
// (19, 11, 'sp4_h_l_43')
// (19, 11, 'sp4_h_r_3')
// (20, 11, 'sp4_h_r_14')
// (21, 10, 'neigh_op_tnr_3')
// (21, 11, 'neigh_op_rgt_3')
// (21, 11, 'sp4_h_r_27')
// (21, 12, 'neigh_op_bnr_3')
// (22, 10, 'neigh_op_top_3')
// (22, 11, 'lutff_3/out')
// (22, 11, 'sp4_h_r_38')
// (22, 12, 'neigh_op_bot_3')
// (23, 10, 'neigh_op_tnl_3')
// (23, 11, 'neigh_op_lft_3')
// (23, 11, 'sp4_h_l_38')
// (23, 12, 'neigh_op_bnl_3')

reg n1609 = 0;
// (11, 11, 'sp4_r_v_b_36')
// (11, 12, 'sp4_r_v_b_25')
// (11, 13, 'sp4_r_v_b_12')
// (11, 14, 'sp4_r_v_b_1')
// (11, 15, 'sp4_r_v_b_36')
// (11, 16, 'neigh_op_tnr_6')
// (11, 16, 'sp4_r_v_b_25')
// (11, 16, 'sp4_r_v_b_41')
// (11, 17, 'neigh_op_rgt_6')
// (11, 17, 'sp4_r_v_b_12')
// (11, 17, 'sp4_r_v_b_28')
// (11, 18, 'neigh_op_bnr_6')
// (11, 18, 'sp4_r_v_b_1')
// (11, 18, 'sp4_r_v_b_17')
// (11, 19, 'sp4_r_v_b_4')
// (12, 10, 'sp4_v_t_36')
// (12, 11, 'local_g3_4')
// (12, 11, 'lutff_0/in_3')
// (12, 11, 'lutff_3/in_2')
// (12, 11, 'sp4_v_b_36')
// (12, 12, 'sp4_v_b_25')
// (12, 13, 'sp4_v_b_12')
// (12, 14, 'sp4_v_b_1')
// (12, 14, 'sp4_v_t_36')
// (12, 15, 'local_g3_4')
// (12, 15, 'lutff_5/in_0')
// (12, 15, 'sp4_h_r_9')
// (12, 15, 'sp4_v_b_36')
// (12, 15, 'sp4_v_t_41')
// (12, 16, 'neigh_op_top_6')
// (12, 16, 'sp4_v_b_25')
// (12, 16, 'sp4_v_b_41')
// (12, 17, 'lutff_6/out')
// (12, 17, 'sp4_v_b_12')
// (12, 17, 'sp4_v_b_28')
// (12, 18, 'local_g1_6')
// (12, 18, 'lutff_1/in_2')
// (12, 18, 'neigh_op_bot_6')
// (12, 18, 'sp4_v_b_1')
// (12, 18, 'sp4_v_b_17')
// (12, 19, 'sp4_v_b_4')
// (13, 15, 'sp4_h_r_20')
// (13, 16, 'neigh_op_tnl_6')
// (13, 17, 'neigh_op_lft_6')
// (13, 18, 'neigh_op_bnl_6')
// (14, 15, 'local_g2_1')
// (14, 15, 'lutff_3/in_0')
// (14, 15, 'sp4_h_r_33')
// (15, 15, 'sp4_h_r_44')
// (16, 15, 'sp4_h_l_44')

wire n1610;
// (11, 12, 'neigh_op_tnr_0')
// (11, 13, 'neigh_op_rgt_0')
// (11, 14, 'neigh_op_bnr_0')
// (12, 12, 'neigh_op_top_0')
// (12, 13, 'lutff_0/out')
// (12, 14, 'local_g1_0')
// (12, 14, 'lutff_7/in_0')
// (12, 14, 'neigh_op_bot_0')
// (13, 12, 'neigh_op_tnl_0')
// (13, 13, 'neigh_op_lft_0')
// (13, 14, 'neigh_op_bnl_0')

reg n1611 = 0;
// (11, 12, 'neigh_op_tnr_1')
// (11, 13, 'neigh_op_rgt_1')
// (11, 14, 'local_g0_1')
// (11, 14, 'lutff_1/in_0')
// (11, 14, 'neigh_op_bnr_1')
// (12, 12, 'neigh_op_top_1')
// (12, 13, 'lutff_1/out')
// (12, 14, 'neigh_op_bot_1')
// (13, 12, 'neigh_op_tnl_1')
// (13, 13, 'neigh_op_lft_1')
// (13, 14, 'neigh_op_bnl_1')

wire n1612;
// (11, 12, 'neigh_op_tnr_2')
// (11, 13, 'neigh_op_rgt_2')
// (11, 14, 'neigh_op_bnr_2')
// (12, 12, 'neigh_op_top_2')
// (12, 13, 'local_g2_2')
// (12, 13, 'lutff_0/in_0')
// (12, 13, 'lutff_2/out')
// (12, 14, 'neigh_op_bot_2')
// (13, 12, 'neigh_op_tnl_2')
// (13, 13, 'neigh_op_lft_2')
// (13, 14, 'neigh_op_bnl_2')

reg n1613 = 0;
// (11, 12, 'neigh_op_tnr_5')
// (11, 13, 'neigh_op_rgt_5')
// (11, 14, 'neigh_op_bnr_5')
// (12, 12, 'neigh_op_top_5')
// (12, 12, 'sp4_r_v_b_38')
// (12, 13, 'lutff_5/out')
// (12, 13, 'sp4_r_v_b_27')
// (12, 14, 'neigh_op_bot_5')
// (12, 14, 'sp4_r_v_b_14')
// (12, 15, 'local_g1_3')
// (12, 15, 'lutff_6/in_0')
// (12, 15, 'sp4_r_v_b_3')
// (13, 11, 'sp4_v_t_38')
// (13, 12, 'neigh_op_tnl_5')
// (13, 12, 'sp4_v_b_38')
// (13, 13, 'neigh_op_lft_5')
// (13, 13, 'sp4_v_b_27')
// (13, 14, 'neigh_op_bnl_5')
// (13, 14, 'sp4_v_b_14')
// (13, 15, 'sp4_v_b_3')

reg n1614 = 0;
// (11, 12, 'neigh_op_tnr_7')
// (11, 13, 'neigh_op_rgt_7')
// (11, 14, 'local_g1_7')
// (11, 14, 'lutff_4/in_2')
// (11, 14, 'neigh_op_bnr_7')
// (12, 12, 'neigh_op_top_7')
// (12, 13, 'lutff_7/out')
// (12, 14, 'neigh_op_bot_7')
// (13, 12, 'neigh_op_tnl_7')
// (13, 13, 'neigh_op_lft_7')
// (13, 14, 'neigh_op_bnl_7')

wire n1615;
// (11, 12, 'sp4_r_v_b_37')
// (11, 13, 'sp4_r_v_b_24')
// (11, 14, 'sp4_r_v_b_13')
// (11, 15, 'sp4_r_v_b_0')
// (12, 11, 'sp4_v_t_37')
// (12, 12, 'sp4_v_b_37')
// (12, 13, 'local_g3_0')
// (12, 13, 'lutff_6/in_3')
// (12, 13, 'sp4_v_b_24')
// (12, 14, 'sp4_v_b_13')
// (12, 15, 'sp4_h_r_7')
// (12, 15, 'sp4_v_b_0')
// (13, 15, 'sp4_h_r_18')
// (14, 15, 'sp4_h_r_31')
// (15, 15, 'sp4_h_r_42')
// (16, 15, 'sp4_h_l_42')
// (16, 15, 'sp4_h_r_11')
// (17, 15, 'sp4_h_r_22')
// (18, 14, 'neigh_op_tnr_7')
// (18, 15, 'neigh_op_rgt_7')
// (18, 15, 'sp4_h_r_35')
// (18, 16, 'neigh_op_bnr_7')
// (19, 14, 'neigh_op_top_7')
// (19, 15, 'ram/RDATA_8')
// (19, 15, 'sp4_h_r_46')
// (19, 16, 'neigh_op_bot_7')
// (20, 14, 'neigh_op_tnl_7')
// (20, 15, 'neigh_op_lft_7')
// (20, 15, 'sp4_h_l_46')
// (20, 16, 'neigh_op_bnl_7')

wire n1616;
// (11, 12, 'sp4_r_v_b_46')
// (11, 13, 'sp4_r_v_b_35')
// (11, 14, 'sp4_r_v_b_22')
// (11, 15, 'sp4_r_v_b_11')
// (12, 11, 'sp4_v_t_46')
// (12, 12, 'sp4_v_b_46')
// (12, 13, 'local_g2_3')
// (12, 13, 'lutff_4/in_1')
// (12, 13, 'sp4_v_b_35')
// (12, 14, 'sp4_v_b_22')
// (12, 15, 'sp4_h_r_11')
// (12, 15, 'sp4_v_b_11')
// (13, 15, 'sp4_h_r_22')
// (14, 15, 'sp4_h_r_35')
// (15, 15, 'sp4_h_r_46')
// (16, 15, 'sp4_h_l_46')
// (16, 15, 'sp4_h_r_3')
// (17, 15, 'sp4_h_r_14')
// (18, 14, 'neigh_op_tnr_3')
// (18, 15, 'neigh_op_rgt_3')
// (18, 15, 'sp4_h_r_27')
// (18, 16, 'neigh_op_bnr_3')
// (19, 14, 'neigh_op_top_3')
// (19, 15, 'ram/RDATA_12')
// (19, 15, 'sp4_h_r_38')
// (19, 16, 'neigh_op_bot_3')
// (20, 14, 'neigh_op_tnl_3')
// (20, 15, 'neigh_op_lft_3')
// (20, 15, 'sp4_h_l_38')
// (20, 16, 'neigh_op_bnl_3')

reg n1617 = 0;
// (11, 13, 'neigh_op_tnr_1')
// (11, 14, 'neigh_op_rgt_1')
// (11, 15, 'neigh_op_bnr_1')
// (12, 13, 'local_g1_1')
// (12, 13, 'lutff_0/in_2')
// (12, 13, 'neigh_op_top_1')
// (12, 14, 'local_g2_1')
// (12, 14, 'lutff_1/in_2')
// (12, 14, 'lutff_1/out')
// (12, 14, 'sp4_h_r_2')
// (12, 15, 'neigh_op_bot_1')
// (13, 13, 'neigh_op_tnl_1')
// (13, 14, 'neigh_op_lft_1')
// (13, 14, 'sp4_h_r_15')
// (13, 15, 'neigh_op_bnl_1')
// (14, 14, 'sp4_h_r_26')
// (15, 11, 'sp4_r_v_b_39')
// (15, 12, 'sp4_r_v_b_26')
// (15, 13, 'sp4_r_v_b_15')
// (15, 14, 'sp4_h_r_39')
// (15, 14, 'sp4_r_v_b_2')
// (16, 10, 'sp4_h_r_2')
// (16, 10, 'sp4_v_t_39')
// (16, 11, 'sp4_v_b_39')
// (16, 12, 'sp4_v_b_26')
// (16, 13, 'sp4_v_b_15')
// (16, 14, 'sp4_h_l_39')
// (16, 14, 'sp4_v_b_2')
// (17, 10, 'local_g0_7')
// (17, 10, 'lutff_1/in_2')
// (17, 10, 'sp4_h_r_15')
// (18, 10, 'sp4_h_r_26')
// (19, 10, 'sp4_h_r_39')
// (20, 10, 'sp4_h_l_39')

reg n1618 = 0;
// (11, 13, 'neigh_op_tnr_2')
// (11, 14, 'neigh_op_rgt_2')
// (11, 15, 'neigh_op_bnr_2')
// (12, 11, 'sp4_r_v_b_40')
// (12, 12, 'sp4_r_v_b_29')
// (12, 13, 'neigh_op_top_2')
// (12, 13, 'sp4_r_v_b_16')
// (12, 14, 'local_g2_2')
// (12, 14, 'lutff_2/in_2')
// (12, 14, 'lutff_2/out')
// (12, 14, 'lutff_4/in_0')
// (12, 14, 'sp4_r_v_b_5')
// (12, 15, 'neigh_op_bot_2')
// (13, 10, 'sp4_h_r_10')
// (13, 10, 'sp4_v_t_40')
// (13, 11, 'sp4_v_b_40')
// (13, 12, 'sp4_v_b_29')
// (13, 13, 'neigh_op_tnl_2')
// (13, 13, 'sp4_v_b_16')
// (13, 14, 'neigh_op_lft_2')
// (13, 14, 'sp4_v_b_5')
// (13, 15, 'neigh_op_bnl_2')
// (14, 10, 'sp4_h_r_23')
// (15, 10, 'sp4_h_r_34')
// (16, 10, 'sp4_h_r_47')
// (17, 10, 'local_g1_2')
// (17, 10, 'lutff_2/in_1')
// (17, 10, 'sp4_h_l_47')
// (17, 10, 'sp4_h_r_10')
// (18, 10, 'sp4_h_r_23')
// (19, 10, 'sp4_h_r_34')
// (20, 10, 'sp4_h_r_47')
// (21, 10, 'sp4_h_l_47')

reg n1619 = 0;
// (11, 13, 'neigh_op_tnr_3')
// (11, 14, 'neigh_op_rgt_3')
// (11, 15, 'neigh_op_bnr_3')
// (12, 13, 'neigh_op_top_3')
// (12, 14, 'local_g0_3')
// (12, 14, 'lutff_3/in_2')
// (12, 14, 'lutff_3/out')
// (12, 14, 'lutff_4/in_1')
// (12, 15, 'neigh_op_bot_3')
// (13, 13, 'neigh_op_tnl_3')
// (13, 14, 'neigh_op_lft_3')
// (13, 15, 'neigh_op_bnl_3')

wire n1620;
// (11, 13, 'neigh_op_tnr_4')
// (11, 14, 'neigh_op_rgt_4')
// (11, 15, 'neigh_op_bnr_4')
// (12, 13, 'neigh_op_top_4')
// (12, 14, 'local_g2_4')
// (12, 14, 'lutff_4/out')
// (12, 14, 'lutff_7/in_1')
// (12, 15, 'neigh_op_bot_4')
// (13, 13, 'neigh_op_tnl_4')
// (13, 14, 'neigh_op_lft_4')
// (13, 15, 'neigh_op_bnl_4')

wire n1621;
// (11, 13, 'neigh_op_tnr_5')
// (11, 14, 'neigh_op_rgt_5')
// (11, 15, 'neigh_op_bnr_5')
// (12, 13, 'neigh_op_top_5')
// (12, 13, 'sp4_r_v_b_38')
// (12, 14, 'lutff_5/out')
// (12, 14, 'sp4_r_v_b_27')
// (12, 15, 'neigh_op_bot_5')
// (12, 15, 'sp4_r_v_b_14')
// (12, 16, 'sp4_r_v_b_3')
// (13, 12, 'sp4_v_t_38')
// (13, 13, 'neigh_op_tnl_5')
// (13, 13, 'sp4_v_b_38')
// (13, 14, 'neigh_op_lft_5')
// (13, 14, 'sp4_v_b_27')
// (13, 15, 'neigh_op_bnl_5')
// (13, 15, 'sp4_v_b_14')
// (13, 16, 'sp4_h_r_9')
// (13, 16, 'sp4_v_b_3')
// (14, 16, 'local_g0_4')
// (14, 16, 'lutff_6/in_2')
// (14, 16, 'sp4_h_r_20')
// (15, 16, 'sp4_h_r_33')
// (16, 16, 'sp4_h_r_44')
// (17, 16, 'sp4_h_l_44')

reg n1622 = 0;
// (11, 13, 'neigh_op_tnr_6')
// (11, 14, 'neigh_op_rgt_6')
// (11, 15, 'neigh_op_bnr_6')
// (12, 12, 'sp4_r_v_b_37')
// (12, 13, 'local_g1_6')
// (12, 13, 'lutff_0/in_3')
// (12, 13, 'neigh_op_top_6')
// (12, 13, 'sp4_r_v_b_24')
// (12, 14, 'local_g0_6')
// (12, 14, 'local_g3_6')
// (12, 14, 'lutff_0/in_1')
// (12, 14, 'lutff_1/in_3')
// (12, 14, 'lutff_6/in_3')
// (12, 14, 'lutff_6/out')
// (12, 14, 'sp4_r_v_b_13')
// (12, 15, 'neigh_op_bot_6')
// (12, 15, 'sp4_r_v_b_0')
// (13, 11, 'sp4_h_r_0')
// (13, 11, 'sp4_v_t_37')
// (13, 12, 'sp4_v_b_37')
// (13, 13, 'neigh_op_tnl_6')
// (13, 13, 'sp4_v_b_24')
// (13, 14, 'neigh_op_lft_6')
// (13, 14, 'sp4_v_b_13')
// (13, 15, 'neigh_op_bnl_6')
// (13, 15, 'sp4_v_b_0')
// (14, 11, 'sp4_h_r_13')
// (15, 11, 'sp4_h_r_24')
// (16, 8, 'sp4_r_v_b_37')
// (16, 9, 'sp4_r_v_b_24')
// (16, 10, 'sp4_r_v_b_13')
// (16, 11, 'sp4_h_r_37')
// (16, 11, 'sp4_r_v_b_0')
// (17, 7, 'sp4_v_t_37')
// (17, 8, 'sp4_v_b_37')
// (17, 9, 'sp4_v_b_24')
// (17, 10, 'local_g1_5')
// (17, 10, 'lutff_0/in_2')
// (17, 10, 'lutff_6/in_2')
// (17, 10, 'sp4_v_b_13')
// (17, 11, 'sp4_h_l_37')
// (17, 11, 'sp4_v_b_0')

wire n1623;
// (11, 13, 'neigh_op_tnr_7')
// (11, 14, 'neigh_op_rgt_7')
// (11, 15, 'local_g1_7')
// (11, 15, 'lutff_4/in_0')
// (11, 15, 'neigh_op_bnr_7')
// (12, 13, 'neigh_op_top_7')
// (12, 13, 'sp4_r_v_b_42')
// (12, 14, 'local_g0_7')
// (12, 14, 'local_g1_7')
// (12, 14, 'lutff_1/in_0')
// (12, 14, 'lutff_2/in_0')
// (12, 14, 'lutff_3/in_0')
// (12, 14, 'lutff_6/in_1')
// (12, 14, 'lutff_7/out')
// (12, 14, 'sp4_r_v_b_31')
// (12, 15, 'local_g1_7')
// (12, 15, 'lutff_4/in_0')
// (12, 15, 'neigh_op_bot_7')
// (12, 15, 'sp4_r_v_b_18')
// (12, 16, 'sp4_r_v_b_7')
// (13, 12, 'sp4_v_t_42')
// (13, 13, 'neigh_op_tnl_7')
// (13, 13, 'sp4_v_b_42')
// (13, 14, 'neigh_op_lft_7')
// (13, 14, 'sp4_v_b_31')
// (13, 15, 'neigh_op_bnl_7')
// (13, 15, 'sp4_v_b_18')
// (13, 16, 'sp4_h_r_1')
// (13, 16, 'sp4_v_b_7')
// (14, 16, 'sp4_h_r_12')
// (15, 16, 'local_g3_1')
// (15, 16, 'lutff_2/in_0')
// (15, 16, 'lutff_4/in_0')
// (15, 16, 'lutff_6/in_2')
// (15, 16, 'lutff_7/in_1')
// (15, 16, 'sp4_h_r_25')
// (16, 16, 'sp4_h_r_36')
// (17, 16, 'sp4_h_l_36')

reg n1624 = 0;
// (11, 13, 'sp4_h_r_3')
// (11, 14, 'sp4_h_r_6')
// (12, 13, 'sp4_h_r_14')
// (12, 14, 'sp4_h_r_19')
// (13, 13, 'local_g3_3')
// (13, 13, 'lutff_0/in_0')
// (13, 13, 'lutff_2/in_2')
// (13, 13, 'sp4_h_r_27')
// (13, 14, 'local_g3_6')
// (13, 14, 'lutff_2/in_1')
// (13, 14, 'sp4_h_r_30')
// (14, 13, 'sp4_h_r_38')
// (14, 14, 'sp4_h_r_43')
// (14, 14, 'sp4_r_v_b_38')
// (14, 15, 'neigh_op_tnr_7')
// (14, 15, 'sp4_r_v_b_27')
// (14, 15, 'sp4_r_v_b_43')
// (14, 16, 'neigh_op_rgt_7')
// (14, 16, 'sp4_r_v_b_14')
// (14, 16, 'sp4_r_v_b_30')
// (14, 17, 'neigh_op_bnr_7')
// (14, 17, 'sp4_r_v_b_19')
// (14, 17, 'sp4_r_v_b_3')
// (14, 18, 'sp4_r_v_b_6')
// (15, 11, 'sp4_r_v_b_42')
// (15, 12, 'sp4_r_v_b_31')
// (15, 13, 'local_g0_3')
// (15, 13, 'lutff_3/in_2')
// (15, 13, 'sp4_h_l_38')
// (15, 13, 'sp4_h_r_3')
// (15, 13, 'sp4_r_v_b_18')
// (15, 13, 'sp4_v_t_38')
// (15, 14, 'local_g3_6')
// (15, 14, 'lutff_3/in_2')
// (15, 14, 'lutff_5/in_0')
// (15, 14, 'sp4_h_l_43')
// (15, 14, 'sp4_r_v_b_39')
// (15, 14, 'sp4_r_v_b_7')
// (15, 14, 'sp4_v_b_38')
// (15, 14, 'sp4_v_t_43')
// (15, 15, 'local_g0_7')
// (15, 15, 'lutff_3/in_2')
// (15, 15, 'lutff_4/in_3')
// (15, 15, 'neigh_op_top_7')
// (15, 15, 'sp4_r_v_b_26')
// (15, 15, 'sp4_r_v_b_42')
// (15, 15, 'sp4_v_b_27')
// (15, 15, 'sp4_v_b_43')
// (15, 16, 'local_g3_7')
// (15, 16, 'lutff_1/in_1')
// (15, 16, 'lutff_5/in_3')
// (15, 16, 'lutff_7/in_3')
// (15, 16, 'lutff_7/out')
// (15, 16, 'sp4_r_v_b_15')
// (15, 16, 'sp4_r_v_b_31')
// (15, 16, 'sp4_v_b_14')
// (15, 16, 'sp4_v_b_30')
// (15, 17, 'neigh_op_bot_7')
// (15, 17, 'sp4_r_v_b_18')
// (15, 17, 'sp4_r_v_b_2')
// (15, 17, 'sp4_v_b_19')
// (15, 17, 'sp4_v_b_3')
// (15, 18, 'sp4_r_v_b_7')
// (15, 18, 'sp4_v_b_6')
// (16, 10, 'sp4_v_t_42')
// (16, 11, 'sp4_v_b_42')
// (16, 12, 'local_g2_7')
// (16, 12, 'lutff_6/in_1')
// (16, 12, 'sp4_v_b_31')
// (16, 13, 'sp4_h_r_14')
// (16, 13, 'sp4_v_b_18')
// (16, 13, 'sp4_v_t_39')
// (16, 14, 'local_g3_7')
// (16, 14, 'lutff_5/in_3')
// (16, 14, 'sp4_v_b_39')
// (16, 14, 'sp4_v_b_7')
// (16, 14, 'sp4_v_t_42')
// (16, 15, 'neigh_op_tnl_7')
// (16, 15, 'sp4_v_b_26')
// (16, 15, 'sp4_v_b_42')
// (16, 16, 'neigh_op_lft_7')
// (16, 16, 'sp4_v_b_15')
// (16, 16, 'sp4_v_b_31')
// (16, 17, 'neigh_op_bnl_7')
// (16, 17, 'sp4_v_b_18')
// (16, 17, 'sp4_v_b_2')
// (16, 18, 'sp4_v_b_7')
// (17, 13, 'sp4_h_r_27')
// (18, 13, 'sp4_h_r_38')
// (19, 13, 'sp4_h_l_38')

wire n1625;
// (11, 13, 'sp4_h_r_7')
// (12, 13, 'local_g1_2')
// (12, 13, 'lutff_1/in_2')
// (12, 13, 'sp4_h_r_18')
// (13, 13, 'sp4_h_r_31')
// (14, 13, 'sp4_h_r_42')
// (15, 13, 'sp4_h_l_42')
// (15, 13, 'sp4_h_r_4')
// (16, 13, 'sp4_h_r_17')
// (17, 13, 'sp4_h_r_28')
// (18, 13, 'sp4_h_r_41')
// (18, 14, 'neigh_op_tnr_1')
// (18, 14, 'sp4_r_v_b_47')
// (18, 15, 'neigh_op_rgt_1')
// (18, 15, 'sp4_r_v_b_34')
// (18, 16, 'neigh_op_bnr_1')
// (18, 16, 'sp4_r_v_b_23')
// (18, 17, 'sp4_r_v_b_10')
// (19, 13, 'sp4_h_l_41')
// (19, 13, 'sp4_v_t_47')
// (19, 14, 'neigh_op_top_1')
// (19, 14, 'sp4_v_b_47')
// (19, 15, 'ram/RDATA_14')
// (19, 15, 'sp4_v_b_34')
// (19, 16, 'neigh_op_bot_1')
// (19, 16, 'sp4_v_b_23')
// (19, 17, 'sp4_v_b_10')
// (20, 14, 'neigh_op_tnl_1')
// (20, 15, 'neigh_op_lft_1')
// (20, 16, 'neigh_op_bnl_1')

wire n1626;
// (11, 13, 'sp4_h_r_8')
// (12, 13, 'local_g0_5')
// (12, 13, 'lutff_7/in_0')
// (12, 13, 'sp4_h_r_21')
// (13, 13, 'sp4_h_r_32')
// (14, 13, 'sp4_h_r_45')
// (15, 13, 'sp4_h_l_45')
// (15, 13, 'sp4_h_r_5')
// (16, 13, 'sp4_h_r_16')
// (17, 13, 'sp4_h_r_29')
// (18, 13, 'sp4_h_r_40')
// (18, 14, 'sp4_r_v_b_46')
// (18, 15, 'neigh_op_tnr_3')
// (18, 15, 'sp4_r_v_b_35')
// (18, 16, 'neigh_op_rgt_3')
// (18, 16, 'sp4_r_v_b_22')
// (18, 17, 'neigh_op_bnr_3')
// (18, 17, 'sp4_r_v_b_11')
// (19, 13, 'sp4_h_l_40')
// (19, 13, 'sp4_v_t_46')
// (19, 14, 'sp4_v_b_46')
// (19, 15, 'neigh_op_top_3')
// (19, 15, 'sp4_v_b_35')
// (19, 16, 'ram/RDATA_4')
// (19, 16, 'sp4_v_b_22')
// (19, 17, 'neigh_op_bot_3')
// (19, 17, 'sp4_v_b_11')
// (20, 15, 'neigh_op_tnl_3')
// (20, 16, 'neigh_op_lft_3')
// (20, 17, 'neigh_op_bnl_3')

wire n1627;
// (11, 13, 'sp4_r_v_b_47')
// (11, 14, 'sp4_r_v_b_34')
// (11, 15, 'sp4_r_v_b_23')
// (11, 16, 'sp4_r_v_b_10')
// (12, 12, 'sp4_v_t_47')
// (12, 13, 'local_g3_7')
// (12, 13, 'lutff_5/in_1')
// (12, 13, 'sp4_v_b_47')
// (12, 14, 'sp4_v_b_34')
// (12, 15, 'sp4_v_b_23')
// (12, 16, 'sp4_h_r_10')
// (12, 16, 'sp4_v_b_10')
// (13, 16, 'sp4_h_r_23')
// (14, 16, 'sp4_h_r_34')
// (15, 16, 'sp4_h_r_47')
// (16, 16, 'sp4_h_l_47')
// (16, 16, 'sp4_h_r_7')
// (17, 16, 'sp4_h_r_18')
// (18, 15, 'neigh_op_tnr_5')
// (18, 16, 'neigh_op_rgt_5')
// (18, 16, 'sp4_h_r_31')
// (18, 17, 'neigh_op_bnr_5')
// (19, 15, 'neigh_op_top_5')
// (19, 16, 'ram/RDATA_2')
// (19, 16, 'sp4_h_r_42')
// (19, 17, 'neigh_op_bot_5')
// (20, 15, 'neigh_op_tnl_5')
// (20, 16, 'neigh_op_lft_5')
// (20, 16, 'sp4_h_l_42')
// (20, 17, 'neigh_op_bnl_5')

reg n1628 = 0;
// (11, 14, 'neigh_op_tnr_0')
// (11, 15, 'neigh_op_rgt_0')
// (11, 16, 'neigh_op_bnr_0')
// (12, 14, 'neigh_op_top_0')
// (12, 14, 'sp4_r_v_b_44')
// (12, 15, 'lutff_0/out')
// (12, 15, 'sp4_r_v_b_33')
// (12, 16, 'neigh_op_bot_0')
// (12, 16, 'sp4_r_v_b_20')
// (12, 17, 'sp4_r_v_b_9')
// (13, 13, 'sp4_v_t_44')
// (13, 14, 'neigh_op_tnl_0')
// (13, 14, 'sp4_v_b_44')
// (13, 15, 'neigh_op_lft_0')
// (13, 15, 'sp4_v_b_33')
// (13, 16, 'neigh_op_bnl_0')
// (13, 16, 'sp4_v_b_20')
// (13, 17, 'sp4_h_r_3')
// (13, 17, 'sp4_v_b_9')
// (14, 17, 'sp4_h_r_14')
// (15, 17, 'sp4_h_r_27')
// (16, 14, 'sp4_r_v_b_44')
// (16, 15, 'sp4_r_v_b_33')
// (16, 16, 'sp4_r_v_b_20')
// (16, 17, 'sp4_h_r_38')
// (16, 17, 'sp4_r_v_b_9')
// (17, 13, 'sp4_v_t_44')
// (17, 14, 'sp4_v_b_44')
// (17, 15, 'sp4_v_b_33')
// (17, 16, 'local_g0_4')
// (17, 16, 'lutff_2/in_0')
// (17, 16, 'sp4_v_b_20')
// (17, 17, 'sp4_h_l_38')
// (17, 17, 'sp4_v_b_9')

reg n1629 = 0;
// (11, 14, 'neigh_op_tnr_1')
// (11, 15, 'neigh_op_rgt_1')
// (11, 16, 'neigh_op_bnr_1')
// (12, 14, 'neigh_op_top_1')
// (12, 15, 'lutff_1/out')
// (12, 15, 'sp4_h_r_2')
// (12, 16, 'neigh_op_bot_1')
// (13, 14, 'neigh_op_tnl_1')
// (13, 15, 'neigh_op_lft_1')
// (13, 15, 'sp4_h_r_15')
// (13, 16, 'neigh_op_bnl_1')
// (14, 15, 'sp4_h_r_26')
// (15, 15, 'sp4_h_r_39')
// (16, 15, 'local_g1_5')
// (16, 15, 'lutff_1/in_1')
// (16, 15, 'sp4_h_l_39')
// (16, 15, 'sp4_h_r_5')
// (17, 15, 'sp4_h_r_16')
// (18, 15, 'sp4_h_r_29')
// (19, 15, 'sp4_h_r_40')
// (20, 15, 'sp4_h_l_40')

wire n1630;
// (11, 14, 'neigh_op_tnr_4')
// (11, 15, 'neigh_op_rgt_4')
// (11, 15, 'sp4_r_v_b_40')
// (11, 16, 'neigh_op_bnr_4')
// (11, 16, 'sp4_r_v_b_29')
// (11, 17, 'sp4_r_v_b_16')
// (11, 18, 'sp4_r_v_b_5')
// (12, 14, 'local_g0_2')
// (12, 14, 'lutff_global/cen')
// (12, 14, 'neigh_op_top_4')
// (12, 14, 'sp4_h_r_10')
// (12, 14, 'sp4_v_t_40')
// (12, 15, 'lutff_4/out')
// (12, 15, 'sp4_v_b_40')
// (12, 16, 'neigh_op_bot_4')
// (12, 16, 'sp4_v_b_29')
// (12, 17, 'sp4_v_b_16')
// (12, 18, 'sp4_v_b_5')
// (13, 14, 'neigh_op_tnl_4')
// (13, 14, 'sp4_h_r_23')
// (13, 15, 'neigh_op_lft_4')
// (13, 16, 'neigh_op_bnl_4')
// (14, 14, 'sp4_h_r_34')
// (15, 14, 'sp4_h_r_47')
// (16, 14, 'sp4_h_l_47')

reg n1631 = 0;
// (11, 14, 'neigh_op_tnr_6')
// (11, 15, 'neigh_op_rgt_6')
// (11, 15, 'sp4_h_r_1')
// (11, 16, 'neigh_op_bnr_6')
// (12, 14, 'neigh_op_top_6')
// (12, 15, 'lutff_6/out')
// (12, 15, 'sp4_h_r_12')
// (12, 16, 'neigh_op_bot_6')
// (13, 14, 'neigh_op_tnl_6')
// (13, 15, 'neigh_op_lft_6')
// (13, 15, 'sp4_h_r_25')
// (13, 16, 'neigh_op_bnl_6')
// (14, 15, 'sp4_h_r_36')
// (15, 15, 'sp4_h_l_36')
// (15, 15, 'sp4_h_r_4')
// (16, 15, 'local_g0_1')
// (16, 15, 'lutff_5/in_0')
// (16, 15, 'sp4_h_r_17')
// (17, 15, 'sp4_h_r_28')
// (18, 15, 'sp4_h_r_41')
// (19, 15, 'sp4_h_l_41')

reg n1632 = 0;
// (11, 14, 'sp4_h_r_4')
// (12, 5, 'sp4_r_v_b_38')
// (12, 5, 'sp4_r_v_b_47')
// (12, 6, 'local_g2_2')
// (12, 6, 'lutff_5/in_1')
// (12, 6, 'sp4_r_v_b_27')
// (12, 6, 'sp4_r_v_b_34')
// (12, 7, 'sp4_r_v_b_14')
// (12, 7, 'sp4_r_v_b_23')
// (12, 8, 'sp4_r_v_b_10')
// (12, 8, 'sp4_r_v_b_3')
// (12, 9, 'sp4_r_v_b_42')
// (12, 10, 'sp4_r_v_b_31')
// (12, 11, 'sp4_r_v_b_18')
// (12, 12, 'sp4_r_v_b_7')
// (12, 13, 'neigh_op_tnr_6')
// (12, 13, 'sp4_r_v_b_41')
// (12, 14, 'neigh_op_rgt_6')
// (12, 14, 'sp4_h_r_17')
// (12, 14, 'sp4_r_v_b_28')
// (12, 15, 'neigh_op_bnr_6')
// (12, 15, 'sp4_r_v_b_17')
// (12, 16, 'sp4_r_v_b_4')
// (13, 4, 'sp4_v_t_38')
// (13, 4, 'sp4_v_t_47')
// (13, 5, 'sp4_v_b_38')
// (13, 5, 'sp4_v_b_47')
// (13, 6, 'local_g3_3')
// (13, 6, 'lutff_1/in_3')
// (13, 6, 'sp4_v_b_27')
// (13, 6, 'sp4_v_b_34')
// (13, 7, 'sp4_v_b_14')
// (13, 7, 'sp4_v_b_23')
// (13, 8, 'sp4_v_b_10')
// (13, 8, 'sp4_v_b_3')
// (13, 8, 'sp4_v_t_42')
// (13, 9, 'sp4_v_b_42')
// (13, 10, 'sp4_v_b_31')
// (13, 11, 'sp4_v_b_18')
// (13, 12, 'local_g2_5')
// (13, 12, 'lutff_6/in_1')
// (13, 12, 'sp4_r_v_b_37')
// (13, 12, 'sp4_v_b_7')
// (13, 12, 'sp4_v_t_41')
// (13, 13, 'neigh_op_top_6')
// (13, 13, 'sp4_r_v_b_24')
// (13, 13, 'sp4_r_v_b_40')
// (13, 13, 'sp4_v_b_41')
// (13, 14, 'lutff_6/out')
// (13, 14, 'sp4_h_r_28')
// (13, 14, 'sp4_r_v_b_13')
// (13, 14, 'sp4_r_v_b_29')
// (13, 14, 'sp4_v_b_28')
// (13, 15, 'neigh_op_bot_6')
// (13, 15, 'sp4_r_v_b_0')
// (13, 15, 'sp4_r_v_b_16')
// (13, 15, 'sp4_v_b_17')
// (13, 16, 'sp4_r_v_b_5')
// (13, 16, 'sp4_v_b_4')
// (14, 7, 'sp4_r_v_b_37')
// (14, 8, 'sp4_r_v_b_24')
// (14, 9, 'sp4_r_v_b_13')
// (14, 10, 'sp4_r_v_b_0')
// (14, 11, 'sp4_r_v_b_41')
// (14, 11, 'sp4_v_t_37')
// (14, 12, 'sp4_h_r_10')
// (14, 12, 'sp4_r_v_b_28')
// (14, 12, 'sp4_v_b_37')
// (14, 12, 'sp4_v_t_40')
// (14, 13, 'neigh_op_tnl_6')
// (14, 13, 'sp4_r_v_b_17')
// (14, 13, 'sp4_v_b_24')
// (14, 13, 'sp4_v_b_40')
// (14, 14, 'neigh_op_lft_6')
// (14, 14, 'sp4_h_r_41')
// (14, 14, 'sp4_r_v_b_4')
// (14, 14, 'sp4_v_b_13')
// (14, 14, 'sp4_v_b_29')
// (14, 15, 'neigh_op_bnl_6')
// (14, 15, 'sp4_v_b_0')
// (14, 15, 'sp4_v_b_16')
// (14, 16, 'sp4_v_b_5')
// (15, 6, 'sp4_v_t_37')
// (15, 7, 'sp4_v_b_37')
// (15, 8, 'sp4_v_b_24')
// (15, 9, 'sp4_v_b_13')
// (15, 10, 'local_g1_0')
// (15, 10, 'lutff_2/in_1')
// (15, 10, 'sp4_v_b_0')
// (15, 10, 'sp4_v_t_41')
// (15, 11, 'sp4_v_b_41')
// (15, 12, 'local_g1_7')
// (15, 12, 'lutff_1/in_1')
// (15, 12, 'sp4_h_r_23')
// (15, 12, 'sp4_v_b_28')
// (15, 13, 'sp4_v_b_17')
// (15, 14, 'sp4_h_l_41')
// (15, 14, 'sp4_v_b_4')
// (16, 12, 'sp4_h_r_34')
// (17, 12, 'local_g2_7')
// (17, 12, 'lutff_4/in_3')
// (17, 12, 'sp4_h_r_47')
// (18, 12, 'sp4_h_l_47')

reg n1633 = 0;
// (11, 15, 'neigh_op_tnr_0')
// (11, 16, 'neigh_op_rgt_0')
// (11, 17, 'neigh_op_bnr_0')
// (12, 15, 'local_g1_0')
// (12, 15, 'lutff_7/in_2')
// (12, 15, 'neigh_op_top_0')
// (12, 16, 'lutff_0/out')
// (12, 17, 'neigh_op_bot_0')
// (13, 15, 'neigh_op_tnl_0')
// (13, 16, 'neigh_op_lft_0')
// (13, 17, 'neigh_op_bnl_0')

reg n1634 = 0;
// (11, 15, 'neigh_op_tnr_1')
// (11, 16, 'neigh_op_rgt_1')
// (11, 17, 'neigh_op_bnr_1')
// (12, 15, 'local_g0_1')
// (12, 15, 'lutff_1/in_2')
// (12, 15, 'neigh_op_top_1')
// (12, 16, 'lutff_1/out')
// (12, 17, 'neigh_op_bot_1')
// (13, 15, 'neigh_op_tnl_1')
// (13, 16, 'neigh_op_lft_1')
// (13, 17, 'neigh_op_bnl_1')

reg n1635 = 0;
// (11, 16, 'neigh_op_tnr_0')
// (11, 17, 'neigh_op_rgt_0')
// (11, 18, 'neigh_op_bnr_0')
// (12, 16, 'neigh_op_top_0')
// (12, 17, 'local_g3_0')
// (12, 17, 'lutff_0/out')
// (12, 17, 'lutff_5/in_0')
// (12, 18, 'neigh_op_bot_0')
// (13, 16, 'neigh_op_tnl_0')
// (13, 17, 'neigh_op_lft_0')
// (13, 18, 'neigh_op_bnl_0')

reg n1636 = 0;
// (11, 16, 'neigh_op_tnr_2')
// (11, 17, 'neigh_op_rgt_2')
// (11, 18, 'neigh_op_bnr_2')
// (12, 16, 'neigh_op_top_2')
// (12, 17, 'local_g2_2')
// (12, 17, 'lutff_2/out')
// (12, 17, 'lutff_7/in_3')
// (12, 17, 'sp4_h_r_4')
// (12, 18, 'neigh_op_bot_2')
// (13, 16, 'neigh_op_tnl_2')
// (13, 17, 'neigh_op_lft_2')
// (13, 17, 'sp4_h_r_17')
// (13, 18, 'neigh_op_bnl_2')
// (14, 17, 'local_g2_4')
// (14, 17, 'lutff_3/in_3')
// (14, 17, 'lutff_6/in_2')
// (14, 17, 'sp4_h_r_28')
// (15, 17, 'sp4_h_r_41')
// (16, 17, 'sp4_h_l_41')

reg n1637 = 0;
// (11, 16, 'neigh_op_tnr_5')
// (11, 17, 'neigh_op_rgt_5')
// (11, 18, 'neigh_op_bnr_5')
// (12, 10, 'sp4_r_v_b_42')
// (12, 11, 'local_g1_7')
// (12, 11, 'lutff_0/in_2')
// (12, 11, 'lutff_3/in_1')
// (12, 11, 'sp4_r_v_b_31')
// (12, 12, 'sp4_r_v_b_18')
// (12, 13, 'sp4_r_v_b_7')
// (12, 14, 'sp4_r_v_b_46')
// (12, 15, 'local_g2_3')
// (12, 15, 'lutff_5/in_2')
// (12, 15, 'sp4_r_v_b_35')
// (12, 16, 'neigh_op_top_5')
// (12, 16, 'sp4_r_v_b_22')
// (12, 16, 'sp4_r_v_b_38')
// (12, 17, 'local_g1_5')
// (12, 17, 'lutff_5/out')
// (12, 17, 'lutff_6/in_0')
// (12, 17, 'sp4_r_v_b_11')
// (12, 17, 'sp4_r_v_b_27')
// (12, 18, 'neigh_op_bot_5')
// (12, 18, 'sp4_r_v_b_14')
// (12, 19, 'sp4_r_v_b_3')
// (13, 9, 'sp4_v_t_42')
// (13, 10, 'sp4_v_b_42')
// (13, 11, 'sp4_v_b_31')
// (13, 12, 'sp4_v_b_18')
// (13, 13, 'sp4_v_b_7')
// (13, 13, 'sp4_v_t_46')
// (13, 14, 'sp4_v_b_46')
// (13, 15, 'sp4_h_r_8')
// (13, 15, 'sp4_v_b_35')
// (13, 15, 'sp4_v_t_38')
// (13, 16, 'neigh_op_tnl_5')
// (13, 16, 'sp4_v_b_22')
// (13, 16, 'sp4_v_b_38')
// (13, 17, 'neigh_op_lft_5')
// (13, 17, 'sp4_v_b_11')
// (13, 17, 'sp4_v_b_27')
// (13, 18, 'neigh_op_bnl_5')
// (13, 18, 'sp4_v_b_14')
// (13, 19, 'sp4_v_b_3')
// (14, 15, 'local_g1_5')
// (14, 15, 'lutff_3/in_1')
// (14, 15, 'sp4_h_r_21')
// (15, 15, 'sp4_h_r_32')
// (16, 15, 'sp4_h_r_45')
// (17, 15, 'sp4_h_l_45')

wire n1638;
// (11, 16, 'neigh_op_tnr_7')
// (11, 17, 'neigh_op_rgt_7')
// (11, 18, 'neigh_op_bnr_7')
// (12, 16, 'neigh_op_top_7')
// (12, 17, 'local_g3_7')
// (12, 17, 'lutff_2/in_2')
// (12, 17, 'lutff_7/out')
// (12, 18, 'neigh_op_bot_7')
// (13, 16, 'neigh_op_tnl_7')
// (13, 17, 'neigh_op_lft_7')
// (13, 18, 'neigh_op_bnl_7')

wire n1639;
// (11, 17, 'local_g3_7')
// (11, 17, 'lutff_6/in_2')
// (11, 17, 'neigh_op_tnr_7')
// (11, 18, 'neigh_op_rgt_7')
// (11, 19, 'neigh_op_bnr_7')
// (12, 17, 'neigh_op_top_7')
// (12, 18, 'local_g1_7')
// (12, 18, 'lutff_2/in_0')
// (12, 18, 'lutff_7/out')
// (12, 19, 'local_g1_7')
// (12, 19, 'lutff_0/in_0')
// (12, 19, 'neigh_op_bot_7')
// (13, 17, 'neigh_op_tnl_7')
// (13, 18, 'neigh_op_lft_7')
// (13, 19, 'neigh_op_bnl_7')

reg n1640 = 0;
// (11, 17, 'neigh_op_tnr_0')
// (11, 18, 'neigh_op_rgt_0')
// (11, 19, 'neigh_op_bnr_0')
// (12, 17, 'neigh_op_top_0')
// (12, 18, 'local_g2_0')
// (12, 18, 'lutff_0/out')
// (12, 18, 'lutff_3/in_1')
// (12, 18, 'lutff_6/in_0')
// (12, 19, 'neigh_op_bot_0')
// (13, 17, 'neigh_op_tnl_0')
// (13, 18, 'neigh_op_lft_0')
// (13, 19, 'neigh_op_bnl_0')

reg n1641 = 0;
// (11, 17, 'neigh_op_tnr_1')
// (11, 18, 'neigh_op_rgt_1')
// (11, 19, 'neigh_op_bnr_1')
// (12, 17, 'neigh_op_top_1')
// (12, 18, 'local_g2_1')
// (12, 18, 'lutff_0/in_1')
// (12, 18, 'lutff_1/out')
// (12, 19, 'neigh_op_bot_1')
// (13, 17, 'neigh_op_tnl_1')
// (13, 18, 'neigh_op_lft_1')
// (13, 19, 'neigh_op_bnl_1')

reg n1642 = 0;
// (11, 17, 'neigh_op_tnr_3')
// (11, 18, 'neigh_op_rgt_3')
// (11, 19, 'neigh_op_bnr_3')
// (12, 17, 'neigh_op_top_3')
// (12, 18, 'local_g0_3')
// (12, 18, 'lutff_3/out')
// (12, 18, 'lutff_5/in_2')
// (12, 18, 'lutff_6/in_3')
// (12, 19, 'neigh_op_bot_3')
// (13, 17, 'neigh_op_tnl_3')
// (13, 18, 'neigh_op_lft_3')
// (13, 19, 'neigh_op_bnl_3')

reg n1643 = 0;
// (11, 17, 'neigh_op_tnr_4')
// (11, 18, 'neigh_op_rgt_4')
// (11, 19, 'neigh_op_bnr_4')
// (12, 17, 'local_g0_4')
// (12, 17, 'lutff_0/in_0')
// (12, 17, 'neigh_op_top_4')
// (12, 18, 'lutff_4/out')
// (12, 19, 'neigh_op_bot_4')
// (13, 17, 'neigh_op_tnl_4')
// (13, 18, 'neigh_op_lft_4')
// (13, 19, 'neigh_op_bnl_4')

reg n1644 = 0;
// (11, 17, 'neigh_op_tnr_5')
// (11, 18, 'neigh_op_rgt_5')
// (11, 19, 'neigh_op_bnr_5')
// (12, 17, 'neigh_op_top_5')
// (12, 18, 'local_g2_5')
// (12, 18, 'lutff_4/in_1')
// (12, 18, 'lutff_5/out')
// (12, 19, 'neigh_op_bot_5')
// (13, 17, 'neigh_op_tnl_5')
// (13, 18, 'neigh_op_lft_5')
// (13, 19, 'neigh_op_bnl_5')

reg n1645 = 0;
// (11, 17, 'sp4_h_r_10')
// (12, 15, 'local_g1_4')
// (12, 15, 'lutff_3/in_2')
// (12, 15, 'sp4_h_r_4')
// (12, 17, 'local_g0_7')
// (12, 17, 'lutff_0/in_3')
// (12, 17, 'sp4_h_r_23')
// (13, 15, 'sp4_h_r_11')
// (13, 15, 'sp4_h_r_17')
// (13, 17, 'sp4_h_r_34')
// (14, 15, 'local_g0_6')
// (14, 15, 'lutff_4/in_0')
// (14, 15, 'sp4_h_r_22')
// (14, 15, 'sp4_h_r_28')
// (14, 17, 'sp4_h_r_47')
// (15, 12, 'sp4_r_v_b_36')
// (15, 13, 'sp4_r_v_b_25')
// (15, 14, 'sp4_r_v_b_12')
// (15, 15, 'local_g1_1')
// (15, 15, 'lutff_7/in_3')
// (15, 15, 'sp4_h_r_35')
// (15, 15, 'sp4_h_r_41')
// (15, 15, 'sp4_r_v_b_1')
// (15, 16, 'neigh_op_tnr_1')
// (15, 16, 'sp4_r_v_b_47')
// (15, 17, 'neigh_op_rgt_1')
// (15, 17, 'sp4_h_l_47')
// (15, 17, 'sp4_h_r_7')
// (15, 17, 'sp4_r_v_b_34')
// (15, 18, 'neigh_op_bnr_1')
// (15, 18, 'sp4_r_v_b_23')
// (15, 19, 'sp4_r_v_b_10')
// (16, 11, 'sp4_v_t_36')
// (16, 12, 'sp4_v_b_36')
// (16, 13, 'sp4_v_b_25')
// (16, 14, 'local_g2_6')
// (16, 14, 'lutff_1/in_3')
// (16, 14, 'sp4_r_v_b_38')
// (16, 14, 'sp4_v_b_12')
// (16, 15, 'sp4_h_l_41')
// (16, 15, 'sp4_h_r_46')
// (16, 15, 'sp4_r_v_b_27')
// (16, 15, 'sp4_v_b_1')
// (16, 15, 'sp4_v_t_47')
// (16, 16, 'neigh_op_top_1')
// (16, 16, 'sp4_r_v_b_14')
// (16, 16, 'sp4_r_v_b_46')
// (16, 16, 'sp4_v_b_47')
// (16, 17, 'local_g0_1')
// (16, 17, 'lutff_1/in_2')
// (16, 17, 'lutff_1/out')
// (16, 17, 'sp4_h_r_18')
// (16, 17, 'sp4_r_v_b_3')
// (16, 17, 'sp4_r_v_b_35')
// (16, 17, 'sp4_v_b_34')
// (16, 18, 'neigh_op_bot_1')
// (16, 18, 'sp4_r_v_b_22')
// (16, 18, 'sp4_v_b_23')
// (16, 19, 'sp4_r_v_b_11')
// (16, 19, 'sp4_v_b_10')
// (17, 13, 'sp4_v_t_38')
// (17, 14, 'sp4_v_b_38')
// (17, 15, 'sp4_h_l_46')
// (17, 15, 'sp4_h_r_11')
// (17, 15, 'sp4_v_b_27')
// (17, 15, 'sp4_v_t_46')
// (17, 16, 'neigh_op_tnl_1')
// (17, 16, 'sp4_v_b_14')
// (17, 16, 'sp4_v_b_46')
// (17, 17, 'neigh_op_lft_1')
// (17, 17, 'sp4_h_r_31')
// (17, 17, 'sp4_v_b_3')
// (17, 17, 'sp4_v_b_35')
// (17, 18, 'neigh_op_bnl_1')
// (17, 18, 'sp4_v_b_22')
// (17, 19, 'sp4_v_b_11')
// (18, 10, 'sp4_r_v_b_41')
// (18, 11, 'sp4_r_v_b_28')
// (18, 12, 'sp4_r_v_b_17')
// (18, 13, 'sp4_r_v_b_4')
// (18, 14, 'sp4_r_v_b_36')
// (18, 15, 'sp4_h_r_22')
// (18, 15, 'sp4_r_v_b_25')
// (18, 16, 'sp4_r_v_b_12')
// (18, 17, 'sp4_h_r_42')
// (18, 17, 'sp4_r_v_b_1')
// (19, 9, 'sp4_h_r_9')
// (19, 9, 'sp4_v_t_41')
// (19, 10, 'sp4_v_b_41')
// (19, 11, 'sp4_v_b_28')
// (19, 12, 'sp4_v_b_17')
// (19, 13, 'sp4_v_b_4')
// (19, 13, 'sp4_v_t_36')
// (19, 14, 'sp4_v_b_36')
// (19, 15, 'sp4_h_r_35')
// (19, 15, 'sp4_v_b_25')
// (19, 16, 'sp4_v_b_12')
// (19, 17, 'sp4_h_l_42')
// (19, 17, 'sp4_v_b_1')
// (20, 9, 'sp4_h_r_20')
// (20, 12, 'sp4_r_v_b_40')
// (20, 13, 'sp4_r_v_b_29')
// (20, 14, 'sp4_r_v_b_16')
// (20, 15, 'sp4_h_r_46')
// (20, 15, 'sp4_r_v_b_5')
// (21, 9, 'sp4_h_r_33')
// (21, 11, 'sp4_h_r_5')
// (21, 11, 'sp4_v_t_40')
// (21, 12, 'sp4_v_b_40')
// (21, 13, 'sp4_v_b_29')
// (21, 14, 'sp4_v_b_16')
// (21, 15, 'sp4_h_l_46')
// (21, 15, 'sp4_v_b_5')
// (22, 6, 'sp4_r_v_b_38')
// (22, 7, 'sp4_r_v_b_27')
// (22, 8, 'local_g2_6')
// (22, 8, 'lutff_0/in_0')
// (22, 8, 'lutff_1/in_1')
// (22, 8, 'lutff_6/in_0')
// (22, 8, 'sp4_r_v_b_14')
// (22, 9, 'sp4_h_r_44')
// (22, 9, 'sp4_r_v_b_3')
// (22, 11, 'local_g0_0')
// (22, 11, 'lutff_2/in_0')
// (22, 11, 'sp4_h_r_16')
// (23, 5, 'sp4_v_t_38')
// (23, 6, 'sp4_v_b_38')
// (23, 7, 'sp4_v_b_27')
// (23, 8, 'sp4_v_b_14')
// (23, 9, 'sp4_h_l_44')
// (23, 9, 'sp4_v_b_3')
// (23, 11, 'sp4_h_r_29')
// (24, 11, 'sp4_h_r_40')
// (25, 11, 'sp4_h_l_40')

wire n1646;
// (11, 18, 'neigh_op_tnr_0')
// (11, 19, 'neigh_op_rgt_0')
// (11, 20, 'neigh_op_bnr_0')
// (12, 17, 'sp4_r_v_b_41')
// (12, 18, 'neigh_op_top_0')
// (12, 18, 'sp4_r_v_b_28')
// (12, 19, 'local_g3_0')
// (12, 19, 'lutff_0/out')
// (12, 19, 'lutff_1/in_2')
// (12, 19, 'lutff_3/in_2')
// (12, 19, 'lutff_7/in_0')
// (12, 19, 'sp4_r_v_b_17')
// (12, 20, 'neigh_op_bot_0')
// (12, 20, 'sp4_r_v_b_4')
// (13, 16, 'sp4_v_t_41')
// (13, 17, 'sp4_v_b_41')
// (13, 18, 'neigh_op_tnl_0')
// (13, 18, 'sp4_v_b_28')
// (13, 19, 'local_g1_0')
// (13, 19, 'lutff_7/in_2')
// (13, 19, 'neigh_op_lft_0')
// (13, 19, 'sp4_v_b_17')
// (13, 20, 'neigh_op_bnl_0')
// (13, 20, 'sp4_h_r_4')
// (13, 20, 'sp4_v_b_4')
// (14, 20, 'sp4_h_r_17')
// (15, 20, 'local_g3_4')
// (15, 20, 'lutff_0/in_3')
// (15, 20, 'lutff_2/in_3')
// (15, 20, 'lutff_6/in_1')
// (15, 20, 'sp4_h_r_28')
// (16, 20, 'sp4_h_r_41')
// (17, 20, 'sp4_h_l_41')

reg n1647 = 0;
// (11, 18, 'neigh_op_tnr_3')
// (11, 19, 'neigh_op_rgt_3')
// (11, 20, 'neigh_op_bnr_3')
// (12, 5, 'sp4_r_v_b_41')
// (12, 6, 'sp4_r_v_b_28')
// (12, 7, 'sp4_r_v_b_17')
// (12, 8, 'sp4_r_v_b_4')
// (12, 9, 'sp4_r_v_b_41')
// (12, 10, 'sp4_r_v_b_28')
// (12, 11, 'sp4_r_v_b_17')
// (12, 12, 'sp4_r_v_b_4')
// (12, 13, 'sp4_r_v_b_36')
// (12, 14, 'sp4_r_v_b_25')
// (12, 15, 'sp4_r_v_b_12')
// (12, 16, 'sp4_r_v_b_1')
// (12, 17, 'sp4_r_v_b_47')
// (12, 18, 'local_g1_3')
// (12, 18, 'lutff_7/in_3')
// (12, 18, 'neigh_op_top_3')
// (12, 18, 'sp4_r_v_b_34')
// (12, 19, 'lutff_3/out')
// (12, 19, 'sp4_h_r_6')
// (12, 19, 'sp4_r_v_b_23')
// (12, 20, 'neigh_op_bot_3')
// (12, 20, 'sp4_r_v_b_10')
// (13, 4, 'sp4_h_r_9')
// (13, 4, 'sp4_v_t_41')
// (13, 5, 'sp4_v_b_41')
// (13, 6, 'sp4_v_b_28')
// (13, 7, 'sp4_v_b_17')
// (13, 8, 'sp4_v_b_4')
// (13, 8, 'sp4_v_t_41')
// (13, 9, 'sp4_v_b_41')
// (13, 10, 'sp4_v_b_28')
// (13, 11, 'sp4_v_b_17')
// (13, 12, 'sp4_v_b_4')
// (13, 12, 'sp4_v_t_36')
// (13, 13, 'sp4_v_b_36')
// (13, 14, 'sp4_v_b_25')
// (13, 15, 'sp4_v_b_12')
// (13, 16, 'sp4_v_b_1')
// (13, 16, 'sp4_v_t_47')
// (13, 17, 'sp4_v_b_47')
// (13, 18, 'neigh_op_tnl_3')
// (13, 18, 'sp4_v_b_34')
// (13, 19, 'local_g0_3')
// (13, 19, 'lutff_6/in_1')
// (13, 19, 'neigh_op_lft_3')
// (13, 19, 'sp4_h_r_19')
// (13, 19, 'sp4_v_b_23')
// (13, 20, 'local_g3_3')
// (13, 20, 'lutff_6/in_2')
// (13, 20, 'neigh_op_bnl_3')
// (13, 20, 'sp4_v_b_10')
// (14, 4, 'local_g0_4')
// (14, 4, 'lutff_4/in_0')
// (14, 4, 'sp4_h_r_20')
// (14, 19, 'local_g3_6')
// (14, 19, 'lutff_6/in_3')
// (14, 19, 'sp4_h_r_30')
// (15, 4, 'sp4_h_r_33')
// (15, 19, 'sp4_h_r_43')
// (16, 4, 'sp4_h_r_44')
// (16, 19, 'sp4_h_l_43')
// (17, 4, 'sp4_h_l_44')

reg n1648 = 0;
// (11, 18, 'neigh_op_tnr_7')
// (11, 19, 'neigh_op_rgt_7')
// (11, 20, 'neigh_op_bnr_7')
// (12, 1, 'sp4_r_v_b_40')
// (12, 2, 'sp4_r_v_b_29')
// (12, 3, 'sp4_r_v_b_16')
// (12, 4, 'sp4_r_v_b_5')
// (12, 5, 'sp4_r_v_b_44')
// (12, 6, 'sp4_r_v_b_33')
// (12, 7, 'sp4_r_v_b_20')
// (12, 8, 'sp4_r_v_b_9')
// (12, 9, 'sp4_r_v_b_43')
// (12, 10, 'sp4_r_v_b_30')
// (12, 11, 'sp4_r_v_b_19')
// (12, 12, 'sp4_r_v_b_6')
// (12, 13, 'sp4_r_v_b_47')
// (12, 14, 'sp4_r_v_b_34')
// (12, 15, 'sp4_r_v_b_23')
// (12, 16, 'sp4_r_v_b_10')
// (12, 17, 'sp4_r_v_b_39')
// (12, 18, 'neigh_op_top_7')
// (12, 18, 'sp4_r_v_b_26')
// (12, 19, 'lutff_7/out')
// (12, 19, 'sp4_r_v_b_15')
// (12, 20, 'neigh_op_bot_7')
// (12, 20, 'sp4_r_v_b_2')
// (13, 0, 'span4_vert_40')
// (13, 1, 'sp4_v_b_40')
// (13, 2, 'sp4_v_b_29')
// (13, 3, 'local_g0_0')
// (13, 3, 'lutff_2/in_0')
// (13, 3, 'sp4_v_b_16')
// (13, 4, 'sp4_v_b_5')
// (13, 4, 'sp4_v_t_44')
// (13, 5, 'sp4_v_b_44')
// (13, 6, 'sp4_v_b_33')
// (13, 7, 'sp4_v_b_20')
// (13, 8, 'sp4_v_b_9')
// (13, 8, 'sp4_v_t_43')
// (13, 9, 'sp4_v_b_43')
// (13, 10, 'sp4_v_b_30')
// (13, 11, 'sp4_v_b_19')
// (13, 12, 'sp4_v_b_6')
// (13, 12, 'sp4_v_t_47')
// (13, 13, 'sp4_v_b_47')
// (13, 14, 'sp4_v_b_34')
// (13, 15, 'sp4_v_b_23')
// (13, 16, 'sp4_v_b_10')
// (13, 16, 'sp4_v_t_39')
// (13, 17, 'sp4_v_b_39')
// (13, 18, 'local_g3_7')
// (13, 18, 'lutff_5/in_3')
// (13, 18, 'neigh_op_tnl_7')
// (13, 18, 'sp4_v_b_26')
// (13, 19, 'local_g1_7')
// (13, 19, 'lutff_5/in_1')
// (13, 19, 'neigh_op_lft_7')
// (13, 19, 'sp4_v_b_15')
// (13, 20, 'local_g3_7')
// (13, 20, 'lutff_5/in_1')
// (13, 20, 'neigh_op_bnl_7')
// (13, 20, 'sp4_v_b_2')

reg n1649 = 0;
// (11, 18, 'sp4_h_r_4')
// (11, 19, 'sp4_h_r_3')
// (12, 18, 'sp4_h_r_17')
// (12, 19, 'sp4_h_r_14')
// (12, 20, 'sp4_h_r_9')
// (13, 18, 'local_g2_4')
// (13, 18, 'lutff_5/in_1')
// (13, 18, 'sp4_h_r_28')
// (13, 19, 'local_g2_3')
// (13, 19, 'lutff_3/in_2')
// (13, 19, 'sp4_h_r_27')
// (13, 20, 'local_g1_4')
// (13, 20, 'lutff_3/in_2')
// (13, 20, 'sp4_h_r_20')
// (14, 2, 'sp4_r_v_b_36')
// (14, 3, 'sp4_r_v_b_25')
// (14, 4, 'sp4_r_v_b_12')
// (14, 5, 'sp4_r_v_b_1')
// (14, 6, 'sp4_r_v_b_36')
// (14, 7, 'sp4_r_v_b_25')
// (14, 8, 'sp4_r_v_b_12')
// (14, 9, 'sp4_r_v_b_1')
// (14, 10, 'sp4_r_v_b_40')
// (14, 11, 'sp4_r_v_b_29')
// (14, 12, 'sp4_r_v_b_16')
// (14, 13, 'sp4_r_v_b_5')
// (14, 14, 'sp4_r_v_b_44')
// (14, 15, 'sp4_r_v_b_33')
// (14, 16, 'sp4_r_v_b_20')
// (14, 17, 'sp4_r_v_b_9')
// (14, 18, 'sp4_h_r_41')
// (14, 18, 'sp4_r_v_b_36')
// (14, 19, 'neigh_op_tnr_6')
// (14, 19, 'sp4_h_r_38')
// (14, 19, 'sp4_r_v_b_25')
// (14, 19, 'sp4_r_v_b_41')
// (14, 20, 'neigh_op_rgt_6')
// (14, 20, 'sp4_h_r_33')
// (14, 20, 'sp4_r_v_b_12')
// (14, 20, 'sp4_r_v_b_28')
// (14, 20, 'sp4_r_v_b_44')
// (14, 21, 'neigh_op_bnr_6')
// (14, 21, 'sp4_r_v_b_1')
// (14, 21, 'sp4_r_v_b_17')
// (14, 21, 'sp4_r_v_b_33')
// (14, 22, 'sp4_r_v_b_20')
// (14, 22, 'sp4_r_v_b_4')
// (14, 23, 'sp4_r_v_b_9')
// (15, 1, 'sp4_v_t_36')
// (15, 2, 'local_g2_4')
// (15, 2, 'lutff_1/in_3')
// (15, 2, 'sp4_v_b_36')
// (15, 3, 'sp4_v_b_25')
// (15, 4, 'sp4_v_b_12')
// (15, 5, 'sp4_v_b_1')
// (15, 5, 'sp4_v_t_36')
// (15, 6, 'sp4_v_b_36')
// (15, 7, 'sp4_v_b_25')
// (15, 8, 'sp4_v_b_12')
// (15, 9, 'sp4_v_b_1')
// (15, 9, 'sp4_v_t_40')
// (15, 10, 'sp4_v_b_40')
// (15, 11, 'sp4_v_b_29')
// (15, 12, 'sp4_v_b_16')
// (15, 13, 'sp4_v_b_5')
// (15, 13, 'sp4_v_t_44')
// (15, 14, 'sp4_v_b_44')
// (15, 15, 'sp4_v_b_33')
// (15, 16, 'sp4_v_b_20')
// (15, 17, 'sp4_v_b_9')
// (15, 17, 'sp4_v_t_36')
// (15, 18, 'sp4_h_l_41')
// (15, 18, 'sp4_v_b_36')
// (15, 18, 'sp4_v_t_41')
// (15, 19, 'neigh_op_top_6')
// (15, 19, 'sp4_h_l_38')
// (15, 19, 'sp4_v_b_25')
// (15, 19, 'sp4_v_b_41')
// (15, 19, 'sp4_v_t_44')
// (15, 20, 'lutff_6/out')
// (15, 20, 'sp4_h_r_44')
// (15, 20, 'sp4_v_b_12')
// (15, 20, 'sp4_v_b_28')
// (15, 20, 'sp4_v_b_44')
// (15, 21, 'neigh_op_bot_6')
// (15, 21, 'sp4_v_b_1')
// (15, 21, 'sp4_v_b_17')
// (15, 21, 'sp4_v_b_33')
// (15, 22, 'sp4_v_b_20')
// (15, 22, 'sp4_v_b_4')
// (15, 23, 'sp4_v_b_9')
// (16, 19, 'neigh_op_tnl_6')
// (16, 20, 'neigh_op_lft_6')
// (16, 20, 'sp4_h_l_44')
// (16, 21, 'neigh_op_bnl_6')

reg n1650 = 0;
// (11, 18, 'sp4_h_r_6')
// (12, 17, 'neigh_op_tnr_7')
// (12, 18, 'neigh_op_rgt_7')
// (12, 18, 'sp4_h_r_19')
// (12, 19, 'neigh_op_bnr_7')
// (13, 14, 'sp4_r_v_b_43')
// (13, 15, 'sp4_r_v_b_30')
// (13, 16, 'sp4_r_v_b_19')
// (13, 17, 'local_g1_7')
// (13, 17, 'lutff_7/in_1')
// (13, 17, 'neigh_op_top_7')
// (13, 17, 'sp4_r_v_b_6')
// (13, 18, 'local_g1_7')
// (13, 18, 'lutff_7/in_1')
// (13, 18, 'lutff_7/out')
// (13, 18, 'sp4_h_r_30')
// (13, 18, 'sp4_r_v_b_47')
// (13, 19, 'neigh_op_bot_7')
// (13, 19, 'sp4_r_v_b_34')
// (13, 20, 'sp4_r_v_b_23')
// (13, 21, 'sp4_r_v_b_10')
// (14, 13, 'sp4_v_t_43')
// (14, 14, 'sp4_v_b_43')
// (14, 15, 'local_g3_6')
// (14, 15, 'lutff_6/in_3')
// (14, 15, 'sp4_v_b_30')
// (14, 16, 'sp4_v_b_19')
// (14, 17, 'neigh_op_tnl_7')
// (14, 17, 'sp4_v_b_6')
// (14, 17, 'sp4_v_t_47')
// (14, 18, 'neigh_op_lft_7')
// (14, 18, 'sp4_h_r_43')
// (14, 18, 'sp4_v_b_47')
// (14, 19, 'neigh_op_bnl_7')
// (14, 19, 'sp4_v_b_34')
// (14, 20, 'sp4_v_b_23')
// (14, 21, 'sp4_v_b_10')
// (15, 18, 'sp4_h_l_43')
// (15, 18, 'sp4_h_r_9')
// (16, 18, 'sp4_h_r_20')
// (17, 18, 'sp4_h_r_33')
// (18, 15, 'sp4_r_v_b_44')
// (18, 16, 'sp4_r_v_b_33')
// (18, 17, 'sp4_r_v_b_20')
// (18, 18, 'sp4_h_r_44')
// (18, 18, 'sp4_r_v_b_9')
// (19, 14, 'sp4_v_t_44')
// (19, 15, 'sp4_v_b_44')
// (19, 16, 'local_g2_1')
// (19, 16, 'ram/WADDR_4')
// (19, 16, 'sp4_v_b_33')
// (19, 17, 'sp4_v_b_20')
// (19, 18, 'sp4_h_l_44')
// (19, 18, 'sp4_v_b_9')

reg n1651 = 0;
// (11, 18, 'sp4_h_r_8')
// (12, 17, 'neigh_op_tnr_0')
// (12, 18, 'neigh_op_rgt_0')
// (12, 18, 'sp4_h_r_21')
// (12, 19, 'neigh_op_bnr_0')
// (13, 15, 'sp4_r_v_b_36')
// (13, 16, 'sp4_r_v_b_25')
// (13, 17, 'neigh_op_top_0')
// (13, 17, 'sp4_r_v_b_12')
// (13, 18, 'local_g2_0')
// (13, 18, 'lutff_0/in_2')
// (13, 18, 'lutff_0/out')
// (13, 18, 'sp4_h_r_32')
// (13, 18, 'sp4_r_v_b_1')
// (13, 19, 'neigh_op_bot_0')
// (14, 14, 'sp4_v_t_36')
// (14, 15, 'local_g2_4')
// (14, 15, 'lutff_7/in_3')
// (14, 15, 'sp4_v_b_36')
// (14, 16, 'sp4_v_b_25')
// (14, 17, 'neigh_op_tnl_0')
// (14, 17, 'sp4_v_b_12')
// (14, 18, 'neigh_op_lft_0')
// (14, 18, 'sp4_h_r_45')
// (14, 18, 'sp4_v_b_1')
// (14, 19, 'neigh_op_bnl_0')
// (15, 18, 'sp4_h_l_45')
// (15, 18, 'sp4_h_r_11')
// (16, 18, 'sp4_h_r_22')
// (17, 18, 'sp4_h_r_35')
// (18, 15, 'sp4_r_v_b_46')
// (18, 16, 'sp4_r_v_b_35')
// (18, 17, 'sp4_r_v_b_22')
// (18, 18, 'sp4_h_r_46')
// (18, 18, 'sp4_r_v_b_11')
// (19, 14, 'sp4_v_t_46')
// (19, 15, 'sp4_v_b_46')
// (19, 16, 'local_g3_3')
// (19, 16, 'ram/WADDR_5')
// (19, 16, 'sp4_v_b_35')
// (19, 17, 'sp4_v_b_22')
// (19, 18, 'sp4_h_l_46')
// (19, 18, 'sp4_v_b_11')

reg n1652 = 0;
// (11, 18, 'sp4_r_v_b_38')
// (11, 19, 'neigh_op_tnr_7')
// (11, 19, 'sp4_r_v_b_27')
// (11, 20, 'neigh_op_rgt_7')
// (11, 20, 'sp4_h_r_3')
// (11, 20, 'sp4_r_v_b_14')
// (11, 21, 'neigh_op_bnr_7')
// (11, 21, 'sp4_r_v_b_3')
// (12, 17, 'local_g0_0')
// (12, 17, 'local_g1_0')
// (12, 17, 'lutff_1/in_1')
// (12, 17, 'lutff_2/in_1')
// (12, 17, 'sp4_h_r_8')
// (12, 17, 'sp4_v_t_38')
// (12, 18, 'local_g3_6')
// (12, 18, 'lutff_2/in_1')
// (12, 18, 'sp4_v_b_38')
// (12, 19, 'local_g0_7')
// (12, 19, 'lutff_0/in_3')
// (12, 19, 'neigh_op_top_7')
// (12, 19, 'sp4_v_b_27')
// (12, 20, 'local_g2_7')
// (12, 20, 'lutff_1/in_2')
// (12, 20, 'lutff_4/in_3')
// (12, 20, 'lutff_7/in_2')
// (12, 20, 'lutff_7/out')
// (12, 20, 'sp4_h_r_14')
// (12, 20, 'sp4_v_b_14')
// (12, 21, 'neigh_op_bot_7')
// (12, 21, 'sp4_v_b_3')
// (13, 17, 'sp4_h_r_21')
// (13, 19, 'neigh_op_tnl_7')
// (13, 20, 'neigh_op_lft_7')
// (13, 20, 'sp4_h_r_27')
// (13, 21, 'local_g3_7')
// (13, 21, 'lutff_4/in_2')
// (13, 21, 'lutff_7/in_1')
// (13, 21, 'neigh_op_bnl_7')
// (14, 17, 'sp4_h_r_32')
// (14, 17, 'sp4_r_v_b_44')
// (14, 18, 'sp4_r_v_b_33')
// (14, 19, 'sp4_r_v_b_20')
// (14, 20, 'sp4_h_r_38')
// (14, 20, 'sp4_r_v_b_9')
// (15, 16, 'sp4_v_t_44')
// (15, 17, 'sp4_h_r_45')
// (15, 17, 'sp4_v_b_44')
// (15, 18, 'sp4_v_b_33')
// (15, 19, 'local_g1_4')
// (15, 19, 'lutff_7/in_0')
// (15, 19, 'sp4_v_b_20')
// (15, 20, 'local_g1_1')
// (15, 20, 'lutff_7/in_1')
// (15, 20, 'sp4_h_l_38')
// (15, 20, 'sp4_v_b_9')
// (16, 17, 'sp4_h_l_45')

reg n1653 = 0;
// (11, 19, 'local_g3_4')
// (11, 19, 'lutff_4/in_1')
// (11, 19, 'neigh_op_tnr_4')
// (11, 20, 'neigh_op_rgt_4')
// (11, 21, 'neigh_op_bnr_4')
// (12, 19, 'neigh_op_top_4')
// (12, 20, 'local_g0_4')
// (12, 20, 'local_g3_4')
// (12, 20, 'lutff_1/in_3')
// (12, 20, 'lutff_4/in_2')
// (12, 20, 'lutff_4/out')
// (12, 20, 'lutff_7/in_0')
// (12, 21, 'neigh_op_bot_4')
// (13, 19, 'neigh_op_tnl_4')
// (13, 20, 'neigh_op_lft_4')
// (13, 21, 'neigh_op_bnl_4')

wire n1654;
// (11, 19, 'neigh_op_tnr_1')
// (11, 20, 'neigh_op_rgt_1')
// (11, 20, 'sp4_h_r_7')
// (11, 21, 'neigh_op_bnr_1')
// (12, 19, 'neigh_op_top_1')
// (12, 20, 'local_g0_2')
// (12, 20, 'lutff_1/out')
// (12, 20, 'lutff_global/cen')
// (12, 20, 'sp4_h_r_18')
// (12, 21, 'neigh_op_bot_1')
// (13, 19, 'neigh_op_tnl_1')
// (13, 20, 'neigh_op_lft_1')
// (13, 20, 'sp4_h_r_31')
// (13, 21, 'neigh_op_bnl_1')
// (14, 20, 'sp4_h_r_42')
// (15, 20, 'sp4_h_l_42')

wire n1655;
// (11, 20, 'neigh_op_tnr_1')
// (11, 21, 'neigh_op_rgt_1')
// (11, 22, 'neigh_op_bnr_1')
// (12, 20, 'neigh_op_top_1')
// (12, 21, 'lutff_1/out')
// (12, 22, 'neigh_op_bot_1')
// (13, 20, 'neigh_op_tnl_1')
// (13, 21, 'local_g0_1')
// (13, 21, 'lutff_1/in_0')
// (13, 21, 'neigh_op_lft_1')
// (13, 22, 'neigh_op_bnl_1')

wire n1656;
// (11, 20, 'neigh_op_tnr_2')
// (11, 21, 'neigh_op_rgt_2')
// (11, 22, 'neigh_op_bnr_2')
// (12, 20, 'neigh_op_top_2')
// (12, 21, 'lutff_2/out')
// (12, 22, 'neigh_op_bot_2')
// (13, 20, 'neigh_op_tnl_2')
// (13, 21, 'local_g1_2')
// (13, 21, 'lutff_6/in_3')
// (13, 21, 'neigh_op_lft_2')
// (13, 22, 'neigh_op_bnl_2')

wire n1657;
// (11, 20, 'neigh_op_tnr_3')
// (11, 21, 'neigh_op_rgt_3')
// (11, 22, 'neigh_op_bnr_3')
// (12, 20, 'neigh_op_top_3')
// (12, 21, 'lutff_3/out')
// (12, 22, 'neigh_op_bot_3')
// (13, 20, 'neigh_op_tnl_3')
// (13, 21, 'local_g0_3')
// (13, 21, 'lutff_2/in_3')
// (13, 21, 'neigh_op_lft_3')
// (13, 22, 'neigh_op_bnl_3')

wire n1658;
// (11, 20, 'neigh_op_tnr_7')
// (11, 21, 'neigh_op_rgt_7')
// (11, 21, 'sp4_h_r_3')
// (11, 21, 'sp4_h_r_6')
// (11, 22, 'neigh_op_bnr_7')
// (12, 20, 'neigh_op_top_7')
// (12, 21, 'local_g1_3')
// (12, 21, 'lutff_7/out')
// (12, 21, 'lutff_global/cen')
// (12, 21, 'sp4_h_r_14')
// (12, 21, 'sp4_h_r_19')
// (12, 22, 'neigh_op_bot_7')
// (13, 20, 'neigh_op_tnl_7')
// (13, 21, 'neigh_op_lft_7')
// (13, 21, 'sp4_h_r_27')
// (13, 21, 'sp4_h_r_30')
// (13, 22, 'neigh_op_bnl_7')
// (14, 21, 'sp4_h_r_38')
// (14, 21, 'sp4_h_r_43')
// (15, 21, 'sp4_h_l_38')
// (15, 21, 'sp4_h_l_43')
// (15, 21, 'sp4_h_r_6')
// (16, 21, 'sp4_h_r_19')
// (17, 21, 'sp4_h_r_30')
// (18, 21, 'sp4_h_r_43')
// (19, 21, 'sp4_h_l_43')

wire n1659;
// (11, 21, 'neigh_op_tnr_1')
// (11, 22, 'neigh_op_rgt_1')
// (11, 23, 'neigh_op_bnr_1')
// (12, 21, 'neigh_op_top_1')
// (12, 22, 'lutff_1/out')
// (12, 23, 'local_g1_1')
// (12, 23, 'lutff_4/in_0')
// (12, 23, 'neigh_op_bot_1')
// (13, 21, 'neigh_op_tnl_1')
// (13, 22, 'neigh_op_lft_1')
// (13, 23, 'neigh_op_bnl_1')

wire n1660;
// (11, 21, 'neigh_op_tnr_2')
// (11, 22, 'neigh_op_rgt_2')
// (11, 23, 'neigh_op_bnr_2')
// (12, 21, 'neigh_op_top_2')
// (12, 22, 'lutff_2/out')
// (12, 23, 'neigh_op_bot_2')
// (13, 21, 'neigh_op_tnl_2')
// (13, 22, 'local_g0_2')
// (13, 22, 'lutff_2/in_2')
// (13, 22, 'neigh_op_lft_2')
// (13, 23, 'neigh_op_bnl_2')

wire n1661;
// (11, 21, 'neigh_op_tnr_3')
// (11, 22, 'neigh_op_rgt_3')
// (11, 23, 'neigh_op_bnr_3')
// (12, 21, 'neigh_op_top_3')
// (12, 22, 'lutff_3/out')
// (12, 23, 'neigh_op_bot_3')
// (13, 21, 'neigh_op_tnl_3')
// (13, 22, 'local_g1_3')
// (13, 22, 'lutff_4/in_0')
// (13, 22, 'neigh_op_lft_3')
// (13, 23, 'neigh_op_bnl_3')

wire n1662;
// (11, 21, 'neigh_op_tnr_4')
// (11, 22, 'neigh_op_rgt_4')
// (11, 23, 'neigh_op_bnr_4')
// (12, 21, 'neigh_op_top_4')
// (12, 22, 'lutff_4/out')
// (12, 23, 'neigh_op_bot_4')
// (13, 21, 'neigh_op_tnl_4')
// (13, 22, 'neigh_op_lft_4')
// (13, 23, 'local_g2_4')
// (13, 23, 'lutff_7/in_3')
// (13, 23, 'neigh_op_bnl_4')

wire n1663;
// (11, 21, 'neigh_op_tnr_5')
// (11, 22, 'neigh_op_rgt_5')
// (11, 23, 'neigh_op_bnr_5')
// (12, 21, 'neigh_op_top_5')
// (12, 22, 'lutff_5/out')
// (12, 23, 'neigh_op_bot_5')
// (13, 21, 'neigh_op_tnl_5')
// (13, 22, 'local_g1_5')
// (13, 22, 'lutff_6/in_0')
// (13, 22, 'neigh_op_lft_5')
// (13, 23, 'neigh_op_bnl_5')

wire n1664;
// (11, 21, 'neigh_op_tnr_6')
// (11, 22, 'neigh_op_rgt_6')
// (11, 23, 'neigh_op_bnr_6')
// (12, 21, 'neigh_op_top_6')
// (12, 22, 'local_g0_6')
// (12, 22, 'lutff_6/out')
// (12, 22, 'lutff_7/in_1')
// (12, 23, 'neigh_op_bot_6')
// (13, 21, 'neigh_op_tnl_6')
// (13, 22, 'neigh_op_lft_6')
// (13, 23, 'neigh_op_bnl_6')

reg n1665 = 0;
// (11, 21, 'neigh_op_tnr_7')
// (11, 22, 'neigh_op_rgt_7')
// (11, 22, 'sp4_h_r_3')
// (11, 23, 'neigh_op_bnr_7')
// (12, 20, 'sp4_r_v_b_39')
// (12, 21, 'neigh_op_top_7')
// (12, 21, 'sp4_r_v_b_26')
// (12, 22, 'local_g3_7')
// (12, 22, 'lutff_6/in_2')
// (12, 22, 'lutff_7/out')
// (12, 22, 'sp4_h_r_14')
// (12, 22, 'sp4_r_v_b_15')
// (12, 23, 'neigh_op_bot_7')
// (12, 23, 'sp4_r_v_b_2')
// (13, 19, 'sp4_v_t_39')
// (13, 20, 'sp4_v_b_39')
// (13, 21, 'local_g2_7')
// (13, 21, 'lutff_4/in_1')
// (13, 21, 'neigh_op_tnl_7')
// (13, 21, 'sp4_v_b_26')
// (13, 22, 'neigh_op_lft_7')
// (13, 22, 'sp4_h_r_27')
// (13, 22, 'sp4_v_b_15')
// (13, 23, 'neigh_op_bnl_7')
// (13, 23, 'sp4_h_r_8')
// (13, 23, 'sp4_v_b_2')
// (14, 19, 'sp4_r_v_b_38')
// (14, 20, 'sp4_r_v_b_27')
// (14, 21, 'local_g2_6')
// (14, 21, 'lutff_3/in_1')
// (14, 21, 'lutff_7/in_1')
// (14, 21, 'sp4_r_v_b_14')
// (14, 22, 'sp4_h_r_38')
// (14, 22, 'sp4_r_v_b_3')
// (14, 23, 'local_g0_5')
// (14, 23, 'lutff_6/in_1')
// (14, 23, 'sp4_h_r_21')
// (15, 18, 'sp4_v_t_38')
// (15, 19, 'sp4_v_b_38')
// (15, 20, 'sp4_v_b_27')
// (15, 21, 'sp4_v_b_14')
// (15, 22, 'sp4_h_l_38')
// (15, 22, 'sp4_v_b_3')
// (15, 23, 'sp4_h_r_32')
// (16, 23, 'sp4_h_r_45')
// (17, 23, 'sp4_h_l_45')

wire n1666;
// (11, 22, 'sp4_h_r_2')
// (11, 22, 'sp4_h_r_6')
// (12, 21, 'neigh_op_tnr_7')
// (12, 21, 'sp4_r_v_b_43')
// (12, 22, 'local_g1_3')
// (12, 22, 'lutff_global/cen')
// (12, 22, 'neigh_op_rgt_7')
// (12, 22, 'sp4_h_r_15')
// (12, 22, 'sp4_h_r_19')
// (12, 22, 'sp4_h_r_3')
// (12, 22, 'sp4_r_v_b_30')
// (12, 23, 'local_g3_3')
// (12, 23, 'lutff_global/cen')
// (12, 23, 'neigh_op_bnr_7')
// (12, 23, 'sp4_r_v_b_19')
// (12, 24, 'sp4_r_v_b_6')
// (13, 20, 'sp4_v_t_43')
// (13, 21, 'neigh_op_top_7')
// (13, 21, 'sp4_v_b_43')
// (13, 22, 'local_g2_2')
// (13, 22, 'lutff_7/out')
// (13, 22, 'lutff_global/cen')
// (13, 22, 'sp4_h_r_14')
// (13, 22, 'sp4_h_r_26')
// (13, 22, 'sp4_h_r_30')
// (13, 22, 'sp4_v_b_30')
// (13, 23, 'local_g1_3')
// (13, 23, 'lutff_global/cen')
// (13, 23, 'neigh_op_bot_7')
// (13, 23, 'sp4_v_b_19')
// (13, 24, 'sp4_v_b_6')
// (14, 21, 'neigh_op_tnl_7')
// (14, 22, 'neigh_op_lft_7')
// (14, 22, 'sp4_h_r_27')
// (14, 22, 'sp4_h_r_39')
// (14, 22, 'sp4_h_r_43')
// (14, 23, 'neigh_op_bnl_7')
// (15, 22, 'sp4_h_l_39')
// (15, 22, 'sp4_h_l_43')
// (15, 22, 'sp4_h_r_2')
// (15, 22, 'sp4_h_r_38')
// (16, 22, 'sp4_h_l_38')
// (16, 22, 'sp4_h_r_15')
// (17, 22, 'sp4_h_r_26')
// (18, 22, 'sp4_h_r_39')
// (19, 22, 'sp4_h_l_39')

wire n1667;
// (12, 1, 'lutff_7/cout')
// (12, 2, 'carry_in')
// (12, 2, 'carry_in_mux')
// (12, 2, 'lutff_0/in_3')

reg n1668 = 0;
// (12, 1, 'neigh_op_tnr_2')
// (12, 2, 'neigh_op_rgt_2')
// (12, 3, 'neigh_op_bnr_2')
// (13, 1, 'neigh_op_top_2')
// (13, 2, 'local_g3_2')
// (13, 2, 'lutff_2/out')
// (13, 2, 'lutff_6/in_1')
// (13, 3, 'neigh_op_bot_2')
// (14, 1, 'neigh_op_tnl_2')
// (14, 2, 'neigh_op_lft_2')
// (14, 3, 'neigh_op_bnl_2')

reg n1669 = 0;
// (12, 1, 'neigh_op_tnr_3')
// (12, 2, 'neigh_op_rgt_3')
// (12, 3, 'neigh_op_bnr_3')
// (13, 1, 'neigh_op_top_3')
// (13, 2, 'local_g0_3')
// (13, 2, 'lutff_3/out')
// (13, 2, 'lutff_5/in_2')
// (13, 3, 'neigh_op_bot_3')
// (14, 1, 'neigh_op_tnl_3')
// (14, 2, 'neigh_op_lft_3')
// (14, 3, 'neigh_op_bnl_3')

wire n1670;
// (12, 1, 'neigh_op_tnr_4')
// (12, 2, 'neigh_op_rgt_4')
// (12, 3, 'neigh_op_bnr_4')
// (13, 1, 'neigh_op_top_4')
// (13, 1, 'sp4_r_v_b_14')
// (13, 1, 'sp4_r_v_b_20')
// (13, 2, 'local_g1_3')
// (13, 2, 'lutff_4/out')
// (13, 2, 'lutff_global/cen')
// (13, 2, 'sp4_r_v_b_3')
// (13, 2, 'sp4_r_v_b_9')
// (13, 3, 'neigh_op_bot_4')
// (14, 0, 'span4_vert_14')
// (14, 0, 'span4_vert_20')
// (14, 1, 'local_g2_4')
// (14, 1, 'lutff_0/in_2')
// (14, 1, 'neigh_op_tnl_4')
// (14, 1, 'sp4_v_b_14')
// (14, 1, 'sp4_v_b_20')
// (14, 2, 'local_g1_3')
// (14, 2, 'lutff_global/cen')
// (14, 2, 'neigh_op_lft_4')
// (14, 2, 'sp4_h_r_3')
// (14, 2, 'sp4_v_b_3')
// (14, 2, 'sp4_v_b_9')
// (14, 3, 'neigh_op_bnl_4')
// (15, 2, 'sp4_h_r_14')
// (16, 2, 'sp4_h_r_27')
// (17, 2, 'sp4_h_r_38')
// (18, 2, 'sp4_h_l_38')

wire n1671;
// (12, 2, 'neigh_op_tnr_0')
// (12, 3, 'neigh_op_rgt_0')
// (12, 4, 'neigh_op_bnr_0')
// (13, 2, 'neigh_op_top_0')
// (13, 3, 'local_g1_0')
// (13, 3, 'lutff_0/out')
// (13, 3, 'lutff_2/in_3')
// (13, 4, 'neigh_op_bot_0')
// (14, 2, 'neigh_op_tnl_0')
// (14, 3, 'neigh_op_lft_0')
// (14, 4, 'neigh_op_bnl_0')

wire n1672;
// (12, 2, 'neigh_op_tnr_1')
// (12, 3, 'neigh_op_rgt_1')
// (12, 4, 'neigh_op_bnr_1')
// (13, 2, 'neigh_op_top_1')
// (13, 3, 'lutff_1/out')
// (13, 4, 'neigh_op_bot_1')
// (14, 2, 'neigh_op_tnl_1')
// (14, 3, 'local_g0_1')
// (14, 3, 'lutff_4/in_1')
// (14, 3, 'neigh_op_lft_1')
// (14, 4, 'neigh_op_bnl_1')

wire n1673;
// (12, 2, 'neigh_op_tnr_2')
// (12, 3, 'neigh_op_rgt_2')
// (12, 4, 'neigh_op_bnr_2')
// (13, 2, 'neigh_op_top_2')
// (13, 3, 'local_g3_2')
// (13, 3, 'lutff_2/out')
// (13, 3, 'lutff_3/in_2')
// (13, 4, 'neigh_op_bot_2')
// (14, 2, 'neigh_op_tnl_2')
// (14, 3, 'neigh_op_lft_2')
// (14, 4, 'neigh_op_bnl_2')

wire n1674;
// (12, 2, 'neigh_op_tnr_3')
// (12, 3, 'neigh_op_rgt_3')
// (12, 4, 'neigh_op_bnr_3')
// (13, 2, 'neigh_op_top_3')
// (13, 3, 'lutff_3/out')
// (13, 4, 'local_g0_3')
// (13, 4, 'lutff_2/in_1')
// (13, 4, 'neigh_op_bot_3')
// (14, 2, 'neigh_op_tnl_3')
// (14, 3, 'neigh_op_lft_3')
// (14, 4, 'neigh_op_bnl_3')

wire n1675;
// (12, 2, 'neigh_op_tnr_4')
// (12, 3, 'neigh_op_rgt_4')
// (12, 4, 'neigh_op_bnr_4')
// (13, 2, 'neigh_op_top_4')
// (13, 3, 'local_g3_4')
// (13, 3, 'lutff_4/out')
// (13, 3, 'lutff_7/in_2')
// (13, 4, 'neigh_op_bot_4')
// (14, 2, 'neigh_op_tnl_4')
// (14, 3, 'neigh_op_lft_4')
// (14, 4, 'neigh_op_bnl_4')

wire n1676;
// (12, 2, 'neigh_op_tnr_6')
// (12, 3, 'neigh_op_rgt_6')
// (12, 4, 'neigh_op_bnr_6')
// (13, 2, 'neigh_op_top_6')
// (13, 3, 'lutff_6/out')
// (13, 4, 'local_g0_6')
// (13, 4, 'lutff_5/in_3')
// (13, 4, 'neigh_op_bot_6')
// (14, 2, 'neigh_op_tnl_6')
// (14, 3, 'neigh_op_lft_6')
// (14, 4, 'neigh_op_bnl_6')

wire n1677;
// (12, 2, 'neigh_op_tnr_7')
// (12, 3, 'neigh_op_rgt_7')
// (12, 4, 'neigh_op_bnr_7')
// (13, 2, 'neigh_op_top_7')
// (13, 3, 'lutff_7/out')
// (13, 4, 'local_g0_7')
// (13, 4, 'lutff_7/in_0')
// (13, 4, 'neigh_op_bot_7')
// (14, 2, 'neigh_op_tnl_7')
// (14, 3, 'neigh_op_lft_7')
// (14, 4, 'neigh_op_bnl_7')

reg n1678 = 0;
// (12, 2, 'sp4_h_r_1')
// (13, 2, 'sp4_h_r_12')
// (14, 2, 'local_g3_1')
// (14, 2, 'lutff_4/in_2')
// (14, 2, 'sp4_h_r_25')
// (14, 4, 'sp4_r_v_b_38')
// (14, 5, 'sp4_r_v_b_27')
// (14, 6, 'sp4_r_v_b_14')
// (14, 7, 'local_g1_3')
// (14, 7, 'lutff_3/in_3')
// (14, 7, 'sp4_r_v_b_3')
// (15, 1, 'sp4_r_v_b_44')
// (15, 2, 'neigh_op_tnr_2')
// (15, 2, 'sp4_h_r_36')
// (15, 2, 'sp4_r_v_b_33')
// (15, 3, 'neigh_op_rgt_2')
// (15, 3, 'sp4_h_r_9')
// (15, 3, 'sp4_r_v_b_20')
// (15, 3, 'sp4_r_v_b_36')
// (15, 3, 'sp4_v_t_38')
// (15, 4, 'neigh_op_bnr_2')
// (15, 4, 'sp4_r_v_b_25')
// (15, 4, 'sp4_r_v_b_9')
// (15, 4, 'sp4_v_b_38')
// (15, 5, 'sp4_r_v_b_12')
// (15, 5, 'sp4_r_v_b_37')
// (15, 5, 'sp4_v_b_27')
// (15, 6, 'sp4_r_v_b_1')
// (15, 6, 'sp4_r_v_b_24')
// (15, 6, 'sp4_v_b_14')
// (15, 7, 'local_g2_5')
// (15, 7, 'lutff_2/in_3')
// (15, 7, 'sp4_r_v_b_13')
// (15, 7, 'sp4_v_b_3')
// (15, 8, 'sp4_r_v_b_0')
// (16, 0, 'span4_vert_44')
// (16, 1, 'sp4_v_b_44')
// (16, 2, 'neigh_op_top_2')
// (16, 2, 'sp4_h_l_36')
// (16, 2, 'sp4_v_b_33')
// (16, 2, 'sp4_v_t_36')
// (16, 3, 'lutff_2/out')
// (16, 3, 'sp4_h_r_20')
// (16, 3, 'sp4_v_b_20')
// (16, 3, 'sp4_v_b_36')
// (16, 4, 'neigh_op_bot_2')
// (16, 4, 'sp4_v_b_25')
// (16, 4, 'sp4_v_b_9')
// (16, 4, 'sp4_v_t_37')
// (16, 5, 'sp4_v_b_12')
// (16, 5, 'sp4_v_b_37')
// (16, 6, 'sp4_v_b_1')
// (16, 6, 'sp4_v_b_24')
// (16, 7, 'sp4_v_b_13')
// (16, 8, 'sp4_v_b_0')
// (17, 2, 'neigh_op_tnl_2')
// (17, 3, 'neigh_op_lft_2')
// (17, 3, 'sp4_h_r_33')
// (17, 4, 'neigh_op_bnl_2')
// (18, 3, 'sp4_h_r_44')
// (19, 3, 'sp4_h_l_44')

reg n1679 = 0;
// (12, 2, 'sp4_r_v_b_42')
// (12, 3, 'neigh_op_tnr_1')
// (12, 3, 'sp4_r_v_b_31')
// (12, 4, 'neigh_op_rgt_1')
// (12, 4, 'sp4_h_r_7')
// (12, 4, 'sp4_r_v_b_18')
// (12, 5, 'neigh_op_bnr_1')
// (12, 5, 'sp4_r_v_b_7')
// (13, 1, 'sp4_v_t_42')
// (13, 2, 'sp4_r_v_b_43')
// (13, 2, 'sp4_v_b_42')
// (13, 3, 'neigh_op_top_1')
// (13, 3, 'sp4_r_v_b_30')
// (13, 3, 'sp4_v_b_31')
// (13, 4, 'lutff_1/out')
// (13, 4, 'sp4_h_r_18')
// (13, 4, 'sp4_r_v_b_19')
// (13, 4, 'sp4_v_b_18')
// (13, 5, 'neigh_op_bot_1')
// (13, 5, 'sp4_h_r_7')
// (13, 5, 'sp4_r_v_b_6')
// (13, 5, 'sp4_v_b_7')
// (13, 6, 'sp4_r_v_b_44')
// (13, 7, 'sp4_r_v_b_33')
// (13, 8, 'local_g3_4')
// (13, 8, 'lutff_3/in_0')
// (13, 8, 'sp4_r_v_b_20')
// (13, 9, 'sp4_r_v_b_9')
// (14, 1, 'sp4_v_t_43')
// (14, 2, 'sp4_v_b_43')
// (14, 3, 'neigh_op_tnl_1')
// (14, 3, 'sp4_v_b_30')
// (14, 4, 'local_g1_1')
// (14, 4, 'lutff_2/in_2')
// (14, 4, 'neigh_op_lft_1')
// (14, 4, 'sp4_h_r_31')
// (14, 4, 'sp4_v_b_19')
// (14, 5, 'neigh_op_bnl_1')
// (14, 5, 'sp4_h_r_18')
// (14, 5, 'sp4_v_b_6')
// (14, 5, 'sp4_v_t_44')
// (14, 6, 'sp4_v_b_44')
// (14, 7, 'sp4_v_b_33')
// (14, 8, 'sp4_v_b_20')
// (14, 9, 'sp4_v_b_9')
// (15, 4, 'sp4_h_r_42')
// (15, 5, 'local_g2_7')
// (15, 5, 'lutff_1/in_2')
// (15, 5, 'sp4_h_r_31')
// (15, 5, 'sp4_r_v_b_42')
// (15, 6, 'sp4_r_v_b_31')
// (15, 7, 'sp4_r_v_b_18')
// (15, 8, 'sp4_r_v_b_7')
// (16, 4, 'sp4_h_l_42')
// (16, 4, 'sp4_v_t_42')
// (16, 5, 'sp4_h_r_42')
// (16, 5, 'sp4_v_b_42')
// (16, 6, 'local_g2_7')
// (16, 6, 'lutff_4/in_1')
// (16, 6, 'sp4_v_b_31')
// (16, 7, 'sp4_v_b_18')
// (16, 8, 'local_g0_7')
// (16, 8, 'lutff_6/in_3')
// (16, 8, 'sp4_v_b_7')
// (17, 5, 'sp4_h_l_42')

wire n1680;
// (12, 3, 'lutff_6/cout')
// (12, 3, 'lutff_7/in_3')

wire n1681;
// (12, 3, 'neigh_op_tnr_0')
// (12, 4, 'neigh_op_rgt_0')
// (12, 5, 'neigh_op_bnr_0')
// (13, 3, 'neigh_op_top_0')
// (13, 4, 'local_g3_0')
// (13, 4, 'lutff_0/out')
// (13, 4, 'lutff_5/in_0')
// (13, 5, 'neigh_op_bot_0')
// (14, 3, 'neigh_op_tnl_0')
// (14, 4, 'neigh_op_lft_0')
// (14, 5, 'neigh_op_bnl_0')

wire n1682;
// (12, 3, 'neigh_op_tnr_2')
// (12, 4, 'neigh_op_rgt_2')
// (12, 5, 'neigh_op_bnr_2')
// (13, 3, 'neigh_op_top_2')
// (13, 4, 'lutff_2/out')
// (13, 5, 'local_g1_2')
// (13, 5, 'lutff_2/in_3')
// (13, 5, 'neigh_op_bot_2')
// (14, 3, 'neigh_op_tnl_2')
// (14, 4, 'neigh_op_lft_2')
// (14, 5, 'neigh_op_bnl_2')

wire n1683;
// (12, 3, 'neigh_op_tnr_3')
// (12, 4, 'neigh_op_rgt_3')
// (12, 5, 'neigh_op_bnr_3')
// (13, 3, 'neigh_op_top_3')
// (13, 4, 'lutff_3/out')
// (13, 5, 'local_g0_3')
// (13, 5, 'lutff_4/in_3')
// (13, 5, 'neigh_op_bot_3')
// (14, 3, 'neigh_op_tnl_3')
// (14, 4, 'neigh_op_lft_3')
// (14, 5, 'neigh_op_bnl_3')

wire n1684;
// (12, 3, 'neigh_op_tnr_4')
// (12, 4, 'neigh_op_rgt_4')
// (12, 5, 'neigh_op_bnr_4')
// (13, 3, 'neigh_op_top_4')
// (13, 4, 'lutff_4/out')
// (13, 5, 'local_g0_4')
// (13, 5, 'lutff_3/in_3')
// (13, 5, 'neigh_op_bot_4')
// (14, 3, 'neigh_op_tnl_4')
// (14, 4, 'neigh_op_lft_4')
// (14, 5, 'neigh_op_bnl_4')

wire n1685;
// (12, 3, 'neigh_op_tnr_5')
// (12, 4, 'neigh_op_rgt_5')
// (12, 5, 'neigh_op_bnr_5')
// (13, 3, 'neigh_op_top_5')
// (13, 4, 'local_g1_5')
// (13, 4, 'lutff_3/in_3')
// (13, 4, 'lutff_5/out')
// (13, 5, 'neigh_op_bot_5')
// (14, 3, 'neigh_op_tnl_5')
// (14, 4, 'neigh_op_lft_5')
// (14, 5, 'neigh_op_bnl_5')

wire n1686;
// (12, 3, 'neigh_op_tnr_6')
// (12, 4, 'local_g2_6')
// (12, 4, 'lutff_4/in_2')
// (12, 4, 'neigh_op_rgt_6')
// (12, 5, 'neigh_op_bnr_6')
// (13, 3, 'neigh_op_top_6')
// (13, 4, 'lutff_6/out')
// (13, 5, 'neigh_op_bot_6')
// (14, 3, 'neigh_op_tnl_6')
// (14, 4, 'neigh_op_lft_6')
// (14, 5, 'neigh_op_bnl_6')

wire n1687;
// (12, 3, 'neigh_op_tnr_7')
// (12, 4, 'neigh_op_rgt_7')
// (12, 5, 'neigh_op_bnr_7')
// (13, 3, 'neigh_op_top_7')
// (13, 4, 'lutff_7/out')
// (13, 5, 'local_g0_7')
// (13, 5, 'lutff_6/in_1')
// (13, 5, 'neigh_op_bot_7')
// (14, 3, 'neigh_op_tnl_7')
// (14, 4, 'neigh_op_lft_7')
// (14, 5, 'neigh_op_bnl_7')

wire n1688;
// (12, 3, 'sp4_h_r_1')
// (13, 3, 'local_g0_4')
// (13, 3, 'lutff_3/in_3')
// (13, 3, 'sp4_h_r_12')
// (14, 0, 'logic_op_tnr_4')
// (14, 1, 'neigh_op_rgt_4')
// (14, 2, 'neigh_op_bnr_4')
// (14, 3, 'sp4_h_r_25')
// (15, 0, 'logic_op_top_4')
// (15, 1, 'lutff_4/out')
// (15, 1, 'sp4_r_v_b_25')
// (15, 2, 'neigh_op_bot_4')
// (15, 2, 'sp4_r_v_b_12')
// (15, 3, 'sp4_h_r_36')
// (15, 3, 'sp4_r_v_b_1')
// (16, 0, 'logic_op_tnl_4')
// (16, 0, 'span4_vert_25')
// (16, 1, 'neigh_op_lft_4')
// (16, 1, 'sp4_v_b_25')
// (16, 2, 'neigh_op_bnl_4')
// (16, 2, 'sp4_v_b_12')
// (16, 3, 'sp4_h_l_36')
// (16, 3, 'sp4_v_b_1')

reg n1689 = 0;
// (12, 3, 'sp4_h_r_11')
// (13, 3, 'local_g0_6')
// (13, 3, 'lutff_0/in_0')
// (13, 3, 'sp4_h_r_22')
// (13, 4, 'sp4_r_v_b_44')
// (13, 5, 'sp4_r_v_b_33')
// (13, 6, 'sp4_r_v_b_20')
// (13, 7, 'local_g2_1')
// (13, 7, 'lutff_0/in_1')
// (13, 7, 'sp4_r_v_b_9')
// (13, 8, 'local_g2_5')
// (13, 8, 'lutff_6/in_3')
// (13, 8, 'sp4_r_v_b_37')
// (13, 9, 'sp4_r_v_b_24')
// (13, 10, 'sp4_r_v_b_13')
// (13, 11, 'sp4_r_v_b_0')
// (14, 2, 'neigh_op_tnr_7')
// (14, 3, 'neigh_op_rgt_7')
// (14, 3, 'sp4_h_r_3')
// (14, 3, 'sp4_h_r_35')
// (14, 3, 'sp4_r_v_b_46')
// (14, 3, 'sp4_v_t_44')
// (14, 4, 'neigh_op_bnr_7')
// (14, 4, 'sp4_r_v_b_35')
// (14, 4, 'sp4_v_b_44')
// (14, 5, 'sp4_r_v_b_22')
// (14, 5, 'sp4_v_b_33')
// (14, 6, 'sp4_r_v_b_11')
// (14, 6, 'sp4_v_b_20')
// (14, 7, 'sp4_v_b_9')
// (14, 7, 'sp4_v_t_37')
// (14, 8, 'sp4_v_b_37')
// (14, 9, 'sp4_v_b_24')
// (14, 10, 'sp4_v_b_13')
// (14, 11, 'sp4_v_b_0')
// (15, 0, 'span12_vert_18')
// (15, 1, 'sp12_v_b_18')
// (15, 2, 'neigh_op_top_7')
// (15, 2, 'sp12_v_b_17')
// (15, 2, 'sp4_v_t_46')
// (15, 3, 'lutff_7/out')
// (15, 3, 'sp12_v_b_14')
// (15, 3, 'sp4_h_r_14')
// (15, 3, 'sp4_h_r_46')
// (15, 3, 'sp4_v_b_46')
// (15, 4, 'neigh_op_bot_7')
// (15, 4, 'sp12_v_b_13')
// (15, 4, 'sp4_v_b_35')
// (15, 5, 'sp12_v_b_10')
// (15, 5, 'sp4_v_b_22')
// (15, 6, 'local_g0_3')
// (15, 6, 'lutff_6/in_1')
// (15, 6, 'sp12_v_b_9')
// (15, 6, 'sp4_v_b_11')
// (15, 7, 'sp12_v_b_6')
// (15, 8, 'local_g3_5')
// (15, 8, 'lutff_7/in_3')
// (15, 8, 'sp12_v_b_5')
// (15, 9, 'sp12_v_b_2')
// (15, 10, 'sp12_v_b_1')
// (16, 2, 'neigh_op_tnl_7')
// (16, 3, 'neigh_op_lft_7')
// (16, 3, 'sp4_h_l_46')
// (16, 3, 'sp4_h_r_27')
// (16, 4, 'neigh_op_bnl_7')
// (17, 3, 'sp4_h_r_38')
// (18, 3, 'sp4_h_l_38')

wire n1690;
// (12, 3, 'sp4_h_r_9')
// (13, 3, 'sp12_h_r_0')
// (13, 3, 'sp4_h_r_20')
// (14, 2, 'neigh_op_tnr_6')
// (14, 3, 'local_g1_3')
// (14, 3, 'lutff_global/cen')
// (14, 3, 'neigh_op_rgt_6')
// (14, 3, 'sp12_h_r_3')
// (14, 3, 'sp4_h_r_33')
// (14, 4, 'neigh_op_bnr_6')
// (15, 1, 'sp4_r_v_b_27')
// (15, 2, 'neigh_op_top_6')
// (15, 2, 'sp4_r_v_b_14')
// (15, 3, 'lutff_6/out')
// (15, 3, 'sp12_h_r_4')
// (15, 3, 'sp4_h_r_44')
// (15, 3, 'sp4_r_v_b_3')
// (15, 4, 'neigh_op_bot_6')
// (16, 0, 'span4_vert_27')
// (16, 1, 'sp4_v_b_27')
// (16, 2, 'neigh_op_tnl_6')
// (16, 2, 'sp4_v_b_14')
// (16, 3, 'local_g1_3')
// (16, 3, 'lutff_global/cen')
// (16, 3, 'neigh_op_lft_6')
// (16, 3, 'sp12_h_r_7')
// (16, 3, 'sp4_h_l_44')
// (16, 3, 'sp4_v_b_3')
// (16, 4, 'neigh_op_bnl_6')
// (17, 3, 'sp12_h_r_8')
// (18, 3, 'sp12_h_r_11')
// (19, 3, 'sp12_h_r_12')
// (20, 3, 'sp12_h_r_15')
// (21, 3, 'sp12_h_r_16')
// (22, 3, 'sp12_h_r_19')
// (23, 3, 'sp12_h_r_20')
// (24, 3, 'sp12_h_r_23')
// (25, 3, 'sp12_h_l_23')

reg n1691 = 0;
// (12, 3, 'sp4_r_v_b_37')
// (12, 4, 'sp4_r_v_b_24')
// (12, 5, 'sp4_r_v_b_13')
// (12, 6, 'sp4_r_v_b_0')
// (12, 7, 'sp4_r_v_b_37')
// (12, 8, 'sp4_r_v_b_24')
// (12, 9, 'sp4_r_v_b_13')
// (12, 10, 'sp4_r_v_b_0')
// (13, 2, 'sp4_h_r_0')
// (13, 2, 'sp4_v_t_37')
// (13, 3, 'local_g2_5')
// (13, 3, 'lutff_0/in_1')
// (13, 3, 'sp4_v_b_37')
// (13, 4, 'sp4_v_b_24')
// (13, 5, 'sp4_v_b_13')
// (13, 6, 'sp4_v_b_0')
// (13, 6, 'sp4_v_t_37')
// (13, 7, 'local_g2_5')
// (13, 7, 'lutff_5/in_2')
// (13, 7, 'lutff_7/in_2')
// (13, 7, 'sp4_v_b_37')
// (13, 8, 'sp4_v_b_24')
// (13, 9, 'sp4_v_b_13')
// (13, 10, 'sp4_v_b_0')
// (14, 1, 'neigh_op_tnr_4')
// (14, 2, 'neigh_op_rgt_4')
// (14, 2, 'sp4_h_r_13')
// (14, 2, 'sp4_r_v_b_40')
// (14, 3, 'neigh_op_bnr_4')
// (14, 3, 'sp4_r_v_b_29')
// (14, 4, 'sp4_r_v_b_16')
// (14, 5, 'sp4_r_v_b_5')
// (14, 6, 'sp4_r_v_b_45')
// (14, 7, 'sp4_r_v_b_32')
// (14, 8, 'sp4_r_v_b_21')
// (14, 9, 'sp4_r_v_b_8')
// (15, 1, 'neigh_op_top_4')
// (15, 1, 'sp4_v_t_40')
// (15, 2, 'lutff_4/out')
// (15, 2, 'sp4_h_r_24')
// (15, 2, 'sp4_v_b_40')
// (15, 3, 'neigh_op_bot_4')
// (15, 3, 'sp4_v_b_29')
// (15, 4, 'sp4_v_b_16')
// (15, 5, 'local_g0_5')
// (15, 5, 'lutff_2/in_3')
// (15, 5, 'sp4_v_b_5')
// (15, 5, 'sp4_v_t_45')
// (15, 6, 'sp4_v_b_45')
// (15, 7, 'local_g3_0')
// (15, 7, 'lutff_4/in_1')
// (15, 7, 'sp4_v_b_32')
// (15, 8, 'sp4_v_b_21')
// (15, 9, 'sp4_v_b_8')
// (16, 1, 'neigh_op_tnl_4')
// (16, 2, 'neigh_op_lft_4')
// (16, 2, 'sp4_h_r_37')
// (16, 3, 'neigh_op_bnl_4')
// (17, 2, 'sp4_h_l_37')

reg n1692 = 0;
// (12, 3, 'sp4_r_v_b_42')
// (12, 4, 'local_g0_7')
// (12, 4, 'lutff_5/in_0')
// (12, 4, 'sp4_r_v_b_31')
// (12, 5, 'sp4_r_v_b_18')
// (12, 6, 'sp4_r_v_b_7')
// (13, 2, 'sp4_v_t_42')
// (13, 3, 'sp4_v_b_42')
// (13, 4, 'sp4_v_b_31')
// (13, 5, 'sp4_v_b_18')
// (13, 6, 'sp4_h_r_7')
// (13, 6, 'sp4_v_b_7')
// (13, 7, 'sp4_r_v_b_39')
// (13, 8, 'sp4_r_v_b_26')
// (13, 9, 'sp4_r_v_b_15')
// (13, 10, 'sp4_r_v_b_2')
// (14, 6, 'sp4_h_r_18')
// (14, 6, 'sp4_h_r_2')
// (14, 6, 'sp4_v_t_39')
// (14, 7, 'local_g2_7')
// (14, 7, 'lutff_0/in_3')
// (14, 7, 'lutff_1/in_2')
// (14, 7, 'sp4_v_b_39')
// (14, 8, 'sp4_v_b_26')
// (14, 9, 'sp4_v_b_15')
// (14, 10, 'sp4_v_b_2')
// (15, 5, 'neigh_op_tnr_5')
// (15, 6, 'neigh_op_rgt_5')
// (15, 6, 'sp4_h_r_15')
// (15, 6, 'sp4_h_r_31')
// (15, 7, 'local_g0_5')
// (15, 7, 'lutff_6/in_3')
// (15, 7, 'neigh_op_bnr_5')
// (16, 5, 'neigh_op_top_5')
// (16, 6, 'lutff_5/out')
// (16, 6, 'sp4_h_r_26')
// (16, 6, 'sp4_h_r_42')
// (16, 7, 'local_g1_5')
// (16, 7, 'lutff_7/in_3')
// (16, 7, 'neigh_op_bot_5')
// (17, 5, 'neigh_op_tnl_5')
// (17, 6, 'neigh_op_lft_5')
// (17, 6, 'sp4_h_l_42')
// (17, 6, 'sp4_h_r_39')
// (17, 7, 'neigh_op_bnl_5')
// (18, 6, 'sp4_h_l_39')

wire n1693;
// (12, 4, 'neigh_op_tnr_0')
// (12, 5, 'neigh_op_rgt_0')
// (12, 6, 'neigh_op_bnr_0')
// (13, 4, 'neigh_op_top_0')
// (13, 5, 'local_g0_0')
// (13, 5, 'lutff_0/out')
// (13, 5, 'lutff_2/in_0')
// (13, 6, 'neigh_op_bot_0')
// (14, 4, 'neigh_op_tnl_0')
// (14, 5, 'neigh_op_lft_0')
// (14, 6, 'neigh_op_bnl_0')

reg n1694 = 0;
// (12, 4, 'neigh_op_tnr_1')
// (12, 5, 'local_g2_1')
// (12, 5, 'lutff_6/in_3')
// (12, 5, 'neigh_op_rgt_1')
// (12, 6, 'neigh_op_bnr_1')
// (13, 4, 'neigh_op_top_1')
// (13, 5, 'lutff_1/out')
// (13, 6, 'local_g0_1')
// (13, 6, 'lutff_3/in_2')
// (13, 6, 'lutff_5/in_2')
// (13, 6, 'neigh_op_bot_1')
// (14, 4, 'neigh_op_tnl_1')
// (14, 5, 'neigh_op_lft_1')
// (14, 6, 'neigh_op_bnl_1')

wire n1695;
// (12, 4, 'neigh_op_tnr_4')
// (12, 5, 'neigh_op_rgt_4')
// (12, 6, 'local_g1_4')
// (12, 6, 'lutff_1/in_2')
// (12, 6, 'neigh_op_bnr_4')
// (13, 4, 'neigh_op_top_4')
// (13, 5, 'lutff_4/out')
// (13, 6, 'neigh_op_bot_4')
// (14, 4, 'neigh_op_tnl_4')
// (14, 5, 'neigh_op_lft_4')
// (14, 6, 'neigh_op_bnl_4')

reg n1696 = 0;
// (12, 4, 'neigh_op_tnr_5')
// (12, 5, 'neigh_op_rgt_5')
// (12, 6, 'neigh_op_bnr_5')
// (13, 4, 'neigh_op_top_5')
// (13, 5, 'local_g3_5')
// (13, 5, 'lutff_0/in_2')
// (13, 5, 'lutff_5/out')
// (13, 6, 'local_g1_5')
// (13, 6, 'lutff_2/in_2')
// (13, 6, 'lutff_6/in_0')
// (13, 6, 'neigh_op_bot_5')
// (14, 4, 'neigh_op_tnl_5')
// (14, 5, 'neigh_op_lft_5')
// (14, 6, 'neigh_op_bnl_5')

wire n1697;
// (12, 4, 'neigh_op_tnr_6')
// (12, 5, 'neigh_op_rgt_6')
// (12, 6, 'local_g0_6')
// (12, 6, 'lutff_0/in_2')
// (12, 6, 'neigh_op_bnr_6')
// (13, 4, 'neigh_op_top_6')
// (13, 5, 'lutff_6/out')
// (13, 6, 'neigh_op_bot_6')
// (14, 4, 'neigh_op_tnl_6')
// (14, 5, 'neigh_op_lft_6')
// (14, 6, 'neigh_op_bnl_6')

reg n1698 = 0;
// (12, 4, 'neigh_op_tnr_7')
// (12, 5, 'neigh_op_rgt_7')
// (12, 6, 'local_g1_7')
// (12, 6, 'lutff_4/in_2')
// (12, 6, 'neigh_op_bnr_7')
// (13, 4, 'neigh_op_top_7')
// (13, 5, 'lutff_7/out')
// (13, 5, 'sp4_r_v_b_47')
// (13, 6, 'neigh_op_bot_7')
// (13, 6, 'sp4_r_v_b_34')
// (13, 7, 'sp4_r_v_b_23')
// (13, 8, 'sp4_r_v_b_10')
// (14, 4, 'local_g2_7')
// (14, 4, 'lutff_2/in_3')
// (14, 4, 'neigh_op_tnl_7')
// (14, 4, 'sp4_v_t_47')
// (14, 5, 'neigh_op_lft_7')
// (14, 5, 'sp4_v_b_47')
// (14, 6, 'neigh_op_bnl_7')
// (14, 6, 'sp4_v_b_34')
// (14, 7, 'sp4_v_b_23')
// (14, 8, 'sp4_h_r_10')
// (14, 8, 'sp4_v_b_10')
// (15, 8, 'local_g0_7')
// (15, 8, 'lutff_3/in_0')
// (15, 8, 'sp4_h_r_23')
// (16, 8, 'sp4_h_r_34')
// (17, 8, 'sp4_h_r_47')
// (18, 8, 'sp4_h_l_47')

reg n1699 = 0;
// (12, 4, 'sp4_h_r_1')
// (12, 7, 'sp4_h_r_0')
// (12, 9, 'sp4_h_r_4')
// (13, 4, 'local_g1_4')
// (13, 4, 'lutff_0/in_1')
// (13, 4, 'sp4_h_r_12')
// (13, 7, 'local_g0_5')
// (13, 7, 'lutff_2/in_3')
// (13, 7, 'sp4_h_r_13')
// (13, 9, 'local_g1_1')
// (13, 9, 'lutff_6/in_2')
// (13, 9, 'sp4_h_r_17')
// (14, 2, 'sp4_r_v_b_44')
// (14, 3, 'neigh_op_tnr_2')
// (14, 3, 'sp4_r_v_b_33')
// (14, 4, 'neigh_op_rgt_2')
// (14, 4, 'sp4_h_r_25')
// (14, 4, 'sp4_r_v_b_20')
// (14, 5, 'neigh_op_bnr_2')
// (14, 5, 'sp4_r_v_b_9')
// (14, 6, 'sp4_r_v_b_37')
// (14, 7, 'sp4_h_r_24')
// (14, 7, 'sp4_r_v_b_24')
// (14, 8, 'sp4_r_v_b_13')
// (14, 9, 'sp4_h_r_28')
// (14, 9, 'sp4_r_v_b_0')
// (15, 1, 'sp4_v_t_44')
// (15, 2, 'sp4_r_v_b_45')
// (15, 2, 'sp4_v_b_44')
// (15, 3, 'neigh_op_top_2')
// (15, 3, 'sp4_r_v_b_32')
// (15, 3, 'sp4_v_b_33')
// (15, 4, 'lutff_2/out')
// (15, 4, 'sp4_h_r_36')
// (15, 4, 'sp4_r_v_b_21')
// (15, 4, 'sp4_r_v_b_37')
// (15, 4, 'sp4_v_b_20')
// (15, 5, 'neigh_op_bot_2')
// (15, 5, 'sp4_r_v_b_24')
// (15, 5, 'sp4_r_v_b_8')
// (15, 5, 'sp4_v_b_9')
// (15, 5, 'sp4_v_t_37')
// (15, 6, 'sp4_r_v_b_13')
// (15, 6, 'sp4_r_v_b_41')
// (15, 6, 'sp4_v_b_37')
// (15, 7, 'local_g1_0')
// (15, 7, 'lutff_3/in_0')
// (15, 7, 'sp4_h_r_37')
// (15, 7, 'sp4_r_v_b_0')
// (15, 7, 'sp4_r_v_b_28')
// (15, 7, 'sp4_v_b_24')
// (15, 8, 'sp4_r_v_b_17')
// (15, 8, 'sp4_v_b_13')
// (15, 9, 'local_g0_0')
// (15, 9, 'lutff_0/in_2')
// (15, 9, 'sp4_h_r_41')
// (15, 9, 'sp4_r_v_b_4')
// (15, 9, 'sp4_v_b_0')
// (16, 1, 'sp4_v_t_45')
// (16, 2, 'sp4_v_b_45')
// (16, 3, 'neigh_op_tnl_2')
// (16, 3, 'sp4_v_b_32')
// (16, 3, 'sp4_v_t_37')
// (16, 4, 'neigh_op_lft_2')
// (16, 4, 'sp4_h_l_36')
// (16, 4, 'sp4_v_b_21')
// (16, 4, 'sp4_v_b_37')
// (16, 5, 'neigh_op_bnl_2')
// (16, 5, 'sp4_v_b_24')
// (16, 5, 'sp4_v_b_8')
// (16, 5, 'sp4_v_t_41')
// (16, 6, 'sp4_v_b_13')
// (16, 6, 'sp4_v_b_41')
// (16, 7, 'sp4_h_l_37')
// (16, 7, 'sp4_v_b_0')
// (16, 7, 'sp4_v_b_28')
// (16, 8, 'sp4_v_b_17')
// (16, 9, 'sp4_h_l_41')
// (16, 9, 'sp4_v_b_4')

reg n1700 = 0;
// (12, 4, 'sp4_h_r_3')
// (13, 4, 'sp4_h_r_14')
// (13, 8, 'sp4_h_r_2')
// (14, 4, 'local_g3_3')
// (14, 4, 'lutff_6/in_0')
// (14, 4, 'sp4_h_r_27')
// (14, 8, 'local_g1_7')
// (14, 8, 'lutff_7/in_1')
// (14, 8, 'sp4_h_r_15')
// (15, 2, 'sp4_r_v_b_43')
// (15, 3, 'sp4_r_v_b_30')
// (15, 4, 'neigh_op_tnr_3')
// (15, 4, 'sp4_h_r_38')
// (15, 4, 'sp4_r_v_b_19')
// (15, 5, 'neigh_op_rgt_3')
// (15, 5, 'sp4_r_v_b_38')
// (15, 5, 'sp4_r_v_b_6')
// (15, 6, 'neigh_op_bnr_3')
// (15, 6, 'sp4_r_v_b_27')
// (15, 6, 'sp4_r_v_b_44')
// (15, 7, 'sp4_r_v_b_14')
// (15, 7, 'sp4_r_v_b_33')
// (15, 8, 'sp4_h_r_26')
// (15, 8, 'sp4_r_v_b_20')
// (15, 8, 'sp4_r_v_b_3')
// (15, 9, 'local_g2_1')
// (15, 9, 'lutff_7/in_0')
// (15, 9, 'sp4_r_v_b_9')
// (16, 1, 'sp4_v_t_43')
// (16, 2, 'sp4_v_b_43')
// (16, 3, 'sp4_v_b_30')
// (16, 4, 'neigh_op_top_3')
// (16, 4, 'sp4_h_l_38')
// (16, 4, 'sp4_v_b_19')
// (16, 4, 'sp4_v_t_38')
// (16, 5, 'local_g2_3')
// (16, 5, 'lutff_3/out')
// (16, 5, 'lutff_7/in_0')
// (16, 5, 'sp4_r_v_b_39')
// (16, 5, 'sp4_v_b_38')
// (16, 5, 'sp4_v_b_6')
// (16, 5, 'sp4_v_t_44')
// (16, 6, 'neigh_op_bot_3')
// (16, 6, 'sp4_r_v_b_26')
// (16, 6, 'sp4_v_b_27')
// (16, 6, 'sp4_v_b_44')
// (16, 7, 'sp4_r_v_b_15')
// (16, 7, 'sp4_v_b_14')
// (16, 7, 'sp4_v_b_33')
// (16, 8, 'local_g1_3')
// (16, 8, 'lutff_1/in_1')
// (16, 8, 'sp4_h_r_39')
// (16, 8, 'sp4_r_v_b_2')
// (16, 8, 'sp4_v_b_20')
// (16, 8, 'sp4_v_b_3')
// (16, 9, 'sp4_v_b_9')
// (17, 4, 'neigh_op_tnl_3')
// (17, 4, 'sp4_v_t_39')
// (17, 5, 'neigh_op_lft_3')
// (17, 5, 'sp4_v_b_39')
// (17, 6, 'neigh_op_bnl_3')
// (17, 6, 'sp4_v_b_26')
// (17, 7, 'sp4_v_b_15')
// (17, 8, 'sp4_h_l_39')
// (17, 8, 'sp4_v_b_2')

reg n1701 = 0;
// (12, 4, 'sp4_r_v_b_37')
// (12, 5, 'sp4_r_v_b_24')
// (12, 6, 'sp4_r_v_b_13')
// (12, 7, 'sp4_r_v_b_0')
// (12, 8, 'sp4_r_v_b_37')
// (12, 9, 'sp4_r_v_b_24')
// (12, 10, 'sp4_r_v_b_13')
// (12, 11, 'sp4_r_v_b_0')
// (13, 3, 'sp4_h_r_0')
// (13, 3, 'sp4_v_t_37')
// (13, 4, 'sp4_v_b_37')
// (13, 5, 'sp4_v_b_24')
// (13, 6, 'sp4_v_b_13')
// (13, 7, 'sp4_v_b_0')
// (13, 7, 'sp4_v_t_37')
// (13, 8, 'local_g3_5')
// (13, 8, 'lutff_3/in_1')
// (13, 8, 'sp4_v_b_37')
// (13, 9, 'sp4_v_b_24')
// (13, 10, 'sp4_v_b_13')
// (13, 11, 'sp4_v_b_0')
// (14, 2, 'neigh_op_tnr_4')
// (14, 3, 'neigh_op_rgt_4')
// (14, 3, 'sp4_h_r_13')
// (14, 4, 'neigh_op_bnr_4')
// (15, 2, 'local_g1_4')
// (15, 2, 'lutff_6/in_3')
// (15, 2, 'neigh_op_top_4')
// (15, 2, 'sp4_r_v_b_36')
// (15, 3, 'lutff_4/out')
// (15, 3, 'sp4_h_r_24')
// (15, 3, 'sp4_r_v_b_25')
// (15, 3, 'sp4_r_v_b_41')
// (15, 4, 'neigh_op_bot_4')
// (15, 4, 'sp4_r_v_b_12')
// (15, 4, 'sp4_r_v_b_28')
// (15, 5, 'local_g1_1')
// (15, 5, 'lutff_1/in_3')
// (15, 5, 'sp4_r_v_b_1')
// (15, 5, 'sp4_r_v_b_17')
// (15, 6, 'sp4_r_v_b_36')
// (15, 6, 'sp4_r_v_b_4')
// (15, 7, 'sp4_r_v_b_25')
// (15, 8, 'sp4_r_v_b_12')
// (15, 9, 'sp4_r_v_b_1')
// (16, 1, 'sp4_v_t_36')
// (16, 2, 'neigh_op_tnl_4')
// (16, 2, 'sp4_v_b_36')
// (16, 2, 'sp4_v_t_41')
// (16, 3, 'neigh_op_lft_4')
// (16, 3, 'sp4_h_r_37')
// (16, 3, 'sp4_v_b_25')
// (16, 3, 'sp4_v_b_41')
// (16, 4, 'neigh_op_bnl_4')
// (16, 4, 'sp4_v_b_12')
// (16, 4, 'sp4_v_b_28')
// (16, 5, 'sp4_v_b_1')
// (16, 5, 'sp4_v_b_17')
// (16, 5, 'sp4_v_t_36')
// (16, 6, 'local_g1_4')
// (16, 6, 'lutff_4/in_3')
// (16, 6, 'sp4_v_b_36')
// (16, 6, 'sp4_v_b_4')
// (16, 7, 'sp4_v_b_25')
// (16, 8, 'local_g0_4')
// (16, 8, 'lutff_6/in_2')
// (16, 8, 'sp4_v_b_12')
// (16, 9, 'sp4_v_b_1')
// (17, 3, 'sp4_h_l_37')

reg n1702 = 0;
// (12, 4, 'sp4_r_v_b_38')
// (12, 5, 'neigh_op_tnr_7')
// (12, 5, 'sp4_r_v_b_27')
// (12, 6, 'local_g2_7')
// (12, 6, 'lutff_3/in_2')
// (12, 6, 'neigh_op_rgt_7')
// (12, 6, 'sp4_r_v_b_14')
// (12, 6, 'sp4_r_v_b_46')
// (12, 7, 'neigh_op_bnr_7')
// (12, 7, 'sp4_r_v_b_3')
// (12, 7, 'sp4_r_v_b_35')
// (12, 8, 'sp4_r_v_b_22')
// (12, 9, 'sp4_r_v_b_11')
// (13, 3, 'sp4_v_t_38')
// (13, 4, 'sp4_v_b_38')
// (13, 5, 'neigh_op_top_7')
// (13, 5, 'sp4_v_b_27')
// (13, 5, 'sp4_v_t_46')
// (13, 6, 'lutff_7/out')
// (13, 6, 'sp4_r_v_b_47')
// (13, 6, 'sp4_v_b_14')
// (13, 6, 'sp4_v_b_46')
// (13, 7, 'neigh_op_bot_7')
// (13, 7, 'sp4_h_r_3')
// (13, 7, 'sp4_r_v_b_34')
// (13, 7, 'sp4_v_b_3')
// (13, 7, 'sp4_v_b_35')
// (13, 8, 'sp4_r_v_b_23')
// (13, 8, 'sp4_v_b_22')
// (13, 9, 'local_g2_2')
// (13, 9, 'lutff_3/in_1')
// (13, 9, 'sp4_h_r_11')
// (13, 9, 'sp4_r_v_b_10')
// (13, 9, 'sp4_v_b_11')
// (14, 5, 'neigh_op_tnl_7')
// (14, 5, 'sp4_v_t_47')
// (14, 6, 'neigh_op_lft_7')
// (14, 6, 'sp4_v_b_47')
// (14, 7, 'neigh_op_bnl_7')
// (14, 7, 'sp4_h_r_14')
// (14, 7, 'sp4_v_b_34')
// (14, 8, 'sp4_v_b_23')
// (14, 9, 'local_g1_2')
// (14, 9, 'lutff_0/in_1')
// (14, 9, 'sp4_h_r_22')
// (14, 9, 'sp4_v_b_10')
// (15, 7, 'local_g2_3')
// (15, 7, 'lutff_1/in_2')
// (15, 7, 'sp4_h_r_27')
// (15, 9, 'local_g2_3')
// (15, 9, 'lutff_2/in_1')
// (15, 9, 'sp4_h_r_35')
// (16, 7, 'sp4_h_r_38')
// (16, 9, 'sp4_h_r_46')
// (17, 7, 'sp4_h_l_38')
// (17, 9, 'sp4_h_l_46')

reg n1703 = 0;
// (12, 4, 'sp4_r_v_b_40')
// (12, 5, 'sp4_r_v_b_29')
// (12, 6, 'local_g3_0')
// (12, 6, 'lutff_5/in_0')
// (12, 6, 'sp4_r_v_b_16')
// (12, 7, 'local_g1_5')
// (12, 7, 'lutff_4/in_2')
// (12, 7, 'sp4_r_v_b_5')
// (13, 2, 'neigh_op_tnr_3')
// (13, 3, 'local_g2_3')
// (13, 3, 'lutff_6/in_3')
// (13, 3, 'neigh_op_rgt_3')
// (13, 3, 'sp4_h_r_11')
// (13, 3, 'sp4_v_t_40')
// (13, 4, 'neigh_op_bnr_3')
// (13, 4, 'sp4_v_b_40')
// (13, 5, 'sp4_v_b_29')
// (13, 6, 'sp4_v_b_16')
// (13, 7, 'sp4_v_b_5')
// (14, 2, 'neigh_op_top_3')
// (14, 3, 'lutff_3/out')
// (14, 3, 'sp4_h_r_22')
// (14, 4, 'neigh_op_bot_3')
// (15, 2, 'neigh_op_tnl_3')
// (15, 3, 'neigh_op_lft_3')
// (15, 3, 'sp4_h_r_35')
// (15, 4, 'neigh_op_bnl_3')
// (16, 3, 'sp4_h_r_46')
// (17, 3, 'sp4_h_l_46')

reg n1704 = 0;
// (12, 4, 'sp4_r_v_b_42')
// (12, 5, 'sp4_r_v_b_31')
// (12, 6, 'sp4_r_v_b_18')
// (12, 7, 'sp4_r_v_b_7')
// (13, 2, 'neigh_op_tnr_1')
// (13, 3, 'neigh_op_rgt_1')
// (13, 3, 'sp4_h_r_7')
// (13, 3, 'sp4_v_t_42')
// (13, 4, 'neigh_op_bnr_1')
// (13, 4, 'sp4_v_b_42')
// (13, 5, 'sp4_v_b_31')
// (13, 6, 'local_g1_2')
// (13, 6, 'lutff_2/in_3')
// (13, 6, 'lutff_6/in_1')
// (13, 6, 'sp4_v_b_18')
// (13, 7, 'sp4_v_b_7')
// (14, 1, 'sp4_r_v_b_27')
// (14, 2, 'neigh_op_top_1')
// (14, 2, 'sp4_r_v_b_14')
// (14, 3, 'lutff_1/out')
// (14, 3, 'sp4_h_r_18')
// (14, 3, 'sp4_r_v_b_3')
// (14, 4, 'neigh_op_bot_1')
// (15, 0, 'span4_vert_27')
// (15, 1, 'local_g3_3')
// (15, 1, 'lutff_4/in_0')
// (15, 1, 'sp4_v_b_27')
// (15, 2, 'neigh_op_tnl_1')
// (15, 2, 'sp4_v_b_14')
// (15, 3, 'neigh_op_lft_1')
// (15, 3, 'sp4_h_r_31')
// (15, 3, 'sp4_v_b_3')
// (15, 4, 'neigh_op_bnl_1')
// (16, 3, 'sp4_h_r_42')
// (17, 3, 'sp4_h_l_42')

reg n1705 = 0;
// (12, 4, 'sp4_r_v_b_43')
// (12, 5, 'sp4_r_v_b_30')
// (12, 6, 'sp4_r_v_b_19')
// (12, 6, 'sp4_r_v_b_39')
// (12, 7, 'sp4_r_v_b_26')
// (12, 7, 'sp4_r_v_b_6')
// (12, 8, 'sp4_r_v_b_15')
// (12, 8, 'sp4_r_v_b_47')
// (12, 9, 'sp4_r_v_b_2')
// (12, 9, 'sp4_r_v_b_34')
// (12, 10, 'neigh_op_tnr_5')
// (12, 10, 'sp4_r_v_b_23')
// (12, 10, 'sp4_r_v_b_39')
// (12, 11, 'neigh_op_rgt_5')
// (12, 11, 'sp4_r_v_b_10')
// (12, 11, 'sp4_r_v_b_26')
// (12, 12, 'neigh_op_bnr_5')
// (12, 12, 'sp4_r_v_b_15')
// (12, 13, 'sp4_r_v_b_2')
// (13, 3, 'sp4_v_t_43')
// (13, 4, 'sp4_v_b_43')
// (13, 5, 'sp4_v_b_30')
// (13, 5, 'sp4_v_t_39')
// (13, 6, 'local_g3_7')
// (13, 6, 'lutff_0/in_0')
// (13, 6, 'sp4_v_b_19')
// (13, 6, 'sp4_v_b_39')
// (13, 7, 'local_g0_6')
// (13, 7, 'lutff_7/in_3')
// (13, 7, 'sp4_h_r_10')
// (13, 7, 'sp4_v_b_26')
// (13, 7, 'sp4_v_b_6')
// (13, 7, 'sp4_v_t_47')
// (13, 8, 'sp4_v_b_15')
// (13, 8, 'sp4_v_b_47')
// (13, 9, 'sp4_v_b_2')
// (13, 9, 'sp4_v_b_34')
// (13, 9, 'sp4_v_t_39')
// (13, 10, 'neigh_op_top_5')
// (13, 10, 'sp4_v_b_23')
// (13, 10, 'sp4_v_b_39')
// (13, 11, 'lutff_5/out')
// (13, 11, 'sp4_h_r_10')
// (13, 11, 'sp4_v_b_10')
// (13, 11, 'sp4_v_b_26')
// (13, 12, 'neigh_op_bot_5')
// (13, 12, 'sp4_v_b_15')
// (13, 13, 'sp4_v_b_2')
// (14, 7, 'sp4_h_r_23')
// (14, 10, 'neigh_op_tnl_5')
// (14, 11, 'local_g1_5')
// (14, 11, 'lutff_5/in_1')
// (14, 11, 'lutff_7/in_3')
// (14, 11, 'neigh_op_lft_5')
// (14, 11, 'sp4_h_r_23')
// (14, 12, 'neigh_op_bnl_5')
// (15, 7, 'sp4_h_r_34')
// (15, 11, 'sp4_h_r_34')
// (16, 4, 'sp4_r_v_b_41')
// (16, 5, 'sp4_r_v_b_28')
// (16, 6, 'local_g3_1')
// (16, 6, 'lutff_7/in_1')
// (16, 6, 'sp4_r_v_b_17')
// (16, 7, 'sp4_h_r_47')
// (16, 7, 'sp4_r_v_b_4')
// (16, 11, 'local_g2_7')
// (16, 11, 'lutff_0/in_1')
// (16, 11, 'sp4_h_r_47')
// (17, 3, 'sp4_v_t_41')
// (17, 4, 'sp4_v_b_41')
// (17, 5, 'sp4_v_b_28')
// (17, 6, 'sp4_v_b_17')
// (17, 7, 'sp4_h_l_47')
// (17, 7, 'sp4_v_b_4')
// (17, 11, 'sp4_h_l_47')

reg n1706 = 0;
// (12, 4, 'sp4_r_v_b_46')
// (12, 5, 'sp4_r_v_b_35')
// (12, 6, 'sp4_r_v_b_22')
// (12, 7, 'sp4_r_v_b_11')
// (12, 8, 'sp4_r_v_b_46')
// (12, 9, 'neigh_op_tnr_3')
// (12, 9, 'sp4_r_v_b_35')
// (12, 10, 'neigh_op_rgt_3')
// (12, 10, 'sp4_r_v_b_22')
// (12, 10, 'sp4_r_v_b_38')
// (12, 11, 'neigh_op_bnr_3')
// (12, 11, 'sp4_r_v_b_11')
// (12, 11, 'sp4_r_v_b_27')
// (12, 12, 'sp4_r_v_b_14')
// (12, 13, 'sp4_r_v_b_3')
// (13, 3, 'sp4_v_t_46')
// (13, 4, 'sp4_v_b_46')
// (13, 5, 'sp4_v_b_35')
// (13, 6, 'local_g0_6')
// (13, 6, 'lutff_6/in_2')
// (13, 6, 'sp4_v_b_22')
// (13, 7, 'local_g3_2')
// (13, 7, 'lutff_5/in_0')
// (13, 7, 'sp4_r_v_b_42')
// (13, 7, 'sp4_v_b_11')
// (13, 7, 'sp4_v_t_46')
// (13, 8, 'sp4_r_v_b_31')
// (13, 8, 'sp4_v_b_46')
// (13, 9, 'neigh_op_top_3')
// (13, 9, 'sp4_r_v_b_18')
// (13, 9, 'sp4_v_b_35')
// (13, 9, 'sp4_v_t_38')
// (13, 10, 'local_g1_3')
// (13, 10, 'lutff_0/in_0')
// (13, 10, 'lutff_3/out')
// (13, 10, 'sp4_r_v_b_7')
// (13, 10, 'sp4_v_b_22')
// (13, 10, 'sp4_v_b_38')
// (13, 11, 'neigh_op_bot_3')
// (13, 11, 'sp4_v_b_11')
// (13, 11, 'sp4_v_b_27')
// (13, 12, 'local_g1_6')
// (13, 12, 'lutff_1/in_2')
// (13, 12, 'sp4_v_b_14')
// (13, 13, 'sp4_v_b_3')
// (14, 6, 'sp4_v_t_42')
// (14, 7, 'sp4_v_b_42')
// (14, 8, 'sp4_v_b_31')
// (14, 9, 'neigh_op_tnl_3')
// (14, 9, 'sp4_v_b_18')
// (14, 10, 'neigh_op_lft_3')
// (14, 10, 'sp4_v_b_7')
// (14, 11, 'neigh_op_bnl_3')

wire n1707;
// (12, 5, 'neigh_op_tnr_0')
// (12, 6, 'neigh_op_rgt_0')
// (12, 7, 'neigh_op_bnr_0')
// (13, 5, 'neigh_op_top_0')
// (13, 6, 'local_g2_0')
// (13, 6, 'lutff_0/out')
// (13, 6, 'lutff_4/in_0')
// (13, 7, 'neigh_op_bot_0')
// (14, 5, 'neigh_op_tnl_0')
// (14, 6, 'neigh_op_lft_0')
// (14, 7, 'neigh_op_bnl_0')

wire n1708;
// (12, 5, 'neigh_op_tnr_1')
// (12, 6, 'neigh_op_rgt_1')
// (12, 7, 'neigh_op_bnr_1')
// (13, 5, 'neigh_op_top_1')
// (13, 6, 'lutff_1/out')
// (13, 7, 'local_g1_1')
// (13, 7, 'lutff_4/in_0')
// (13, 7, 'neigh_op_bot_1')
// (14, 5, 'neigh_op_tnl_1')
// (14, 6, 'neigh_op_lft_1')
// (14, 7, 'neigh_op_bnl_1')

wire n1709;
// (12, 5, 'neigh_op_tnr_2')
// (12, 6, 'neigh_op_rgt_2')
// (12, 7, 'neigh_op_bnr_2')
// (13, 5, 'neigh_op_top_2')
// (13, 6, 'local_g0_2')
// (13, 6, 'lutff_2/out')
// (13, 6, 'lutff_4/in_2')
// (13, 7, 'neigh_op_bot_2')
// (14, 5, 'neigh_op_tnl_2')
// (14, 6, 'neigh_op_lft_2')
// (14, 7, 'neigh_op_bnl_2')

wire n1710;
// (12, 5, 'neigh_op_tnr_3')
// (12, 6, 'neigh_op_rgt_3')
// (12, 7, 'local_g1_3')
// (12, 7, 'lutff_0/in_0')
// (12, 7, 'neigh_op_bnr_3')
// (13, 5, 'neigh_op_top_3')
// (13, 6, 'lutff_3/out')
// (13, 7, 'neigh_op_bot_3')
// (14, 5, 'neigh_op_tnl_3')
// (14, 6, 'neigh_op_lft_3')
// (14, 7, 'neigh_op_bnl_3')

wire n1711;
// (12, 5, 'neigh_op_tnr_4')
// (12, 6, 'neigh_op_rgt_4')
// (12, 7, 'neigh_op_bnr_4')
// (13, 5, 'neigh_op_top_4')
// (13, 6, 'lutff_4/out')
// (13, 6, 'sp4_r_v_b_41')
// (13, 7, 'neigh_op_bot_4')
// (13, 7, 'sp4_r_v_b_28')
// (13, 8, 'sp4_r_v_b_17')
// (13, 9, 'local_g1_4')
// (13, 9, 'lutff_0/in_1')
// (13, 9, 'sp4_r_v_b_4')
// (14, 5, 'neigh_op_tnl_4')
// (14, 5, 'sp4_v_t_41')
// (14, 6, 'neigh_op_lft_4')
// (14, 6, 'sp4_v_b_41')
// (14, 7, 'neigh_op_bnl_4')
// (14, 7, 'sp4_v_b_28')
// (14, 8, 'sp4_v_b_17')
// (14, 9, 'sp4_v_b_4')

wire n1712;
// (12, 5, 'neigh_op_tnr_5')
// (12, 6, 'neigh_op_rgt_5')
// (12, 7, 'neigh_op_bnr_5')
// (13, 5, 'neigh_op_top_5')
// (13, 6, 'local_g2_5')
// (13, 6, 'lutff_4/in_1')
// (13, 6, 'lutff_5/out')
// (13, 7, 'neigh_op_bot_5')
// (14, 5, 'neigh_op_tnl_5')
// (14, 6, 'neigh_op_lft_5')
// (14, 7, 'neigh_op_bnl_5')

wire n1713;
// (12, 5, 'neigh_op_tnr_6')
// (12, 6, 'neigh_op_rgt_6')
// (12, 7, 'local_g0_6')
// (12, 7, 'lutff_0/in_2')
// (12, 7, 'neigh_op_bnr_6')
// (13, 5, 'neigh_op_top_6')
// (13, 6, 'lutff_6/out')
// (13, 7, 'neigh_op_bot_6')
// (14, 5, 'neigh_op_tnl_6')
// (14, 6, 'neigh_op_lft_6')
// (14, 7, 'neigh_op_bnl_6')

reg n1714 = 0;
// (12, 5, 'sp4_h_r_9')
// (13, 5, 'local_g1_4')
// (13, 5, 'lutff_3/in_0')
// (13, 5, 'sp4_h_r_20')
// (14, 3, 'sp4_r_v_b_36')
// (14, 4, 'neigh_op_tnr_6')
// (14, 4, 'sp4_r_v_b_25')
// (14, 4, 'sp4_r_v_b_41')
// (14, 5, 'neigh_op_rgt_6')
// (14, 5, 'sp4_h_r_33')
// (14, 5, 'sp4_r_v_b_12')
// (14, 5, 'sp4_r_v_b_28')
// (14, 6, 'local_g0_6')
// (14, 6, 'lutff_4/in_2')
// (14, 6, 'neigh_op_bnr_6')
// (14, 6, 'sp4_r_v_b_1')
// (14, 6, 'sp4_r_v_b_17')
// (14, 7, 'sp4_r_v_b_4')
// (14, 7, 'sp4_r_v_b_41')
// (14, 8, 'sp4_r_v_b_28')
// (14, 8, 'sp4_r_v_b_42')
// (14, 9, 'sp4_r_v_b_17')
// (14, 9, 'sp4_r_v_b_31')
// (14, 10, 'local_g1_4')
// (14, 10, 'lutff_7/in_0')
// (14, 10, 'sp4_r_v_b_18')
// (14, 10, 'sp4_r_v_b_4')
// (14, 11, 'sp4_r_v_b_7')
// (15, 2, 'sp4_v_t_36')
// (15, 3, 'sp4_v_b_36')
// (15, 3, 'sp4_v_t_41')
// (15, 4, 'neigh_op_top_6')
// (15, 4, 'sp4_v_b_25')
// (15, 4, 'sp4_v_b_41')
// (15, 5, 'lutff_6/out')
// (15, 5, 'sp4_h_r_44')
// (15, 5, 'sp4_v_b_12')
// (15, 5, 'sp4_v_b_28')
// (15, 6, 'neigh_op_bot_6')
// (15, 6, 'sp4_r_v_b_39')
// (15, 6, 'sp4_v_b_1')
// (15, 6, 'sp4_v_b_17')
// (15, 6, 'sp4_v_t_41')
// (15, 7, 'sp4_r_v_b_26')
// (15, 7, 'sp4_v_b_4')
// (15, 7, 'sp4_v_b_41')
// (15, 7, 'sp4_v_t_42')
// (15, 8, 'sp4_r_v_b_15')
// (15, 8, 'sp4_v_b_28')
// (15, 8, 'sp4_v_b_42')
// (15, 9, 'local_g1_2')
// (15, 9, 'lutff_1/in_0')
// (15, 9, 'sp4_r_v_b_2')
// (15, 9, 'sp4_v_b_17')
// (15, 9, 'sp4_v_b_31')
// (15, 10, 'local_g0_2')
// (15, 10, 'lutff_7/in_1')
// (15, 10, 'sp4_v_b_18')
// (15, 10, 'sp4_v_b_4')
// (15, 11, 'sp4_v_b_7')
// (16, 4, 'neigh_op_tnl_6')
// (16, 5, 'neigh_op_lft_6')
// (16, 5, 'sp4_h_l_44')
// (16, 5, 'sp4_v_t_39')
// (16, 6, 'neigh_op_bnl_6')
// (16, 6, 'sp4_v_b_39')
// (16, 7, 'sp4_v_b_26')
// (16, 8, 'sp4_v_b_15')
// (16, 9, 'sp4_v_b_2')

reg n1715 = 0;
// (12, 5, 'sp4_r_v_b_40')
// (12, 6, 'sp4_r_v_b_29')
// (12, 7, 'sp4_r_v_b_16')
// (12, 8, 'sp4_r_v_b_5')
// (12, 9, 'sp4_r_v_b_39')
// (12, 10, 'sp4_r_v_b_26')
// (12, 11, 'sp4_r_v_b_15')
// (12, 12, 'sp4_r_v_b_2')
// (12, 13, 'sp4_r_v_b_43')
// (12, 14, 'sp4_r_v_b_30')
// (12, 15, 'sp4_r_v_b_19')
// (12, 16, 'sp4_r_v_b_6')
// (12, 17, 'sp4_r_v_b_38')
// (12, 18, 'neigh_op_tnr_7')
// (12, 18, 'sp4_r_v_b_27')
// (12, 19, 'neigh_op_rgt_7')
// (12, 19, 'sp4_r_v_b_14')
// (12, 20, 'neigh_op_bnr_7')
// (12, 20, 'sp4_r_v_b_3')
// (13, 4, 'local_g0_5')
// (13, 4, 'lutff_0/in_3')
// (13, 4, 'sp4_h_r_5')
// (13, 4, 'sp4_v_t_40')
// (13, 5, 'sp4_v_b_40')
// (13, 6, 'sp4_v_b_29')
// (13, 7, 'sp4_v_b_16')
// (13, 8, 'sp4_v_b_5')
// (13, 8, 'sp4_v_t_39')
// (13, 9, 'sp4_v_b_39')
// (13, 10, 'sp4_v_b_26')
// (13, 11, 'sp4_v_b_15')
// (13, 12, 'sp4_v_b_2')
// (13, 12, 'sp4_v_t_43')
// (13, 13, 'sp4_v_b_43')
// (13, 14, 'sp4_v_b_30')
// (13, 15, 'sp4_v_b_19')
// (13, 16, 'sp4_v_b_6')
// (13, 16, 'sp4_v_t_38')
// (13, 17, 'sp4_v_b_38')
// (13, 18, 'local_g0_7')
// (13, 18, 'lutff_5/in_0')
// (13, 18, 'neigh_op_top_7')
// (13, 18, 'sp4_v_b_27')
// (13, 19, 'local_g0_7')
// (13, 19, 'lutff_4/in_1')
// (13, 19, 'lutff_7/out')
// (13, 19, 'sp4_v_b_14')
// (13, 20, 'local_g1_7')
// (13, 20, 'lutff_4/in_2')
// (13, 20, 'neigh_op_bot_7')
// (13, 20, 'sp4_v_b_3')
// (14, 4, 'sp4_h_r_16')
// (14, 18, 'neigh_op_tnl_7')
// (14, 19, 'neigh_op_lft_7')
// (14, 20, 'neigh_op_bnl_7')
// (15, 4, 'sp4_h_r_29')
// (16, 4, 'sp4_h_r_40')
// (17, 4, 'sp4_h_l_40')

reg n1716 = 0;
// (12, 5, 'sp4_r_v_b_45')
// (12, 6, 'sp4_r_v_b_32')
// (12, 7, 'sp4_r_v_b_21')
// (12, 8, 'sp4_r_v_b_8')
// (13, 3, 'local_g3_5')
// (13, 3, 'lutff_6/in_2')
// (13, 3, 'sp4_r_v_b_45')
// (13, 4, 'sp4_h_r_8')
// (13, 4, 'sp4_r_v_b_32')
// (13, 4, 'sp4_v_t_45')
// (13, 5, 'sp4_r_v_b_21')
// (13, 5, 'sp4_v_b_45')
// (13, 6, 'sp4_r_v_b_8')
// (13, 6, 'sp4_v_b_32')
// (13, 7, 'local_g1_5')
// (13, 7, 'lutff_4/in_2')
// (13, 7, 'sp4_v_b_21')
// (13, 8, 'sp4_v_b_8')
// (14, 2, 'sp4_h_r_2')
// (14, 2, 'sp4_v_t_45')
// (14, 3, 'sp4_v_b_45')
// (14, 4, 'sp4_h_r_21')
// (14, 4, 'sp4_v_b_32')
// (14, 5, 'sp4_v_b_21')
// (14, 6, 'local_g0_0')
// (14, 6, 'lutff_1/in_1')
// (14, 6, 'sp4_v_b_8')
// (15, 1, 'neigh_op_tnr_5')
// (15, 2, 'neigh_op_rgt_5')
// (15, 2, 'sp4_h_r_15')
// (15, 3, 'neigh_op_bnr_5')
// (15, 4, 'sp4_h_r_32')
// (16, 0, 'span12_vert_13')
// (16, 1, 'neigh_op_top_5')
// (16, 1, 'sp12_v_b_13')
// (16, 1, 'sp4_r_v_b_38')
// (16, 2, 'lutff_5/out')
// (16, 2, 'sp12_v_b_10')
// (16, 2, 'sp4_h_r_26')
// (16, 2, 'sp4_r_v_b_27')
// (16, 3, 'neigh_op_bot_5')
// (16, 3, 'sp12_v_b_9')
// (16, 3, 'sp4_r_v_b_14')
// (16, 4, 'sp12_v_b_6')
// (16, 4, 'sp4_h_r_45')
// (16, 4, 'sp4_r_v_b_3')
// (16, 5, 'sp12_v_b_5')
// (16, 6, 'sp12_v_b_2')
// (16, 7, 'local_g2_1')
// (16, 7, 'lutff_0/in_3')
// (16, 7, 'sp12_v_b_1')
// (17, 0, 'span4_vert_38')
// (17, 1, 'neigh_op_tnl_5')
// (17, 1, 'sp4_v_b_38')
// (17, 2, 'neigh_op_lft_5')
// (17, 2, 'sp4_h_r_39')
// (17, 2, 'sp4_v_b_27')
// (17, 3, 'neigh_op_bnl_5')
// (17, 3, 'sp4_v_b_14')
// (17, 4, 'sp4_h_l_45')
// (17, 4, 'sp4_v_b_3')
// (18, 2, 'sp4_h_l_39')

wire n1717;
// (12, 6, 'local_g2_6')
// (12, 6, 'lutff_4/in_0')
// (12, 6, 'sp4_r_v_b_38')
// (12, 7, 'neigh_op_tnr_7')
// (12, 7, 'sp4_r_v_b_27')
// (12, 8, 'neigh_op_rgt_7')
// (12, 8, 'sp4_r_v_b_14')
// (12, 9, 'neigh_op_bnr_7')
// (12, 9, 'sp4_r_v_b_3')
// (13, 5, 'sp4_v_t_38')
// (13, 6, 'sp4_v_b_38')
// (13, 7, 'neigh_op_top_7')
// (13, 7, 'sp4_v_b_27')
// (13, 8, 'lutff_7/out')
// (13, 8, 'sp4_v_b_14')
// (13, 9, 'neigh_op_bot_7')
// (13, 9, 'sp4_v_b_3')
// (14, 7, 'neigh_op_tnl_7')
// (14, 8, 'neigh_op_lft_7')
// (14, 9, 'neigh_op_bnl_7')

reg n1718 = 0;
// (12, 6, 'local_g3_1')
// (12, 6, 'lutff_2/in_2')
// (12, 6, 'sp4_r_v_b_41')
// (12, 7, 'sp4_r_v_b_28')
// (12, 8, 'neigh_op_tnr_2')
// (12, 8, 'sp4_r_v_b_17')
// (12, 9, 'neigh_op_rgt_2')
// (12, 9, 'sp4_r_v_b_36')
// (12, 9, 'sp4_r_v_b_4')
// (12, 10, 'neigh_op_bnr_2')
// (12, 10, 'sp4_r_v_b_25')
// (12, 11, 'sp4_r_v_b_12')
// (12, 12, 'sp4_r_v_b_1')
// (13, 5, 'sp4_v_t_41')
// (13, 6, 'sp4_r_v_b_40')
// (13, 6, 'sp4_v_b_41')
// (13, 7, 'sp4_r_v_b_29')
// (13, 7, 'sp4_v_b_28')
// (13, 8, 'neigh_op_top_2')
// (13, 8, 'sp4_r_v_b_16')
// (13, 8, 'sp4_v_b_17')
// (13, 8, 'sp4_v_t_36')
// (13, 9, 'lutff_2/out')
// (13, 9, 'sp4_r_v_b_5')
// (13, 9, 'sp4_v_b_36')
// (13, 9, 'sp4_v_b_4')
// (13, 10, 'neigh_op_bot_2')
// (13, 10, 'sp4_v_b_25')
// (13, 11, 'local_g0_4')
// (13, 11, 'lutff_4/in_0')
// (13, 11, 'sp4_v_b_12')
// (13, 12, 'local_g0_1')
// (13, 12, 'lutff_4/in_1')
// (13, 12, 'sp4_v_b_1')
// (14, 5, 'sp4_v_t_40')
// (14, 6, 'sp4_v_b_40')
// (14, 7, 'local_g2_5')
// (14, 7, 'lutff_1/in_0')
// (14, 7, 'sp4_v_b_29')
// (14, 8, 'neigh_op_tnl_2')
// (14, 8, 'sp4_v_b_16')
// (14, 9, 'neigh_op_lft_2')
// (14, 9, 'sp4_v_b_5')
// (14, 10, 'neigh_op_bnl_2')

wire n1719;
// (12, 6, 'neigh_op_tnr_0')
// (12, 7, 'neigh_op_rgt_0')
// (12, 8, 'neigh_op_bnr_0')
// (13, 6, 'neigh_op_top_0')
// (13, 7, 'local_g1_0')
// (13, 7, 'lutff_0/out')
// (13, 7, 'lutff_7/in_0')
// (13, 8, 'neigh_op_bot_0')
// (14, 6, 'neigh_op_tnl_0')
// (14, 7, 'neigh_op_lft_0')
// (14, 8, 'neigh_op_bnl_0')

wire n1720;
// (12, 6, 'neigh_op_tnr_2')
// (12, 7, 'neigh_op_rgt_2')
// (12, 8, 'neigh_op_bnr_2')
// (13, 6, 'neigh_op_top_2')
// (13, 7, 'local_g1_2')
// (13, 7, 'lutff_2/out')
// (13, 7, 'lutff_4/in_1')
// (13, 8, 'neigh_op_bot_2')
// (14, 6, 'neigh_op_tnl_2')
// (14, 7, 'neigh_op_lft_2')
// (14, 8, 'neigh_op_bnl_2')

wire n1721;
// (12, 6, 'neigh_op_tnr_3')
// (12, 7, 'neigh_op_rgt_3')
// (12, 8, 'neigh_op_bnr_3')
// (13, 6, 'neigh_op_top_3')
// (13, 7, 'lutff_3/out')
// (13, 8, 'local_g0_3')
// (13, 8, 'lutff_2/in_1')
// (13, 8, 'neigh_op_bot_3')
// (14, 6, 'neigh_op_tnl_3')
// (14, 7, 'neigh_op_lft_3')
// (14, 8, 'neigh_op_bnl_3')

wire n1722;
// (12, 6, 'neigh_op_tnr_4')
// (12, 7, 'neigh_op_rgt_4')
// (12, 8, 'neigh_op_bnr_4')
// (13, 6, 'neigh_op_top_4')
// (13, 7, 'local_g3_4')
// (13, 7, 'lutff_4/out')
// (13, 7, 'lutff_6/in_1')
// (13, 8, 'neigh_op_bot_4')
// (14, 6, 'neigh_op_tnl_4')
// (14, 7, 'neigh_op_lft_4')
// (14, 8, 'neigh_op_bnl_4')

wire n1723;
// (12, 6, 'neigh_op_tnr_5')
// (12, 7, 'neigh_op_rgt_5')
// (12, 8, 'neigh_op_bnr_5')
// (13, 6, 'neigh_op_top_5')
// (13, 7, 'lutff_5/out')
// (13, 8, 'neigh_op_bot_5')
// (14, 6, 'neigh_op_tnl_5')
// (14, 7, 'neigh_op_lft_5')
// (14, 8, 'local_g3_5')
// (14, 8, 'lutff_0/in_2')
// (14, 8, 'neigh_op_bnl_5')

wire n1724;
// (12, 6, 'neigh_op_tnr_6')
// (12, 7, 'neigh_op_rgt_6')
// (12, 8, 'neigh_op_bnr_6')
// (13, 6, 'neigh_op_top_6')
// (13, 7, 'lutff_6/out')
// (13, 8, 'local_g1_6')
// (13, 8, 'lutff_1/in_0')
// (13, 8, 'neigh_op_bot_6')
// (14, 6, 'neigh_op_tnl_6')
// (14, 7, 'neigh_op_lft_6')
// (14, 8, 'neigh_op_bnl_6')

wire n1725;
// (12, 6, 'neigh_op_tnr_7')
// (12, 7, 'neigh_op_rgt_7')
// (12, 8, 'neigh_op_bnr_7')
// (13, 6, 'neigh_op_top_7')
// (13, 7, 'lutff_7/out')
// (13, 8, 'neigh_op_bot_7')
// (14, 6, 'neigh_op_tnl_7')
// (14, 7, 'local_g0_7')
// (14, 7, 'lutff_7/in_0')
// (14, 7, 'neigh_op_lft_7')
// (14, 8, 'neigh_op_bnl_7')

wire n1726;
// (12, 6, 'sp12_h_r_1')
// (13, 6, 'sp12_h_r_2')
// (14, 6, 'sp12_h_r_5')
// (15, 6, 'local_g0_6')
// (15, 6, 'lutff_0/in_2')
// (15, 6, 'sp12_h_r_6')
// (16, 5, 'neigh_op_tnr_1')
// (16, 6, 'neigh_op_rgt_1')
// (16, 6, 'sp12_h_r_9')
// (16, 7, 'neigh_op_bnr_1')
// (17, 5, 'neigh_op_top_1')
// (17, 6, 'lutff_1/out')
// (17, 6, 'sp12_h_r_10')
// (17, 7, 'neigh_op_bot_1')
// (18, 5, 'neigh_op_tnl_1')
// (18, 6, 'neigh_op_lft_1')
// (18, 6, 'sp12_h_r_13')
// (18, 7, 'neigh_op_bnl_1')
// (19, 6, 'sp12_h_r_14')
// (20, 6, 'sp12_h_r_17')
// (21, 6, 'sp12_h_r_18')
// (22, 6, 'sp12_h_r_21')
// (23, 6, 'sp12_h_r_22')
// (24, 6, 'sp12_h_l_22')

reg n1727 = 0;
// (12, 6, 'sp4_h_r_11')
// (13, 6, 'sp4_h_r_22')
// (14, 3, 'local_g0_6')
// (14, 3, 'lutff_4/in_2')
// (14, 3, 'sp4_h_r_6')
// (14, 6, 'local_g2_3')
// (14, 6, 'lutff_2/in_3')
// (14, 6, 'sp4_h_r_35')
// (15, 2, 'neigh_op_tnr_7')
// (15, 3, 'neigh_op_rgt_7')
// (15, 3, 'sp4_h_r_19')
// (15, 3, 'sp4_r_v_b_46')
// (15, 4, 'neigh_op_bnr_7')
// (15, 4, 'sp4_r_v_b_35')
// (15, 5, 'sp4_r_v_b_22')
// (15, 6, 'local_g2_3')
// (15, 6, 'lutff_7/in_0')
// (15, 6, 'sp4_h_r_46')
// (15, 6, 'sp4_r_v_b_11')
// (16, 2, 'neigh_op_top_7')
// (16, 2, 'sp4_v_t_46')
// (16, 3, 'lutff_7/out')
// (16, 3, 'sp4_h_r_30')
// (16, 3, 'sp4_v_b_46')
// (16, 4, 'neigh_op_bot_7')
// (16, 4, 'sp4_v_b_35')
// (16, 5, 'sp4_v_b_22')
// (16, 6, 'sp4_h_l_46')
// (16, 6, 'sp4_v_b_11')
// (17, 2, 'neigh_op_tnl_7')
// (17, 3, 'neigh_op_lft_7')
// (17, 3, 'sp4_h_r_43')
// (17, 4, 'neigh_op_bnl_7')
// (18, 3, 'sp4_h_l_43')

reg n1728 = 0;
// (12, 6, 'sp4_h_r_9')
// (12, 9, 'local_g3_7')
// (12, 9, 'lutff_5/in_3')
// (12, 9, 'neigh_op_tnr_7')
// (12, 10, 'neigh_op_rgt_7')
// (12, 10, 'sp4_h_r_3')
// (12, 11, 'neigh_op_bnr_7')
// (13, 6, 'sp4_h_r_20')
// (13, 8, 'sp4_r_v_b_39')
// (13, 9, 'neigh_op_top_7')
// (13, 9, 'sp4_r_v_b_26')
// (13, 10, 'lutff_7/out')
// (13, 10, 'sp4_h_r_14')
// (13, 10, 'sp4_r_v_b_15')
// (13, 11, 'local_g0_7')
// (13, 11, 'lutff_7/in_0')
// (13, 11, 'neigh_op_bot_7')
// (13, 11, 'sp4_r_v_b_2')
// (14, 6, 'sp4_h_r_33')
// (14, 7, 'sp4_v_t_39')
// (14, 8, 'sp4_v_b_39')
// (14, 9, 'neigh_op_tnl_7')
// (14, 9, 'sp4_v_b_26')
// (14, 10, 'neigh_op_lft_7')
// (14, 10, 'sp4_h_r_27')
// (14, 10, 'sp4_v_b_15')
// (14, 11, 'neigh_op_bnl_7')
// (14, 11, 'sp4_h_r_2')
// (14, 11, 'sp4_v_b_2')
// (15, 3, 'sp4_r_v_b_38')
// (15, 4, 'sp4_r_v_b_27')
// (15, 5, 'local_g2_6')
// (15, 5, 'lutff_1/in_1')
// (15, 5, 'sp4_r_v_b_14')
// (15, 6, 'local_g2_4')
// (15, 6, 'lutff_6/in_2')
// (15, 6, 'sp4_h_r_44')
// (15, 6, 'sp4_r_v_b_3')
// (15, 7, 'sp4_r_v_b_38')
// (15, 8, 'sp4_r_v_b_27')
// (15, 9, 'sp4_r_v_b_14')
// (15, 10, 'sp4_h_r_38')
// (15, 10, 'sp4_r_v_b_3')
// (15, 11, 'local_g1_7')
// (15, 11, 'lutff_3/in_3')
// (15, 11, 'sp4_h_r_15')
// (15, 11, 'sp4_r_v_b_38')
// (15, 12, 'sp4_r_v_b_27')
// (15, 13, 'local_g2_6')
// (15, 13, 'lutff_0/in_2')
// (15, 13, 'sp4_r_v_b_14')
// (15, 14, 'sp4_r_v_b_3')
// (16, 2, 'sp4_v_t_38')
// (16, 3, 'sp4_v_b_38')
// (16, 4, 'sp4_v_b_27')
// (16, 5, 'sp4_v_b_14')
// (16, 6, 'sp4_h_l_44')
// (16, 6, 'sp4_v_b_3')
// (16, 6, 'sp4_v_t_38')
// (16, 7, 'sp4_v_b_38')
// (16, 8, 'sp4_v_b_27')
// (16, 9, 'sp4_v_b_14')
// (16, 10, 'sp4_h_l_38')
// (16, 10, 'sp4_v_b_3')
// (16, 10, 'sp4_v_t_38')
// (16, 11, 'sp4_h_r_26')
// (16, 11, 'sp4_v_b_38')
// (16, 12, 'sp4_v_b_27')
// (16, 13, 'sp4_v_b_14')
// (16, 14, 'sp4_v_b_3')
// (17, 11, 'sp4_h_r_39')
// (18, 11, 'sp4_h_l_39')

wire n1729;
// (12, 6, 'sp4_r_v_b_44')
// (12, 7, 'neigh_op_tnr_2')
// (12, 7, 'sp4_r_v_b_33')
// (12, 8, 'neigh_op_rgt_2')
// (12, 8, 'sp4_r_v_b_20')
// (12, 9, 'neigh_op_bnr_2')
// (12, 9, 'sp4_r_v_b_9')
// (13, 5, 'sp4_v_t_44')
// (13, 6, 'sp4_v_b_44')
// (13, 7, 'neigh_op_top_2')
// (13, 7, 'sp4_v_b_33')
// (13, 8, 'lutff_2/out')
// (13, 8, 'sp4_v_b_20')
// (13, 9, 'local_g0_1')
// (13, 9, 'lutff_5/in_2')
// (13, 9, 'neigh_op_bot_2')
// (13, 9, 'sp4_v_b_9')
// (14, 7, 'neigh_op_tnl_2')
// (14, 8, 'neigh_op_lft_2')
// (14, 9, 'neigh_op_bnl_2')

reg n1730 = 0;
// (12, 7, 'local_g2_7')
// (12, 7, 'lutff_4/in_3')
// (12, 7, 'sp4_r_v_b_39')
// (12, 8, 'sp4_r_v_b_26')
// (12, 9, 'neigh_op_tnr_1')
// (12, 9, 'sp4_r_v_b_15')
// (12, 10, 'neigh_op_rgt_1')
// (12, 10, 'sp4_r_v_b_2')
// (12, 11, 'neigh_op_bnr_1')
// (13, 5, 'sp4_r_v_b_39')
// (13, 6, 'sp4_r_v_b_26')
// (13, 6, 'sp4_v_t_39')
// (13, 7, 'sp4_r_v_b_15')
// (13, 7, 'sp4_v_b_39')
// (13, 8, 'sp4_r_v_b_2')
// (13, 8, 'sp4_v_b_26')
// (13, 9, 'neigh_op_top_1')
// (13, 9, 'sp4_r_v_b_46')
// (13, 9, 'sp4_v_b_15')
// (13, 10, 'local_g1_1')
// (13, 10, 'lutff_1/out')
// (13, 10, 'lutff_3/in_1')
// (13, 10, 'sp4_r_v_b_35')
// (13, 10, 'sp4_v_b_2')
// (13, 11, 'neigh_op_bot_1')
// (13, 11, 'sp4_r_v_b_22')
// (13, 12, 'sp4_r_v_b_11')
// (14, 4, 'sp4_v_t_39')
// (14, 5, 'sp4_v_b_39')
// (14, 6, 'local_g3_2')
// (14, 6, 'lutff_1/in_2')
// (14, 6, 'sp4_v_b_26')
// (14, 7, 'sp4_v_b_15')
// (14, 8, 'sp4_v_b_2')
// (14, 8, 'sp4_v_t_46')
// (14, 9, 'neigh_op_tnl_1')
// (14, 9, 'sp4_v_b_46')
// (14, 10, 'neigh_op_lft_1')
// (14, 10, 'sp4_v_b_35')
// (14, 11, 'neigh_op_bnl_1')
// (14, 11, 'sp4_v_b_22')
// (14, 12, 'local_g1_3')
// (14, 12, 'lutff_4/in_2')
// (14, 12, 'sp4_v_b_11')

reg n1731 = 0;
// (12, 7, 'local_g3_4')
// (12, 7, 'lutff_7/in_2')
// (12, 7, 'sp4_r_v_b_44')
// (12, 8, 'sp4_r_v_b_33')
// (12, 9, 'sp4_h_r_8')
// (12, 9, 'sp4_r_v_b_20')
// (12, 10, 'sp4_r_v_b_9')
// (13, 6, 'sp4_h_r_3')
// (13, 6, 'sp4_v_t_44')
// (13, 7, 'sp4_v_b_44')
// (13, 8, 'sp4_v_b_33')
// (13, 9, 'local_g1_5')
// (13, 9, 'lutff_1/in_3')
// (13, 9, 'sp4_h_r_21')
// (13, 9, 'sp4_v_b_20')
// (13, 10, 'sp4_v_b_9')
// (14, 6, 'sp4_h_r_14')
// (14, 9, 'sp4_h_r_32')
// (15, 5, 'neigh_op_tnr_3')
// (15, 6, 'neigh_op_rgt_3')
// (15, 6, 'sp4_h_r_27')
// (15, 6, 'sp4_r_v_b_38')
// (15, 7, 'neigh_op_bnr_3')
// (15, 7, 'sp4_r_v_b_27')
// (15, 8, 'sp4_r_v_b_14')
// (15, 9, 'local_g1_3')
// (15, 9, 'lutff_5/in_1')
// (15, 9, 'sp4_h_r_45')
// (15, 9, 'sp4_r_v_b_3')
// (16, 5, 'neigh_op_top_3')
// (16, 5, 'sp4_v_t_38')
// (16, 6, 'local_g1_3')
// (16, 6, 'lutff_2/in_2')
// (16, 6, 'lutff_3/out')
// (16, 6, 'lutff_6/in_0')
// (16, 6, 'sp4_h_r_38')
// (16, 6, 'sp4_v_b_38')
// (16, 7, 'neigh_op_bot_3')
// (16, 7, 'sp4_v_b_27')
// (16, 8, 'sp4_v_b_14')
// (16, 9, 'sp4_h_l_45')
// (16, 9, 'sp4_v_b_3')
// (17, 5, 'neigh_op_tnl_3')
// (17, 6, 'neigh_op_lft_3')
// (17, 6, 'sp4_h_l_38')
// (17, 7, 'neigh_op_bnl_3')

reg n1732 = 0;
// (12, 7, 'local_g3_7')
// (12, 7, 'lutff_5/in_1')
// (12, 7, 'sp4_r_v_b_47')
// (12, 8, 'sp4_r_v_b_34')
// (12, 9, 'neigh_op_tnr_5')
// (12, 9, 'sp4_r_v_b_23')
// (12, 10, 'neigh_op_rgt_5')
// (12, 10, 'sp4_r_v_b_10')
// (12, 11, 'local_g1_5')
// (12, 11, 'lutff_1/in_1')
// (12, 11, 'neigh_op_bnr_5')
// (13, 6, 'sp4_v_t_47')
// (13, 7, 'sp4_v_b_47')
// (13, 8, 'sp4_v_b_34')
// (13, 9, 'local_g0_5')
// (13, 9, 'lutff_6/in_1')
// (13, 9, 'neigh_op_top_5')
// (13, 9, 'sp4_v_b_23')
// (13, 10, 'lutff_5/out')
// (13, 10, 'sp4_r_v_b_43')
// (13, 10, 'sp4_v_b_10')
// (13, 11, 'neigh_op_bot_5')
// (13, 11, 'sp4_r_v_b_30')
// (13, 12, 'sp4_r_v_b_19')
// (13, 13, 'sp4_r_v_b_6')
// (14, 9, 'neigh_op_tnl_5')
// (14, 9, 'sp4_v_t_43')
// (14, 10, 'neigh_op_lft_5')
// (14, 10, 'sp4_v_b_43')
// (14, 11, 'neigh_op_bnl_5')
// (14, 11, 'sp4_v_b_30')
// (14, 12, 'sp4_v_b_19')
// (14, 13, 'local_g0_6')
// (14, 13, 'lutff_1/in_1')
// (14, 13, 'sp4_v_b_6')

wire n1733;
// (12, 7, 'neigh_op_tnr_1')
// (12, 8, 'neigh_op_rgt_1')
// (12, 9, 'local_g1_1')
// (12, 9, 'lutff_6/in_0')
// (12, 9, 'neigh_op_bnr_1')
// (13, 7, 'neigh_op_top_1')
// (13, 8, 'lutff_1/out')
// (13, 9, 'neigh_op_bot_1')
// (14, 7, 'neigh_op_tnl_1')
// (14, 8, 'neigh_op_lft_1')
// (14, 9, 'neigh_op_bnl_1')

wire n1734;
// (12, 7, 'neigh_op_tnr_3')
// (12, 8, 'neigh_op_rgt_3')
// (12, 9, 'neigh_op_bnr_3')
// (13, 7, 'neigh_op_top_3')
// (13, 8, 'lutff_3/out')
// (13, 9, 'local_g0_3')
// (13, 9, 'lutff_4/in_1')
// (13, 9, 'neigh_op_bot_3')
// (14, 7, 'neigh_op_tnl_3')
// (14, 8, 'neigh_op_lft_3')
// (14, 9, 'neigh_op_bnl_3')

wire n1735;
// (12, 7, 'neigh_op_tnr_4')
// (12, 8, 'neigh_op_rgt_4')
// (12, 9, 'local_g1_4')
// (12, 9, 'lutff_2/in_1')
// (12, 9, 'neigh_op_bnr_4')
// (13, 7, 'neigh_op_top_4')
// (13, 8, 'lutff_4/out')
// (13, 9, 'neigh_op_bot_4')
// (14, 7, 'neigh_op_tnl_4')
// (14, 8, 'neigh_op_lft_4')
// (14, 9, 'neigh_op_bnl_4')

wire n1736;
// (12, 7, 'neigh_op_tnr_5')
// (12, 8, 'neigh_op_rgt_5')
// (12, 9, 'neigh_op_bnr_5')
// (13, 7, 'neigh_op_top_5')
// (13, 8, 'local_g1_5')
// (13, 8, 'lutff_1/in_1')
// (13, 8, 'lutff_5/out')
// (13, 9, 'neigh_op_bot_5')
// (14, 7, 'neigh_op_tnl_5')
// (14, 8, 'neigh_op_lft_5')
// (14, 9, 'neigh_op_bnl_5')

wire n1737;
// (12, 7, 'neigh_op_tnr_6')
// (12, 8, 'neigh_op_rgt_6')
// (12, 9, 'neigh_op_bnr_6')
// (13, 7, 'neigh_op_top_6')
// (13, 8, 'local_g3_6')
// (13, 8, 'lutff_5/in_0')
// (13, 8, 'lutff_6/out')
// (13, 9, 'neigh_op_bot_6')
// (14, 7, 'neigh_op_tnl_6')
// (14, 8, 'neigh_op_lft_6')
// (14, 9, 'neigh_op_bnl_6')

wire n1738;
// (12, 7, 'sp4_h_r_1')
// (13, 7, 'local_g1_4')
// (13, 7, 'lutff_1/in_2')
// (13, 7, 'sp4_h_r_12')
// (14, 3, 'neigh_op_tnr_6')
// (14, 4, 'neigh_op_rgt_6')
// (14, 5, 'neigh_op_bnr_6')
// (14, 7, 'sp4_h_r_25')
// (15, 3, 'neigh_op_top_6')
// (15, 4, 'lutff_6/out')
// (15, 4, 'sp4_r_v_b_45')
// (15, 5, 'neigh_op_bot_6')
// (15, 5, 'sp4_r_v_b_32')
// (15, 6, 'sp4_r_v_b_21')
// (15, 7, 'sp4_h_r_36')
// (15, 7, 'sp4_r_v_b_8')
// (16, 3, 'neigh_op_tnl_6')
// (16, 3, 'sp4_v_t_45')
// (16, 4, 'neigh_op_lft_6')
// (16, 4, 'sp4_v_b_45')
// (16, 5, 'neigh_op_bnl_6')
// (16, 5, 'sp4_v_b_32')
// (16, 6, 'sp4_v_b_21')
// (16, 7, 'sp4_h_l_36')
// (16, 7, 'sp4_v_b_8')

wire n1739;
// (12, 7, 'sp4_h_r_9')
// (13, 7, 'sp4_h_r_20')
// (14, 7, 'sp4_h_r_33')
// (14, 9, 'local_g0_2')
// (14, 9, 'lutff_global/cen')
// (14, 9, 'sp4_h_r_10')
// (15, 4, 'sp4_r_v_b_38')
// (15, 5, 'sp4_r_v_b_27')
// (15, 6, 'sp4_r_v_b_14')
// (15, 7, 'local_g1_3')
// (15, 7, 'lutff_global/cen')
// (15, 7, 'sp4_h_r_44')
// (15, 7, 'sp4_r_v_b_3')
// (15, 9, 'sp4_h_r_23')
// (16, 3, 'sp4_v_t_38')
// (16, 4, 'sp4_v_b_38')
// (16, 5, 'sp4_v_b_27')
// (16, 6, 'neigh_op_tnr_6')
// (16, 6, 'sp4_v_b_14')
// (16, 7, 'neigh_op_rgt_6')
// (16, 7, 'sp4_h_l_44')
// (16, 7, 'sp4_h_r_1')
// (16, 7, 'sp4_v_b_3')
// (16, 8, 'neigh_op_bnr_6')
// (16, 9, 'sp4_h_r_34')
// (17, 6, 'neigh_op_top_6')
// (17, 6, 'sp4_r_v_b_40')
// (17, 7, 'lutff_6/out')
// (17, 7, 'sp4_h_r_12')
// (17, 7, 'sp4_r_v_b_29')
// (17, 8, 'neigh_op_bot_6')
// (17, 8, 'sp4_r_v_b_16')
// (17, 9, 'sp4_h_r_47')
// (17, 9, 'sp4_r_v_b_5')
// (18, 5, 'sp4_v_t_40')
// (18, 6, 'neigh_op_tnl_6')
// (18, 6, 'sp4_v_b_40')
// (18, 7, 'neigh_op_lft_6')
// (18, 7, 'sp4_h_r_25')
// (18, 7, 'sp4_v_b_29')
// (18, 8, 'neigh_op_bnl_6')
// (18, 8, 'sp4_v_b_16')
// (18, 9, 'sp4_h_l_47')
// (18, 9, 'sp4_v_b_5')
// (19, 7, 'sp4_h_r_36')
// (20, 7, 'sp4_h_l_36')

reg n1740 = 0;
// (12, 7, 'sp4_r_v_b_36')
// (12, 8, 'sp4_r_v_b_25')
// (12, 8, 'sp4_r_v_b_41')
// (12, 9, 'sp4_r_v_b_12')
// (12, 9, 'sp4_r_v_b_28')
// (12, 9, 'sp4_r_v_b_44')
// (12, 10, 'neigh_op_tnr_2')
// (12, 10, 'sp4_r_v_b_1')
// (12, 10, 'sp4_r_v_b_17')
// (12, 10, 'sp4_r_v_b_33')
// (12, 11, 'neigh_op_rgt_2')
// (12, 11, 'sp4_r_v_b_20')
// (12, 11, 'sp4_r_v_b_36')
// (12, 11, 'sp4_r_v_b_4')
// (12, 12, 'neigh_op_bnr_2')
// (12, 12, 'sp4_r_v_b_25')
// (12, 12, 'sp4_r_v_b_9')
// (12, 13, 'sp4_r_v_b_12')
// (12, 14, 'sp4_r_v_b_1')
// (13, 4, 'sp4_r_v_b_36')
// (13, 5, 'sp4_r_v_b_25')
// (13, 6, 'sp4_h_r_1')
// (13, 6, 'sp4_r_v_b_12')
// (13, 6, 'sp4_v_t_36')
// (13, 7, 'sp4_r_v_b_1')
// (13, 7, 'sp4_v_b_36')
// (13, 7, 'sp4_v_t_41')
// (13, 8, 'local_g3_1')
// (13, 8, 'lutff_4/in_0')
// (13, 8, 'sp4_r_v_b_40')
// (13, 8, 'sp4_v_b_25')
// (13, 8, 'sp4_v_b_41')
// (13, 8, 'sp4_v_t_44')
// (13, 9, 'sp4_r_v_b_29')
// (13, 9, 'sp4_v_b_12')
// (13, 9, 'sp4_v_b_28')
// (13, 9, 'sp4_v_b_44')
// (13, 10, 'neigh_op_top_2')
// (13, 10, 'sp4_r_v_b_16')
// (13, 10, 'sp4_v_b_1')
// (13, 10, 'sp4_v_b_17')
// (13, 10, 'sp4_v_b_33')
// (13, 10, 'sp4_v_t_36')
// (13, 11, 'lutff_2/out')
// (13, 11, 'sp4_r_v_b_5')
// (13, 11, 'sp4_v_b_20')
// (13, 11, 'sp4_v_b_36')
// (13, 11, 'sp4_v_b_4')
// (13, 12, 'neigh_op_bot_2')
// (13, 12, 'sp4_h_r_9')
// (13, 12, 'sp4_v_b_25')
// (13, 12, 'sp4_v_b_9')
// (13, 13, 'sp4_v_b_12')
// (13, 14, 'sp4_v_b_1')
// (14, 3, 'sp4_v_t_36')
// (14, 4, 'sp4_v_b_36')
// (14, 5, 'sp4_v_b_25')
// (14, 6, 'local_g0_4')
// (14, 6, 'lutff_6/in_0')
// (14, 6, 'sp4_h_r_12')
// (14, 6, 'sp4_v_b_12')
// (14, 7, 'sp4_v_b_1')
// (14, 7, 'sp4_v_t_40')
// (14, 8, 'sp4_v_b_40')
// (14, 9, 'sp4_v_b_29')
// (14, 10, 'local_g3_2')
// (14, 10, 'lutff_3/in_2')
// (14, 10, 'neigh_op_tnl_2')
// (14, 10, 'sp4_v_b_16')
// (14, 11, 'neigh_op_lft_2')
// (14, 11, 'sp4_v_b_5')
// (14, 12, 'local_g2_2')
// (14, 12, 'lutff_5/in_3')
// (14, 12, 'neigh_op_bnl_2')
// (14, 12, 'sp4_h_r_20')
// (15, 6, 'local_g3_1')
// (15, 6, 'lutff_1/in_3')
// (15, 6, 'sp4_h_r_25')
// (15, 12, 'local_g3_1')
// (15, 12, 'lutff_7/in_1')
// (15, 12, 'sp4_h_r_33')
// (16, 6, 'sp4_h_r_36')
// (16, 12, 'sp4_h_r_44')
// (17, 6, 'sp4_h_l_36')
// (17, 12, 'sp4_h_l_44')

reg n1741 = 0;
// (12, 8, 'local_g3_7')
// (12, 8, 'lutff_5/in_3')
// (12, 8, 'neigh_op_tnr_7')
// (12, 9, 'neigh_op_rgt_7')
// (12, 10, 'neigh_op_bnr_7')
// (13, 4, 'sp12_v_t_22')
// (13, 5, 'sp12_v_b_22')
// (13, 6, 'sp12_v_b_21')
// (13, 7, 'sp12_v_b_18')
// (13, 8, 'local_g0_7')
// (13, 8, 'lutff_3/in_2')
// (13, 8, 'neigh_op_top_7')
// (13, 8, 'sp12_v_b_17')
// (13, 9, 'lutff_7/out')
// (13, 9, 'sp12_v_b_14')
// (13, 10, 'local_g0_7')
// (13, 10, 'lutff_5/in_0')
// (13, 10, 'neigh_op_bot_7')
// (13, 10, 'sp12_v_b_13')
// (13, 11, 'sp12_v_b_10')
// (13, 12, 'sp12_v_b_9')
// (13, 13, 'sp12_v_b_6')
// (13, 14, 'local_g3_5')
// (13, 14, 'lutff_0/in_0')
// (13, 14, 'sp12_v_b_5')
// (13, 15, 'sp12_v_b_2')
// (13, 16, 'sp12_v_b_1')
// (14, 8, 'neigh_op_tnl_7')
// (14, 9, 'neigh_op_lft_7')
// (14, 10, 'neigh_op_bnl_7')

wire n1742;
// (12, 8, 'neigh_op_tnr_0')
// (12, 9, 'local_g3_0')
// (12, 9, 'lutff_6/in_1')
// (12, 9, 'neigh_op_rgt_0')
// (12, 10, 'neigh_op_bnr_0')
// (13, 8, 'neigh_op_top_0')
// (13, 9, 'lutff_0/out')
// (13, 10, 'neigh_op_bot_0')
// (14, 8, 'neigh_op_tnl_0')
// (14, 9, 'neigh_op_lft_0')
// (14, 10, 'neigh_op_bnl_0')

wire n1743;
// (12, 8, 'neigh_op_tnr_1')
// (12, 9, 'neigh_op_rgt_1')
// (12, 10, 'neigh_op_bnr_1')
// (13, 8, 'neigh_op_top_1')
// (13, 9, 'local_g2_1')
// (13, 9, 'lutff_1/out')
// (13, 9, 'lutff_4/in_3')
// (13, 10, 'neigh_op_bot_1')
// (14, 8, 'neigh_op_tnl_1')
// (14, 9, 'neigh_op_lft_1')
// (14, 10, 'neigh_op_bnl_1')

wire n1744;
// (12, 8, 'neigh_op_tnr_3')
// (12, 9, 'neigh_op_rgt_3')
// (12, 10, 'neigh_op_bnr_3')
// (13, 8, 'neigh_op_top_3')
// (13, 9, 'local_g1_3')
// (13, 9, 'lutff_3/out')
// (13, 9, 'lutff_4/in_0')
// (13, 10, 'neigh_op_bot_3')
// (14, 8, 'neigh_op_tnl_3')
// (14, 9, 'neigh_op_lft_3')
// (14, 10, 'neigh_op_bnl_3')

wire n1745;
// (12, 8, 'neigh_op_tnr_4')
// (12, 9, 'neigh_op_rgt_4')
// (12, 10, 'neigh_op_bnr_4')
// (13, 8, 'local_g0_4')
// (13, 8, 'lutff_5/in_3')
// (13, 8, 'neigh_op_top_4')
// (13, 9, 'lutff_4/out')
// (13, 10, 'neigh_op_bot_4')
// (14, 8, 'neigh_op_tnl_4')
// (14, 9, 'neigh_op_lft_4')
// (14, 10, 'neigh_op_bnl_4')

wire n1746;
// (12, 8, 'neigh_op_tnr_5')
// (12, 9, 'neigh_op_rgt_5')
// (12, 10, 'neigh_op_bnr_5')
// (13, 8, 'local_g0_5')
// (13, 8, 'lutff_5/in_2')
// (13, 8, 'neigh_op_top_5')
// (13, 9, 'lutff_5/out')
// (13, 10, 'neigh_op_bot_5')
// (14, 8, 'neigh_op_tnl_5')
// (14, 9, 'neigh_op_lft_5')
// (14, 10, 'neigh_op_bnl_5')

wire n1747;
// (12, 8, 'neigh_op_tnr_6')
// (12, 9, 'neigh_op_rgt_6')
// (12, 10, 'neigh_op_bnr_6')
// (13, 8, 'neigh_op_top_6')
// (13, 9, 'local_g0_6')
// (13, 9, 'lutff_4/in_2')
// (13, 9, 'lutff_6/out')
// (13, 10, 'neigh_op_bot_6')
// (14, 8, 'neigh_op_tnl_6')
// (14, 9, 'neigh_op_lft_6')
// (14, 10, 'neigh_op_bnl_6')

reg n1748 = 0;
// (12, 8, 'sp4_h_r_2')
// (13, 7, 'neigh_op_tnr_5')
// (13, 8, 'neigh_op_rgt_5')
// (13, 8, 'sp4_h_r_15')
// (13, 9, 'neigh_op_bnr_5')
// (14, 7, 'neigh_op_top_5')
// (14, 8, 'lutff_5/out')
// (14, 8, 'sp4_h_r_26')
// (14, 9, 'neigh_op_bot_5')
// (15, 7, 'neigh_op_tnl_5')
// (15, 8, 'neigh_op_lft_5')
// (15, 8, 'sp4_h_r_39')
// (15, 9, 'neigh_op_bnl_5')
// (15, 9, 'sp4_r_v_b_39')
// (15, 10, 'sp4_r_v_b_26')
// (15, 11, 'sp4_r_v_b_15')
// (15, 12, 'sp4_r_v_b_2')
// (16, 8, 'sp4_h_l_39')
// (16, 8, 'sp4_v_t_39')
// (16, 9, 'local_g3_7')
// (16, 9, 'lutff_6/in_0')
// (16, 9, 'sp4_v_b_39')
// (16, 10, 'sp4_v_b_26')
// (16, 11, 'sp4_v_b_15')
// (16, 12, 'sp4_v_b_2')

reg n1749 = 0;
// (12, 8, 'sp4_r_v_b_36')
// (12, 9, 'local_g3_6')
// (12, 9, 'lutff_4/in_1')
// (12, 9, 'neigh_op_tnr_6')
// (12, 9, 'sp4_r_v_b_25')
// (12, 10, 'neigh_op_rgt_6')
// (12, 10, 'sp4_r_v_b_12')
// (12, 11, 'neigh_op_bnr_6')
// (12, 11, 'sp4_r_v_b_1')
// (13, 7, 'local_g1_6')
// (13, 7, 'lutff_0/in_3')
// (13, 7, 'sp4_h_r_1')
// (13, 7, 'sp4_h_r_6')
// (13, 7, 'sp4_v_t_36')
// (13, 8, 'sp4_v_b_36')
// (13, 9, 'neigh_op_top_6')
// (13, 9, 'sp4_v_b_25')
// (13, 10, 'lutff_6/out')
// (13, 10, 'sp4_v_b_12')
// (13, 11, 'neigh_op_bot_6')
// (13, 11, 'sp4_h_r_7')
// (13, 11, 'sp4_v_b_1')
// (14, 7, 'sp4_h_r_12')
// (14, 7, 'sp4_h_r_19')
// (14, 9, 'neigh_op_tnl_6')
// (14, 10, 'neigh_op_lft_6')
// (14, 11, 'local_g2_6')
// (14, 11, 'lutff_2/in_0')
// (14, 11, 'lutff_4/in_0')
// (14, 11, 'neigh_op_bnl_6')
// (14, 11, 'sp4_h_r_18')
// (15, 7, 'local_g3_1')
// (15, 7, 'lutff_1/in_3')
// (15, 7, 'sp4_h_r_25')
// (15, 7, 'sp4_h_r_30')
// (15, 11, 'local_g3_7')
// (15, 11, 'lutff_6/in_0')
// (15, 11, 'sp4_h_r_31')
// (16, 7, 'sp4_h_r_36')
// (16, 7, 'sp4_h_r_43')
// (16, 11, 'sp4_h_r_42')
// (17, 7, 'sp4_h_l_36')
// (17, 7, 'sp4_h_l_43')
// (17, 11, 'sp4_h_l_42')

reg n1750 = 0;
// (12, 8, 'sp4_r_v_b_39')
// (12, 9, 'sp4_r_v_b_26')
// (12, 10, 'neigh_op_tnr_1')
// (12, 10, 'sp4_r_v_b_15')
// (12, 11, 'neigh_op_rgt_1')
// (12, 11, 'sp4_r_v_b_2')
// (12, 12, 'neigh_op_bnr_1')
// (13, 7, 'sp4_v_t_39')
// (13, 8, 'local_g3_7')
// (13, 8, 'lutff_7/in_1')
// (13, 8, 'sp4_v_b_39')
// (13, 9, 'sp4_r_v_b_43')
// (13, 9, 'sp4_v_b_26')
// (13, 10, 'local_g0_1')
// (13, 10, 'lutff_2/in_1')
// (13, 10, 'neigh_op_top_1')
// (13, 10, 'sp4_r_v_b_30')
// (13, 10, 'sp4_v_b_15')
// (13, 11, 'lutff_1/out')
// (13, 11, 'sp4_r_v_b_19')
// (13, 11, 'sp4_v_b_2')
// (13, 12, 'neigh_op_bot_1')
// (13, 12, 'sp4_r_v_b_6')
// (14, 8, 'local_g0_6')
// (14, 8, 'lutff_3/in_1')
// (14, 8, 'sp4_h_r_6')
// (14, 8, 'sp4_v_t_43')
// (14, 9, 'sp4_v_b_43')
// (14, 10, 'neigh_op_tnl_1')
// (14, 10, 'sp4_v_b_30')
// (14, 11, 'neigh_op_lft_1')
// (14, 11, 'sp4_v_b_19')
// (14, 12, 'local_g3_1')
// (14, 12, 'lutff_3/in_3')
// (14, 12, 'neigh_op_bnl_1')
// (14, 12, 'sp4_v_b_6')
// (15, 8, 'sp4_h_r_19')
// (16, 8, 'sp4_h_r_30')
// (17, 8, 'sp4_h_r_43')
// (18, 8, 'sp4_h_l_43')

reg n1751 = 0;
// (12, 8, 'sp4_r_v_b_45')
// (12, 9, 'sp4_r_v_b_32')
// (12, 10, 'neigh_op_tnr_4')
// (12, 10, 'sp4_r_v_b_21')
// (12, 11, 'neigh_op_rgt_4')
// (12, 11, 'sp4_r_v_b_8')
// (12, 12, 'neigh_op_bnr_4')
// (13, 7, 'sp4_v_t_45')
// (13, 8, 'sp4_v_b_45')
// (13, 9, 'local_g2_0')
// (13, 9, 'lutff_3/in_3')
// (13, 9, 'lutff_5/in_3')
// (13, 9, 'sp4_v_b_32')
// (13, 10, 'neigh_op_top_4')
// (13, 10, 'sp4_v_b_21')
// (13, 11, 'lutff_4/out')
// (13, 11, 'sp4_v_b_8')
// (13, 12, 'local_g0_4')
// (13, 12, 'lutff_0/in_0')
// (13, 12, 'neigh_op_bot_4')
// (14, 10, 'neigh_op_tnl_4')
// (14, 11, 'neigh_op_lft_4')
// (14, 12, 'neigh_op_bnl_4')

reg n1752 = 0;
// (12, 9, 'local_g3_2')
// (12, 9, 'lutff_0/in_3')
// (12, 9, 'neigh_op_tnr_2')
// (12, 10, 'neigh_op_rgt_2')
// (12, 11, 'neigh_op_bnr_2')
// (13, 7, 'sp4_r_v_b_40')
// (13, 8, 'sp4_r_v_b_29')
// (13, 9, 'local_g3_0')
// (13, 9, 'lutff_7/in_2')
// (13, 9, 'neigh_op_top_2')
// (13, 9, 'sp4_r_v_b_16')
// (13, 10, 'lutff_2/out')
// (13, 10, 'sp4_r_v_b_37')
// (13, 10, 'sp4_r_v_b_5')
// (13, 11, 'neigh_op_bot_2')
// (13, 11, 'sp4_r_v_b_24')
// (13, 12, 'sp4_r_v_b_13')
// (13, 13, 'sp4_r_v_b_0')
// (14, 6, 'sp4_v_t_40')
// (14, 7, 'sp4_v_b_40')
// (14, 8, 'local_g2_5')
// (14, 8, 'lutff_2/in_3')
// (14, 8, 'sp4_v_b_29')
// (14, 9, 'neigh_op_tnl_2')
// (14, 9, 'sp4_v_b_16')
// (14, 9, 'sp4_v_t_37')
// (14, 10, 'neigh_op_lft_2')
// (14, 10, 'sp4_v_b_37')
// (14, 10, 'sp4_v_b_5')
// (14, 11, 'neigh_op_bnl_2')
// (14, 11, 'sp4_v_b_24')
// (14, 12, 'local_g1_5')
// (14, 12, 'lutff_6/in_0')
// (14, 12, 'sp4_v_b_13')
// (14, 13, 'sp4_v_b_0')

reg n1753 = 0;
// (12, 9, 'neigh_op_tnr_0')
// (12, 10, 'neigh_op_rgt_0')
// (12, 11, 'neigh_op_bnr_0')
// (13, 3, 'sp4_r_v_b_41')
// (13, 4, 'sp4_r_v_b_28')
// (13, 5, 'sp4_r_v_b_17')
// (13, 6, 'local_g1_4')
// (13, 6, 'lutff_3/in_0')
// (13, 6, 'sp4_r_v_b_4')
// (13, 7, 'sp4_r_v_b_36')
// (13, 8, 'sp4_r_v_b_25')
// (13, 9, 'neigh_op_top_0')
// (13, 9, 'sp4_r_v_b_12')
// (13, 9, 'sp4_r_v_b_44')
// (13, 10, 'local_g0_0')
// (13, 10, 'lutff_0/out')
// (13, 10, 'lutff_4/in_2')
// (13, 10, 'sp4_r_v_b_1')
// (13, 10, 'sp4_r_v_b_33')
// (13, 11, 'neigh_op_bot_0')
// (13, 11, 'sp4_r_v_b_20')
// (13, 12, 'sp4_r_v_b_9')
// (14, 2, 'sp4_v_t_41')
// (14, 3, 'sp4_v_b_41')
// (14, 4, 'sp4_v_b_28')
// (14, 5, 'sp4_v_b_17')
// (14, 6, 'local_g1_1')
// (14, 6, 'lutff_3/in_1')
// (14, 6, 'sp4_h_r_1')
// (14, 6, 'sp4_v_b_4')
// (14, 6, 'sp4_v_t_36')
// (14, 7, 'sp4_v_b_36')
// (14, 8, 'sp4_v_b_25')
// (14, 8, 'sp4_v_t_44')
// (14, 9, 'neigh_op_tnl_0')
// (14, 9, 'sp4_v_b_12')
// (14, 9, 'sp4_v_b_44')
// (14, 10, 'neigh_op_lft_0')
// (14, 10, 'sp4_v_b_1')
// (14, 10, 'sp4_v_b_33')
// (14, 11, 'neigh_op_bnl_0')
// (14, 11, 'sp4_v_b_20')
// (14, 12, 'local_g1_1')
// (14, 12, 'lutff_7/in_1')
// (14, 12, 'sp4_v_b_9')
// (15, 6, 'sp4_h_r_12')
// (16, 6, 'sp4_h_r_25')
// (17, 6, 'sp4_h_r_36')
// (18, 6, 'sp4_h_l_36')

reg n1754 = 0;
// (12, 9, 'sp4_h_r_0')
// (13, 9, 'sp4_h_r_13')
// (13, 12, 'sp4_h_r_4')
// (14, 9, 'local_g3_0')
// (14, 9, 'lutff_6/in_1')
// (14, 9, 'sp4_h_r_24')
// (14, 11, 'neigh_op_tnr_6')
// (14, 12, 'neigh_op_rgt_6')
// (14, 12, 'sp4_h_r_17')
// (14, 13, 'neigh_op_bnr_6')
// (15, 9, 'sp4_h_r_37')
// (15, 10, 'sp4_r_v_b_37')
// (15, 11, 'local_g1_6')
// (15, 11, 'lutff_7/in_2')
// (15, 11, 'neigh_op_top_6')
// (15, 11, 'sp4_r_v_b_24')
// (15, 11, 'sp4_r_v_b_40')
// (15, 12, 'lutff_6/out')
// (15, 12, 'sp4_h_r_28')
// (15, 12, 'sp4_r_v_b_13')
// (15, 12, 'sp4_r_v_b_29')
// (15, 13, 'neigh_op_bot_6')
// (15, 13, 'sp4_r_v_b_0')
// (15, 13, 'sp4_r_v_b_16')
// (15, 14, 'sp4_r_v_b_5')
// (16, 9, 'sp4_h_l_37')
// (16, 9, 'sp4_r_v_b_47')
// (16, 9, 'sp4_v_t_37')
// (16, 10, 'sp4_h_r_10')
// (16, 10, 'sp4_h_r_5')
// (16, 10, 'sp4_r_v_b_34')
// (16, 10, 'sp4_v_b_37')
// (16, 10, 'sp4_v_t_40')
// (16, 11, 'local_g2_6')
// (16, 11, 'lutff_2/in_2')
// (16, 11, 'neigh_op_tnl_6')
// (16, 11, 'sp4_r_v_b_23')
// (16, 11, 'sp4_v_b_24')
// (16, 11, 'sp4_v_b_40')
// (16, 12, 'local_g1_6')
// (16, 12, 'lutff_1/in_2')
// (16, 12, 'neigh_op_lft_6')
// (16, 12, 'sp4_h_r_41')
// (16, 12, 'sp4_r_v_b_10')
// (16, 12, 'sp4_v_b_13')
// (16, 12, 'sp4_v_b_29')
// (16, 13, 'neigh_op_bnl_6')
// (16, 13, 'sp4_v_b_0')
// (16, 13, 'sp4_v_b_16')
// (16, 14, 'sp4_v_b_5')
// (17, 8, 'local_g0_2')
// (17, 8, 'lutff_3/in_1')
// (17, 8, 'sp4_h_r_10')
// (17, 8, 'sp4_v_t_47')
// (17, 9, 'local_g3_7')
// (17, 9, 'lutff_6/in_2')
// (17, 9, 'sp4_v_b_47')
// (17, 10, 'local_g1_0')
// (17, 10, 'lutff_3/in_2')
// (17, 10, 'sp4_h_r_16')
// (17, 10, 'sp4_h_r_23')
// (17, 10, 'sp4_v_b_34')
// (17, 11, 'sp4_v_b_23')
// (17, 12, 'sp4_h_l_41')
// (17, 12, 'sp4_v_b_10')
// (18, 8, 'sp4_h_r_23')
// (18, 10, 'sp4_h_r_29')
// (18, 10, 'sp4_h_r_34')
// (19, 7, 'sp4_r_v_b_47')
// (19, 8, 'sp4_h_r_34')
// (19, 8, 'sp4_r_v_b_34')
// (19, 9, 'sp4_r_v_b_23')
// (19, 10, 'sp4_h_r_40')
// (19, 10, 'sp4_h_r_47')
// (19, 10, 'sp4_r_v_b_10')
// (20, 6, 'sp4_v_t_47')
// (20, 7, 'sp4_v_b_47')
// (20, 8, 'sp4_h_r_47')
// (20, 8, 'sp4_v_b_34')
// (20, 9, 'local_g1_7')
// (20, 9, 'lutff_4/in_2')
// (20, 9, 'sp4_v_b_23')
// (20, 10, 'sp4_h_l_40')
// (20, 10, 'sp4_h_l_47')
// (20, 10, 'sp4_v_b_10')
// (21, 8, 'sp4_h_l_47')

reg n1755 = 0;
// (12, 9, 'sp4_h_r_10')
// (13, 9, 'sp4_h_r_23')
// (14, 9, 'local_g3_2')
// (14, 9, 'lutff_5/in_0')
// (14, 9, 'sp4_h_r_34')
// (15, 7, 'sp4_r_v_b_37')
// (15, 8, 'sp4_r_v_b_24')
// (15, 9, 'sp4_h_r_47')
// (15, 9, 'sp4_r_v_b_13')
// (15, 10, 'local_g3_1')
// (15, 10, 'lutff_6/in_0')
// (15, 10, 'sp4_r_v_b_0')
// (15, 10, 'sp4_r_v_b_41')
// (15, 11, 'sp4_r_v_b_28')
// (15, 11, 'sp4_r_v_b_44')
// (15, 12, 'neigh_op_tnr_2')
// (15, 12, 'sp4_r_v_b_17')
// (15, 12, 'sp4_r_v_b_33')
// (15, 13, 'neigh_op_rgt_2')
// (15, 13, 'sp4_r_v_b_20')
// (15, 13, 'sp4_r_v_b_4')
// (15, 14, 'neigh_op_bnr_2')
// (15, 14, 'sp4_r_v_b_9')
// (16, 6, 'sp4_v_t_37')
// (16, 7, 'sp4_r_v_b_41')
// (16, 7, 'sp4_v_b_37')
// (16, 8, 'sp4_r_v_b_28')
// (16, 8, 'sp4_v_b_24')
// (16, 9, 'local_g0_5')
// (16, 9, 'lutff_4/in_3')
// (16, 9, 'sp4_h_l_47')
// (16, 9, 'sp4_r_v_b_17')
// (16, 9, 'sp4_v_b_13')
// (16, 9, 'sp4_v_t_41')
// (16, 10, 'sp4_r_v_b_4')
// (16, 10, 'sp4_v_b_0')
// (16, 10, 'sp4_v_b_41')
// (16, 10, 'sp4_v_t_44')
// (16, 11, 'local_g2_4')
// (16, 11, 'lutff_1/in_3')
// (16, 11, 'sp4_r_v_b_45')
// (16, 11, 'sp4_v_b_28')
// (16, 11, 'sp4_v_b_44')
// (16, 12, 'neigh_op_top_2')
// (16, 12, 'sp4_r_v_b_32')
// (16, 12, 'sp4_v_b_17')
// (16, 12, 'sp4_v_b_33')
// (16, 13, 'local_g0_2')
// (16, 13, 'lutff_2/out')
// (16, 13, 'lutff_3/in_1')
// (16, 13, 'sp4_h_r_4')
// (16, 13, 'sp4_r_v_b_21')
// (16, 13, 'sp4_r_v_b_37')
// (16, 13, 'sp4_v_b_20')
// (16, 13, 'sp4_v_b_4')
// (16, 14, 'neigh_op_bot_2')
// (16, 14, 'sp4_r_v_b_24')
// (16, 14, 'sp4_r_v_b_8')
// (16, 14, 'sp4_v_b_9')
// (16, 15, 'sp4_r_v_b_13')
// (16, 16, 'sp4_r_v_b_0')
// (17, 6, 'sp4_v_t_41')
// (17, 7, 'sp4_v_b_41')
// (17, 8, 'local_g3_4')
// (17, 8, 'lutff_6/in_1')
// (17, 8, 'sp4_v_b_28')
// (17, 9, 'sp4_v_b_17')
// (17, 10, 'sp4_h_r_8')
// (17, 10, 'sp4_v_b_4')
// (17, 10, 'sp4_v_t_45')
// (17, 11, 'sp4_v_b_45')
// (17, 12, 'neigh_op_tnl_2')
// (17, 12, 'sp4_h_r_5')
// (17, 12, 'sp4_v_b_32')
// (17, 12, 'sp4_v_t_37')
// (17, 13, 'neigh_op_lft_2')
// (17, 13, 'sp4_h_r_17')
// (17, 13, 'sp4_v_b_21')
// (17, 13, 'sp4_v_b_37')
// (17, 14, 'neigh_op_bnl_2')
// (17, 14, 'sp4_v_b_24')
// (17, 14, 'sp4_v_b_8')
// (17, 15, 'sp4_v_b_13')
// (17, 16, 'sp4_v_b_0')
// (18, 10, 'local_g0_5')
// (18, 10, 'lutff_7/in_0')
// (18, 10, 'sp4_h_r_21')
// (18, 12, 'sp4_h_r_16')
// (18, 13, 'sp4_h_r_28')
// (19, 10, 'sp4_h_r_32')
// (19, 10, 'sp4_r_v_b_47')
// (19, 11, 'sp4_r_v_b_34')
// (19, 12, 'sp4_h_r_29')
// (19, 12, 'sp4_r_v_b_23')
// (19, 13, 'sp4_h_r_41')
// (19, 13, 'sp4_r_v_b_10')
// (20, 9, 'sp4_r_v_b_40')
// (20, 9, 'sp4_v_t_47')
// (20, 10, 'sp4_h_r_45')
// (20, 10, 'sp4_r_v_b_29')
// (20, 10, 'sp4_v_b_47')
// (20, 11, 'sp4_r_v_b_16')
// (20, 11, 'sp4_v_b_34')
// (20, 12, 'local_g1_7')
// (20, 12, 'lutff_7/in_1')
// (20, 12, 'sp4_h_r_40')
// (20, 12, 'sp4_r_v_b_5')
// (20, 12, 'sp4_v_b_23')
// (20, 13, 'sp4_h_l_41')
// (20, 13, 'sp4_v_b_10')
// (21, 8, 'sp4_v_t_40')
// (21, 9, 'sp4_v_b_40')
// (21, 10, 'sp4_h_l_45')
// (21, 10, 'sp4_v_b_29')
// (21, 11, 'local_g1_0')
// (21, 11, 'lutff_6/in_1')
// (21, 11, 'sp4_v_b_16')
// (21, 12, 'sp4_h_l_40')
// (21, 12, 'sp4_v_b_5')

reg n1756 = 0;
// (12, 9, 'sp4_h_r_2')
// (13, 8, 'neigh_op_tnr_5')
// (13, 9, 'neigh_op_rgt_5')
// (13, 9, 'sp4_h_r_15')
// (13, 10, 'neigh_op_bnr_5')
// (14, 8, 'neigh_op_top_5')
// (14, 9, 'lutff_5/out')
// (14, 9, 'sp4_h_r_26')
// (14, 10, 'neigh_op_bot_5')
// (15, 8, 'neigh_op_tnl_5')
// (15, 9, 'local_g0_5')
// (15, 9, 'lutff_1/in_2')
// (15, 9, 'neigh_op_lft_5')
// (15, 9, 'sp4_h_r_39')
// (15, 10, 'local_g2_5')
// (15, 10, 'lutff_1/in_2')
// (15, 10, 'neigh_op_bnl_5')
// (15, 10, 'sp4_r_v_b_42')
// (15, 11, 'sp4_r_v_b_31')
// (15, 12, 'sp4_r_v_b_18')
// (15, 13, 'sp4_r_v_b_7')
// (16, 9, 'sp4_h_l_39')
// (16, 9, 'sp4_v_t_42')
// (16, 10, 'local_g3_2')
// (16, 10, 'lutff_2/in_3')
// (16, 10, 'sp4_v_b_42')
// (16, 11, 'sp4_v_b_31')
// (16, 12, 'sp4_v_b_18')
// (16, 13, 'sp4_v_b_7')

reg n1757 = 0;
// (12, 9, 'sp4_h_r_6')
// (13, 9, 'sp4_h_r_19')
// (14, 9, 'local_g3_6')
// (14, 9, 'lutff_1/in_2')
// (14, 9, 'sp4_h_r_30')
// (15, 9, 'sp4_h_r_43')
// (15, 10, 'local_g3_3')
// (15, 10, 'lutff_0/in_2')
// (15, 10, 'sp4_r_v_b_43')
// (15, 11, 'sp4_r_v_b_30')
// (15, 12, 'neigh_op_tnr_3')
// (15, 12, 'sp4_r_v_b_19')
// (15, 13, 'local_g2_3')
// (15, 13, 'lutff_7/in_2')
// (15, 13, 'neigh_op_rgt_3')
// (15, 13, 'sp4_h_r_11')
// (15, 13, 'sp4_r_v_b_6')
// (15, 14, 'neigh_op_bnr_3')
// (16, 7, 'sp4_r_v_b_43')
// (16, 8, 'sp4_r_v_b_30')
// (16, 9, 'sp4_h_l_43')
// (16, 9, 'sp4_r_v_b_19')
// (16, 9, 'sp4_r_v_b_39')
// (16, 9, 'sp4_v_t_43')
// (16, 10, 'sp4_r_v_b_26')
// (16, 10, 'sp4_r_v_b_6')
// (16, 10, 'sp4_v_b_43')
// (16, 11, 'sp4_r_v_b_15')
// (16, 11, 'sp4_r_v_b_47')
// (16, 11, 'sp4_v_b_30')
// (16, 12, 'neigh_op_top_3')
// (16, 12, 'sp4_r_v_b_2')
// (16, 12, 'sp4_r_v_b_34')
// (16, 12, 'sp4_v_b_19')
// (16, 13, 'lutff_3/out')
// (16, 13, 'sp4_h_r_22')
// (16, 13, 'sp4_h_r_6')
// (16, 13, 'sp4_r_v_b_23')
// (16, 13, 'sp4_r_v_b_39')
// (16, 13, 'sp4_v_b_6')
// (16, 14, 'neigh_op_bot_3')
// (16, 14, 'sp4_r_v_b_10')
// (16, 14, 'sp4_r_v_b_26')
// (16, 15, 'sp4_r_v_b_15')
// (16, 16, 'sp4_r_v_b_2')
// (17, 6, 'sp4_v_t_43')
// (17, 7, 'sp4_v_b_43')
// (17, 8, 'local_g3_6')
// (17, 8, 'lutff_7/in_2')
// (17, 8, 'sp4_h_r_2')
// (17, 8, 'sp4_v_b_30')
// (17, 8, 'sp4_v_t_39')
// (17, 9, 'sp4_v_b_19')
// (17, 9, 'sp4_v_b_39')
// (17, 10, 'sp4_v_b_26')
// (17, 10, 'sp4_v_b_6')
// (17, 10, 'sp4_v_t_47')
// (17, 11, 'sp4_v_b_15')
// (17, 11, 'sp4_v_b_47')
// (17, 12, 'neigh_op_tnl_3')
// (17, 12, 'sp4_h_r_7')
// (17, 12, 'sp4_v_b_2')
// (17, 12, 'sp4_v_b_34')
// (17, 12, 'sp4_v_t_39')
// (17, 13, 'neigh_op_lft_3')
// (17, 13, 'sp4_h_r_19')
// (17, 13, 'sp4_h_r_35')
// (17, 13, 'sp4_v_b_23')
// (17, 13, 'sp4_v_b_39')
// (17, 14, 'neigh_op_bnl_3')
// (17, 14, 'sp4_v_b_10')
// (17, 14, 'sp4_v_b_26')
// (17, 15, 'sp4_v_b_15')
// (17, 16, 'sp4_v_b_2')
// (18, 6, 'sp4_r_v_b_46')
// (18, 7, 'local_g0_0')
// (18, 7, 'lutff_3/in_1')
// (18, 7, 'sp4_r_v_b_35')
// (18, 8, 'local_g1_7')
// (18, 8, 'lutff_6/in_0')
// (18, 8, 'sp4_h_r_15')
// (18, 8, 'sp4_r_v_b_22')
// (18, 9, 'sp4_r_v_b_11')
// (18, 10, 'sp4_r_v_b_46')
// (18, 11, 'sp4_r_v_b_35')
// (18, 12, 'sp4_h_r_18')
// (18, 12, 'sp4_r_v_b_22')
// (18, 13, 'sp4_h_r_30')
// (18, 13, 'sp4_h_r_46')
// (18, 13, 'sp4_r_v_b_11')
// (19, 5, 'sp4_v_t_46')
// (19, 6, 'sp4_v_b_46')
// (19, 7, 'sp4_v_b_35')
// (19, 8, 'sp4_h_r_26')
// (19, 8, 'sp4_v_b_22')
// (19, 9, 'sp4_v_b_11')
// (19, 9, 'sp4_v_t_46')
// (19, 10, 'sp4_r_v_b_37')
// (19, 10, 'sp4_v_b_46')
// (19, 11, 'sp4_r_v_b_24')
// (19, 11, 'sp4_v_b_35')
// (19, 12, 'sp4_h_r_31')
// (19, 12, 'sp4_r_v_b_13')
// (19, 12, 'sp4_v_b_22')
// (19, 13, 'sp4_h_l_46')
// (19, 13, 'sp4_h_r_43')
// (19, 13, 'sp4_r_v_b_0')
// (19, 13, 'sp4_v_b_11')
// (20, 8, 'sp4_h_r_39')
// (20, 9, 'local_g0_0')
// (20, 9, 'lutff_2/in_2')
// (20, 9, 'sp4_h_r_0')
// (20, 9, 'sp4_r_v_b_42')
// (20, 9, 'sp4_v_t_37')
// (20, 10, 'local_g2_5')
// (20, 10, 'lutff_5/in_0')
// (20, 10, 'sp4_r_v_b_31')
// (20, 10, 'sp4_v_b_37')
// (20, 11, 'sp4_r_v_b_18')
// (20, 11, 'sp4_v_b_24')
// (20, 12, 'sp4_h_r_42')
// (20, 12, 'sp4_r_v_b_7')
// (20, 12, 'sp4_v_b_13')
// (20, 13, 'sp4_h_l_43')
// (20, 13, 'sp4_v_b_0')
// (21, 8, 'sp4_h_l_39')
// (21, 8, 'sp4_v_t_42')
// (21, 9, 'sp4_h_r_13')
// (21, 9, 'sp4_v_b_42')
// (21, 10, 'sp4_v_b_31')
// (21, 11, 'local_g1_2')
// (21, 11, 'lutff_0/in_3')
// (21, 11, 'sp4_v_b_18')
// (21, 12, 'sp4_h_l_42')
// (21, 12, 'sp4_v_b_7')
// (22, 9, 'sp4_h_r_24')
// (23, 9, 'sp4_h_r_37')
// (24, 9, 'sp4_h_l_37')

wire n1758;
// (12, 11, 'neigh_op_tnr_0')
// (12, 12, 'neigh_op_rgt_0')
// (12, 13, 'neigh_op_bnr_0')
// (13, 11, 'neigh_op_top_0')
// (13, 12, 'lutff_0/out')
// (13, 13, 'neigh_op_bot_0')
// (14, 11, 'neigh_op_tnl_0')
// (14, 12, 'neigh_op_lft_0')
// (14, 13, 'local_g2_0')
// (14, 13, 'lutff_7/in_1')
// (14, 13, 'neigh_op_bnl_0')

wire n1759;
// (12, 11, 'neigh_op_tnr_1')
// (12, 12, 'neigh_op_rgt_1')
// (12, 13, 'neigh_op_bnr_1')
// (13, 11, 'neigh_op_top_1')
// (13, 12, 'local_g3_1')
// (13, 12, 'lutff_1/out')
// (13, 12, 'lutff_3/in_3')
// (13, 13, 'neigh_op_bot_1')
// (14, 11, 'neigh_op_tnl_1')
// (14, 12, 'neigh_op_lft_1')
// (14, 13, 'neigh_op_bnl_1')

wire n1760;
// (12, 11, 'neigh_op_tnr_3')
// (12, 12, 'neigh_op_rgt_3')
// (12, 13, 'neigh_op_bnr_3')
// (13, 11, 'neigh_op_top_3')
// (13, 12, 'lutff_3/out')
// (13, 12, 'sp4_r_v_b_39')
// (13, 13, 'local_g1_3')
// (13, 13, 'lutff_1/in_3')
// (13, 13, 'neigh_op_bot_3')
// (13, 13, 'sp4_r_v_b_26')
// (13, 14, 'sp4_r_v_b_15')
// (13, 15, 'sp4_r_v_b_2')
// (14, 11, 'neigh_op_tnl_3')
// (14, 11, 'sp4_v_t_39')
// (14, 12, 'neigh_op_lft_3')
// (14, 12, 'sp4_v_b_39')
// (14, 13, 'neigh_op_bnl_3')
// (14, 13, 'sp4_v_b_26')
// (14, 14, 'sp4_v_b_15')
// (14, 15, 'sp4_h_r_2')
// (14, 15, 'sp4_v_b_2')
// (15, 15, 'sp4_h_r_15')
// (16, 15, 'sp4_h_r_26')
// (17, 15, 'sp4_h_r_39')
// (18, 15, 'sp4_h_l_39')
// (18, 15, 'sp4_h_r_10')
// (19, 15, 'local_g1_7')
// (19, 15, 'ram/WDATA_10')
// (19, 15, 'sp4_h_r_23')
// (20, 15, 'sp4_h_r_34')
// (21, 15, 'sp4_h_r_47')
// (22, 15, 'sp4_h_l_47')

wire n1761;
// (12, 11, 'neigh_op_tnr_4')
// (12, 12, 'neigh_op_rgt_4')
// (12, 13, 'neigh_op_bnr_4')
// (13, 11, 'neigh_op_top_4')
// (13, 12, 'lutff_4/out')
// (13, 13, 'neigh_op_bot_4')
// (14, 11, 'neigh_op_tnl_4')
// (14, 12, 'neigh_op_lft_4')
// (14, 13, 'local_g3_4')
// (14, 13, 'lutff_6/in_1')
// (14, 13, 'neigh_op_bnl_4')

wire n1762;
// (12, 11, 'neigh_op_tnr_5')
// (12, 12, 'neigh_op_rgt_5')
// (12, 13, 'neigh_op_bnr_5')
// (13, 11, 'neigh_op_top_5')
// (13, 12, 'local_g1_5')
// (13, 12, 'lutff_3/in_1')
// (13, 12, 'lutff_5/out')
// (13, 13, 'neigh_op_bot_5')
// (14, 11, 'neigh_op_tnl_5')
// (14, 12, 'neigh_op_lft_5')
// (14, 13, 'neigh_op_bnl_5')

reg n1763 = 0;
// (12, 11, 'neigh_op_tnr_7')
// (12, 12, 'neigh_op_rgt_7')
// (12, 13, 'neigh_op_bnr_7')
// (13, 10, 'sp4_r_v_b_39')
// (13, 11, 'neigh_op_top_7')
// (13, 11, 'sp4_r_v_b_26')
// (13, 12, 'local_g0_7')
// (13, 12, 'lutff_4/in_3')
// (13, 12, 'lutff_6/in_3')
// (13, 12, 'lutff_7/out')
// (13, 12, 'sp4_r_v_b_15')
// (13, 13, 'neigh_op_bot_7')
// (13, 13, 'sp4_r_v_b_2')
// (14, 9, 'sp4_v_t_39')
// (14, 10, 'local_g3_7')
// (14, 10, 'lutff_7/in_1')
// (14, 10, 'sp4_v_b_39')
// (14, 11, 'neigh_op_tnl_7')
// (14, 11, 'sp4_v_b_26')
// (14, 12, 'neigh_op_lft_7')
// (14, 12, 'sp4_v_b_15')
// (14, 13, 'neigh_op_bnl_7')
// (14, 13, 'sp4_v_b_2')

wire n1764;
// (12, 11, 'sp12_h_r_0')
// (13, 10, 'neigh_op_tnr_6')
// (13, 11, 'neigh_op_rgt_6')
// (13, 11, 'sp12_h_r_3')
// (13, 12, 'neigh_op_bnr_6')
// (14, 10, 'neigh_op_top_6')
// (14, 11, 'lutff_6/out')
// (14, 11, 'sp12_h_r_4')
// (14, 12, 'neigh_op_bot_6')
// (15, 10, 'neigh_op_tnl_6')
// (15, 11, 'neigh_op_lft_6')
// (15, 11, 'sp12_h_r_7')
// (15, 12, 'neigh_op_bnl_6')
// (16, 11, 'sp12_h_r_8')
// (17, 11, 'local_g1_3')
// (17, 11, 'lutff_global/cen')
// (17, 11, 'sp12_h_r_11')
// (18, 11, 'sp12_h_r_12')
// (19, 11, 'sp12_h_r_15')
// (20, 11, 'sp12_h_r_16')
// (21, 11, 'sp12_h_r_19')
// (22, 11, 'sp12_h_r_20')
// (23, 11, 'sp12_h_r_23')
// (24, 11, 'sp12_h_l_23')

wire n1765;
// (12, 11, 'sp4_r_v_b_38')
// (12, 12, 'local_g1_3')
// (12, 12, 'lutff_1/in_1')
// (12, 12, 'sp4_r_v_b_27')
// (12, 13, 'sp4_r_v_b_14')
// (12, 14, 'sp4_r_v_b_3')
// (13, 10, 'sp4_v_t_38')
// (13, 11, 'sp4_v_b_38')
// (13, 12, 'sp4_v_b_27')
// (13, 13, 'sp4_v_b_14')
// (13, 14, 'sp4_h_r_3')
// (13, 14, 'sp4_v_b_3')
// (14, 14, 'sp4_h_r_14')
// (15, 11, 'sp4_r_v_b_43')
// (15, 12, 'sp4_r_v_b_30')
// (15, 13, 'neigh_op_tnr_3')
// (15, 13, 'sp4_r_v_b_19')
// (15, 14, 'neigh_op_rgt_3')
// (15, 14, 'sp4_h_r_27')
// (15, 14, 'sp4_r_v_b_6')
// (15, 15, 'local_g0_3')
// (15, 15, 'lutff_1/in_2')
// (15, 15, 'neigh_op_bnr_3')
// (16, 10, 'sp4_h_r_11')
// (16, 10, 'sp4_v_t_43')
// (16, 11, 'sp4_v_b_43')
// (16, 12, 'sp4_v_b_30')
// (16, 13, 'neigh_op_top_3')
// (16, 13, 'sp4_v_b_19')
// (16, 14, 'lutff_3/out')
// (16, 14, 'sp4_h_r_38')
// (16, 14, 'sp4_v_b_6')
// (16, 15, 'neigh_op_bot_3')
// (17, 10, 'local_g0_6')
// (17, 10, 'lutff_2/in_2')
// (17, 10, 'sp4_h_r_22')
// (17, 13, 'neigh_op_tnl_3')
// (17, 14, 'neigh_op_lft_3')
// (17, 14, 'sp4_h_l_38')
// (17, 15, 'neigh_op_bnl_3')
// (18, 10, 'sp4_h_r_35')
// (19, 10, 'sp4_h_r_46')
// (20, 10, 'sp4_h_l_46')

wire n1766;
// (12, 11, 'sp4_r_v_b_46')
// (12, 12, 'local_g2_3')
// (12, 12, 'lutff_2/in_1')
// (12, 12, 'sp4_r_v_b_35')
// (12, 13, 'sp4_r_v_b_22')
// (12, 14, 'sp4_r_v_b_11')
// (13, 10, 'sp4_v_t_46')
// (13, 11, 'sp4_v_b_46')
// (13, 12, 'sp4_v_b_35')
// (13, 13, 'sp4_v_b_22')
// (13, 14, 'sp4_h_r_11')
// (13, 14, 'sp4_v_b_11')
// (14, 14, 'local_g1_6')
// (14, 14, 'lutff_3/in_2')
// (14, 14, 'sp4_h_r_22')
// (15, 13, 'neigh_op_tnr_7')
// (15, 14, 'neigh_op_rgt_7')
// (15, 14, 'sp4_h_r_35')
// (15, 15, 'local_g1_7')
// (15, 15, 'lutff_2/in_2')
// (15, 15, 'neigh_op_bnr_7')
// (16, 8, 'sp4_r_v_b_39')
// (16, 9, 'sp4_r_v_b_26')
// (16, 10, 'sp4_r_v_b_15')
// (16, 11, 'sp4_r_v_b_2')
// (16, 12, 'sp4_r_v_b_39')
// (16, 13, 'neigh_op_top_7')
// (16, 13, 'sp4_r_v_b_26')
// (16, 14, 'local_g2_7')
// (16, 14, 'lutff_0/in_3')
// (16, 14, 'lutff_3/in_0')
// (16, 14, 'lutff_7/out')
// (16, 14, 'sp4_h_r_46')
// (16, 14, 'sp4_r_v_b_15')
// (16, 15, 'neigh_op_bot_7')
// (16, 15, 'sp4_r_v_b_2')
// (17, 7, 'sp4_v_t_39')
// (17, 8, 'sp4_v_b_39')
// (17, 9, 'sp4_v_b_26')
// (17, 10, 'local_g1_7')
// (17, 10, 'lutff_1/in_1')
// (17, 10, 'sp4_v_b_15')
// (17, 11, 'sp4_v_b_2')
// (17, 11, 'sp4_v_t_39')
// (17, 12, 'sp4_v_b_39')
// (17, 13, 'neigh_op_tnl_7')
// (17, 13, 'sp4_v_b_26')
// (17, 14, 'neigh_op_lft_7')
// (17, 14, 'sp4_h_l_46')
// (17, 14, 'sp4_v_b_15')
// (17, 15, 'neigh_op_bnl_7')
// (17, 15, 'sp4_v_b_2')

wire n1767;
// (12, 12, 'lutff_0/cout')
// (12, 12, 'lutff_1/in_3')

wire n1768;
// (12, 12, 'lutff_1/cout')
// (12, 12, 'lutff_2/in_3')

wire n1769;
// (12, 12, 'lutff_2/cout')
// (12, 12, 'lutff_3/in_3')

wire n1770;
// (12, 12, 'neigh_op_tnr_0')
// (12, 13, 'neigh_op_rgt_0')
// (12, 14, 'neigh_op_bnr_0')
// (13, 12, 'local_g1_0')
// (13, 12, 'lutff_5/in_2')
// (13, 12, 'neigh_op_top_0')
// (13, 13, 'lutff_0/out')
// (13, 14, 'neigh_op_bot_0')
// (14, 12, 'local_g3_0')
// (14, 12, 'lutff_0/in_3')
// (14, 12, 'lutff_2/in_3')
// (14, 12, 'lutff_3/in_0')
// (14, 12, 'lutff_4/in_1')
// (14, 12, 'lutff_6/in_1')
// (14, 12, 'lutff_7/in_0')
// (14, 12, 'neigh_op_tnl_0')
// (14, 13, 'local_g1_0')
// (14, 13, 'lutff_3/in_2')
// (14, 13, 'lutff_4/in_3')
// (14, 13, 'neigh_op_lft_0')
// (14, 14, 'local_g3_0')
// (14, 14, 'lutff_0/in_1')
// (14, 14, 'lutff_1/in_2')
// (14, 14, 'lutff_5/in_0')
// (14, 14, 'neigh_op_bnl_0')

reg n1771 = 0;
// (12, 12, 'neigh_op_tnr_1')
// (12, 13, 'local_g2_1')
// (12, 13, 'lutff_3/in_2')
// (12, 13, 'neigh_op_rgt_1')
// (12, 14, 'neigh_op_bnr_1')
// (13, 12, 'neigh_op_top_1')
// (13, 13, 'lutff_1/out')
// (13, 14, 'neigh_op_bot_1')
// (14, 12, 'neigh_op_tnl_1')
// (14, 13, 'neigh_op_lft_1')
// (14, 14, 'neigh_op_bnl_1')

wire n1772;
// (12, 12, 'neigh_op_tnr_2')
// (12, 13, 'neigh_op_rgt_2')
// (12, 14, 'neigh_op_bnr_2')
// (13, 12, 'local_g0_2')
// (13, 12, 'lutff_0/in_2')
// (13, 12, 'lutff_1/in_3')
// (13, 12, 'lutff_5/in_1')
// (13, 12, 'neigh_op_top_2')
// (13, 13, 'lutff_2/out')
// (13, 14, 'local_g0_2')
// (13, 14, 'lutff_3/in_1')
// (13, 14, 'lutff_4/in_2')
// (13, 14, 'neigh_op_bot_2')
// (14, 12, 'local_g3_2')
// (14, 12, 'lutff_3/in_2')
// (14, 12, 'lutff_4/in_3')
// (14, 12, 'lutff_6/in_3')
// (14, 12, 'neigh_op_tnl_2')
// (14, 13, 'local_g1_2')
// (14, 13, 'lutff_1/in_2')
// (14, 13, 'lutff_4/in_1')
// (14, 13, 'lutff_5/in_0')
// (14, 13, 'lutff_6/in_3')
// (14, 13, 'neigh_op_lft_2')
// (14, 14, 'local_g2_2')
// (14, 14, 'lutff_2/in_0')
// (14, 14, 'lutff_7/in_3')
// (14, 14, 'neigh_op_bnl_2')

reg n1773 = 0;
// (12, 12, 'neigh_op_tnr_3')
// (12, 13, 'local_g3_3')
// (12, 13, 'lutff_7/in_1')
// (12, 13, 'neigh_op_rgt_3')
// (12, 14, 'neigh_op_bnr_3')
// (13, 12, 'neigh_op_top_3')
// (13, 13, 'lutff_3/out')
// (13, 14, 'neigh_op_bot_3')
// (14, 12, 'neigh_op_tnl_3')
// (14, 13, 'neigh_op_lft_3')
// (14, 14, 'neigh_op_bnl_3')

reg n1774 = 0;
// (12, 12, 'neigh_op_tnr_4')
// (12, 13, 'local_g3_4')
// (12, 13, 'lutff_5/in_2')
// (12, 13, 'neigh_op_rgt_4')
// (12, 14, 'neigh_op_bnr_4')
// (13, 12, 'neigh_op_top_4')
// (13, 13, 'lutff_4/out')
// (13, 14, 'neigh_op_bot_4')
// (14, 12, 'neigh_op_tnl_4')
// (14, 13, 'neigh_op_lft_4')
// (14, 14, 'neigh_op_bnl_4')

reg n1775 = 0;
// (12, 12, 'neigh_op_tnr_5')
// (12, 13, 'local_g2_5')
// (12, 13, 'lutff_4/in_3')
// (12, 13, 'neigh_op_rgt_5')
// (12, 14, 'neigh_op_bnr_5')
// (13, 12, 'neigh_op_top_5')
// (13, 13, 'lutff_5/out')
// (13, 14, 'neigh_op_bot_5')
// (14, 12, 'neigh_op_tnl_5')
// (14, 13, 'neigh_op_lft_5')
// (14, 14, 'neigh_op_bnl_5')

reg n1776 = 0;
// (12, 12, 'neigh_op_tnr_6')
// (12, 13, 'local_g3_6')
// (12, 13, 'lutff_1/in_0')
// (12, 13, 'neigh_op_rgt_6')
// (12, 14, 'neigh_op_bnr_6')
// (13, 12, 'neigh_op_top_6')
// (13, 13, 'lutff_6/out')
// (13, 14, 'neigh_op_bot_6')
// (14, 12, 'neigh_op_tnl_6')
// (14, 13, 'neigh_op_lft_6')
// (14, 14, 'neigh_op_bnl_6')

reg n1777 = 0;
// (12, 12, 'neigh_op_tnr_7')
// (12, 13, 'local_g2_7')
// (12, 13, 'lutff_6/in_1')
// (12, 13, 'neigh_op_rgt_7')
// (12, 14, 'neigh_op_bnr_7')
// (13, 12, 'neigh_op_top_7')
// (13, 13, 'lutff_7/out')
// (13, 14, 'neigh_op_bot_7')
// (14, 12, 'neigh_op_tnl_7')
// (14, 13, 'neigh_op_lft_7')
// (14, 14, 'neigh_op_bnl_7')

wire n1778;
// (12, 12, 'sp4_h_r_1')
// (13, 12, 'sp4_h_r_12')
// (14, 11, 'neigh_op_tnr_2')
// (14, 12, 'neigh_op_rgt_2')
// (14, 12, 'sp4_h_r_25')
// (14, 13, 'neigh_op_bnr_2')
// (15, 11, 'neigh_op_top_2')
// (15, 12, 'local_g2_4')
// (15, 12, 'lutff_2/out')
// (15, 12, 'lutff_4/in_2')
// (15, 12, 'sp4_h_r_36')
// (15, 13, 'neigh_op_bot_2')
// (16, 11, 'neigh_op_tnl_2')
// (16, 12, 'neigh_op_lft_2')
// (16, 12, 'sp4_h_l_36')
// (16, 13, 'neigh_op_bnl_2')

wire n1779;
// (12, 12, 'sp4_r_v_b_39')
// (12, 13, 'sp4_r_v_b_26')
// (12, 14, 'local_g2_7')
// (12, 14, 'lutff_5/in_0')
// (12, 14, 'sp4_r_v_b_15')
// (12, 15, 'sp4_r_v_b_2')
// (13, 11, 'sp4_v_t_39')
// (13, 12, 'sp4_v_b_39')
// (13, 13, 'sp4_v_b_26')
// (13, 14, 'neigh_op_tnr_2')
// (13, 14, 'sp4_v_b_15')
// (13, 15, 'neigh_op_rgt_2')
// (13, 15, 'sp4_h_r_9')
// (13, 15, 'sp4_v_b_2')
// (13, 16, 'neigh_op_bnr_2')
// (14, 14, 'neigh_op_top_2')
// (14, 15, 'lutff_2/out')
// (14, 15, 'sp4_h_r_20')
// (14, 16, 'neigh_op_bot_2')
// (15, 14, 'neigh_op_tnl_2')
// (15, 15, 'neigh_op_lft_2')
// (15, 15, 'sp4_h_r_33')
// (15, 16, 'neigh_op_bnl_2')
// (16, 15, 'sp4_h_r_44')
// (17, 15, 'sp4_h_l_44')

reg n1780 = 0;
// (12, 12, 'sp4_r_v_b_41')
// (12, 13, 'sp4_r_v_b_28')
// (12, 14, 'local_g3_1')
// (12, 14, 'lutff_5/in_1')
// (12, 14, 'sp4_r_v_b_17')
// (12, 15, 'sp4_r_v_b_4')
// (12, 16, 'sp4_r_v_b_36')
// (12, 17, 'neigh_op_tnr_6')
// (12, 17, 'sp4_r_v_b_25')
// (12, 18, 'neigh_op_rgt_6')
// (12, 18, 'sp4_r_v_b_12')
// (12, 19, 'neigh_op_bnr_6')
// (12, 19, 'sp4_r_v_b_1')
// (13, 11, 'sp4_v_t_41')
// (13, 12, 'sp4_v_b_41')
// (13, 13, 'sp4_v_b_28')
// (13, 14, 'sp4_v_b_17')
// (13, 15, 'sp4_v_b_4')
// (13, 15, 'sp4_v_t_36')
// (13, 16, 'sp4_v_b_36')
// (13, 17, 'local_g1_6')
// (13, 17, 'lutff_5/in_2')
// (13, 17, 'neigh_op_top_6')
// (13, 17, 'sp4_r_v_b_40')
// (13, 17, 'sp4_v_b_25')
// (13, 18, 'local_g0_6')
// (13, 18, 'lutff_6/in_2')
// (13, 18, 'lutff_6/out')
// (13, 18, 'sp4_r_v_b_29')
// (13, 18, 'sp4_v_b_12')
// (13, 19, 'neigh_op_bot_6')
// (13, 19, 'sp4_r_v_b_16')
// (13, 19, 'sp4_v_b_1')
// (13, 20, 'sp4_r_v_b_5')
// (14, 16, 'sp4_h_r_10')
// (14, 16, 'sp4_v_t_40')
// (14, 17, 'neigh_op_tnl_6')
// (14, 17, 'sp4_v_b_40')
// (14, 18, 'neigh_op_lft_6')
// (14, 18, 'sp4_v_b_29')
// (14, 19, 'neigh_op_bnl_6')
// (14, 19, 'sp4_v_b_16')
// (14, 20, 'sp4_v_b_5')
// (15, 16, 'sp4_h_r_23')
// (16, 16, 'sp4_h_r_34')
// (17, 16, 'sp4_h_r_47')
// (18, 16, 'sp4_h_l_47')
// (18, 16, 'sp4_h_r_10')
// (19, 16, 'local_g1_7')
// (19, 16, 'ram/WADDR_3')
// (19, 16, 'sp4_h_r_23')
// (20, 16, 'sp4_h_r_34')
// (21, 16, 'sp4_h_r_47')
// (22, 16, 'sp4_h_l_47')

wire n1781;
// (12, 12, 'sp4_r_v_b_43')
// (12, 13, 'sp4_r_v_b_30')
// (12, 14, 'local_g3_3')
// (12, 14, 'lutff_5/in_3')
// (12, 14, 'sp4_r_v_b_19')
// (12, 15, 'sp4_r_v_b_6')
// (13, 11, 'sp4_v_t_43')
// (13, 12, 'sp4_v_b_43')
// (13, 13, 'sp4_v_b_30')
// (13, 14, 'neigh_op_tnr_6')
// (13, 14, 'sp4_v_b_19')
// (13, 15, 'neigh_op_rgt_6')
// (13, 15, 'sp4_h_r_1')
// (13, 15, 'sp4_v_b_6')
// (13, 16, 'neigh_op_bnr_6')
// (14, 14, 'neigh_op_top_6')
// (14, 15, 'lutff_6/out')
// (14, 15, 'sp4_h_r_12')
// (14, 16, 'neigh_op_bot_6')
// (15, 14, 'neigh_op_tnl_6')
// (15, 15, 'neigh_op_lft_6')
// (15, 15, 'sp4_h_r_25')
// (15, 16, 'neigh_op_bnl_6')
// (16, 15, 'sp4_h_r_36')
// (17, 15, 'sp4_h_l_36')

wire n1782;
// (12, 13, 'local_g0_3')
// (12, 13, 'lutff_3/in_0')
// (12, 13, 'sp4_h_r_3')
// (13, 13, 'sp4_h_r_14')
// (14, 13, 'sp4_h_r_27')
// (15, 13, 'sp4_h_r_38')
// (16, 13, 'sp4_h_l_38')
// (16, 13, 'sp4_h_r_3')
// (17, 13, 'sp4_h_r_14')
// (18, 13, 'sp4_h_r_27')
// (18, 14, 'neigh_op_tnr_5')
// (18, 15, 'neigh_op_rgt_5')
// (18, 16, 'neigh_op_bnr_5')
// (19, 13, 'sp4_h_r_38')
// (19, 14, 'neigh_op_top_5')
// (19, 14, 'sp4_r_v_b_38')
// (19, 15, 'ram/RDATA_10')
// (19, 15, 'sp4_r_v_b_27')
// (19, 16, 'neigh_op_bot_5')
// (19, 16, 'sp4_r_v_b_14')
// (19, 17, 'sp4_r_v_b_3')
// (20, 13, 'sp4_h_l_38')
// (20, 13, 'sp4_v_t_38')
// (20, 14, 'neigh_op_tnl_5')
// (20, 14, 'sp4_v_b_38')
// (20, 15, 'neigh_op_lft_5')
// (20, 15, 'sp4_v_b_27')
// (20, 16, 'neigh_op_bnl_5')
// (20, 16, 'sp4_v_b_14')
// (20, 17, 'sp4_v_b_3')

reg n1783 = 0;
// (12, 13, 'local_g3_5')
// (12, 13, 'lutff_1/in_3')
// (12, 13, 'lutff_3/in_3')
// (12, 13, 'lutff_4/in_2')
// (12, 13, 'lutff_5/in_3')
// (12, 13, 'lutff_6/in_0')
// (12, 13, 'lutff_7/in_3')
// (12, 13, 'sp4_r_v_b_45')
// (12, 14, 'sp4_r_v_b_32')
// (12, 15, 'neigh_op_tnr_4')
// (12, 15, 'sp4_r_v_b_21')
// (12, 16, 'local_g2_4')
// (12, 16, 'lutff_0/in_0')
// (12, 16, 'lutff_1/in_3')
// (12, 16, 'neigh_op_rgt_4')
// (12, 16, 'sp4_r_v_b_8')
// (12, 17, 'neigh_op_bnr_4')
// (13, 12, 'sp4_v_t_45')
// (13, 13, 'sp4_v_b_45')
// (13, 14, 'sp4_v_b_32')
// (13, 15, 'neigh_op_top_4')
// (13, 15, 'sp4_v_b_21')
// (13, 16, 'lutff_4/out')
// (13, 16, 'sp4_v_b_8')
// (13, 17, 'neigh_op_bot_4')
// (14, 15, 'neigh_op_tnl_4')
// (14, 16, 'neigh_op_lft_4')
// (14, 17, 'neigh_op_bnl_4')

wire n1784;
// (12, 13, 'neigh_op_tnr_0')
// (12, 14, 'neigh_op_rgt_0')
// (12, 15, 'neigh_op_bnr_0')
// (13, 13, 'neigh_op_top_0')
// (13, 14, 'lutff_0/out')
// (13, 15, 'neigh_op_bot_0')
// (14, 13, 'neigh_op_tnl_0')
// (14, 14, 'local_g1_0')
// (14, 14, 'lutff_7/in_0')
// (14, 14, 'neigh_op_lft_0')
// (14, 15, 'neigh_op_bnl_0')

wire n1785;
// (12, 13, 'neigh_op_tnr_3')
// (12, 14, 'neigh_op_rgt_3')
// (12, 15, 'neigh_op_bnr_3')
// (13, 13, 'neigh_op_top_3')
// (13, 14, 'local_g0_3')
// (13, 14, 'lutff_3/out')
// (13, 14, 'lutff_4/in_3')
// (13, 15, 'neigh_op_bot_3')
// (14, 13, 'neigh_op_tnl_3')
// (14, 14, 'neigh_op_lft_3')
// (14, 15, 'neigh_op_bnl_3')

wire n1786;
// (12, 13, 'neigh_op_tnr_4')
// (12, 14, 'neigh_op_rgt_4')
// (12, 15, 'neigh_op_bnr_4')
// (13, 13, 'neigh_op_top_4')
// (13, 13, 'sp4_r_v_b_36')
// (13, 14, 'lutff_4/out')
// (13, 14, 'sp4_r_v_b_25')
// (13, 15, 'local_g1_4')
// (13, 15, 'lutff_6/in_3')
// (13, 15, 'neigh_op_bot_4')
// (13, 15, 'sp4_r_v_b_12')
// (13, 16, 'sp4_r_v_b_1')
// (14, 12, 'sp4_v_t_36')
// (14, 13, 'neigh_op_tnl_4')
// (14, 13, 'sp4_v_b_36')
// (14, 14, 'neigh_op_lft_4')
// (14, 14, 'sp4_v_b_25')
// (14, 15, 'neigh_op_bnl_4')
// (14, 15, 'sp4_v_b_12')
// (14, 16, 'sp4_h_r_7')
// (14, 16, 'sp4_v_b_1')
// (15, 16, 'sp4_h_r_18')
// (16, 16, 'sp4_h_r_31')
// (17, 16, 'sp4_h_r_42')
// (18, 16, 'sp4_h_l_42')
// (18, 16, 'sp4_h_r_3')
// (19, 16, 'local_g0_6')
// (19, 16, 'ram/WDATA_0')
// (19, 16, 'sp4_h_r_14')
// (20, 16, 'sp4_h_r_27')
// (21, 16, 'sp4_h_r_38')
// (22, 16, 'sp4_h_l_38')

wire n1787;
// (12, 13, 'neigh_op_tnr_5')
// (12, 14, 'neigh_op_rgt_5')
// (12, 15, 'neigh_op_bnr_5')
// (13, 13, 'neigh_op_top_5')
// (13, 14, 'lutff_5/out')
// (13, 15, 'local_g1_5')
// (13, 15, 'lutff_1/in_1')
// (13, 15, 'neigh_op_bot_5')
// (14, 13, 'neigh_op_tnl_5')
// (14, 14, 'neigh_op_lft_5')
// (14, 15, 'neigh_op_bnl_5')

wire n1788;
// (12, 13, 'neigh_op_tnr_7')
// (12, 14, 'neigh_op_rgt_7')
// (12, 15, 'neigh_op_bnr_7')
// (13, 13, 'neigh_op_top_7')
// (13, 14, 'lutff_7/out')
// (13, 15, 'local_g1_7')
// (13, 15, 'lutff_2/in_2')
// (13, 15, 'neigh_op_bot_7')
// (14, 13, 'neigh_op_tnl_7')
// (14, 14, 'neigh_op_lft_7')
// (14, 15, 'neigh_op_bnl_7')

reg n1789 = 0;
// (12, 13, 'sp4_h_r_8')
// (13, 12, 'neigh_op_tnr_0')
// (13, 13, 'neigh_op_rgt_0')
// (13, 13, 'sp4_h_r_21')
// (13, 13, 'sp4_h_r_5')
// (13, 14, 'neigh_op_bnr_0')
// (14, 1, 'sp12_v_t_23')
// (14, 2, 'sp12_v_b_23')
// (14, 3, 'sp12_v_b_20')
// (14, 4, 'sp12_v_b_19')
// (14, 5, 'sp12_v_b_16')
// (14, 6, 'sp12_v_b_15')
// (14, 7, 'sp12_v_b_12')
// (14, 8, 'sp12_v_b_11')
// (14, 9, 'local_g2_0')
// (14, 9, 'lutff_2/in_2')
// (14, 9, 'sp12_v_b_8')
// (14, 10, 'sp12_v_b_7')
// (14, 11, 'sp12_v_b_4')
// (14, 12, 'neigh_op_top_0')
// (14, 12, 'sp12_v_b_3')
// (14, 13, 'lutff_0/out')
// (14, 13, 'sp12_v_b_0')
// (14, 13, 'sp4_h_r_0')
// (14, 13, 'sp4_h_r_16')
// (14, 13, 'sp4_h_r_32')
// (14, 14, 'neigh_op_bot_0')
// (15, 12, 'neigh_op_tnl_0')
// (15, 13, 'neigh_op_lft_0')
// (15, 13, 'sp4_h_r_13')
// (15, 13, 'sp4_h_r_29')
// (15, 13, 'sp4_h_r_45')
// (15, 14, 'neigh_op_bnl_0')
// (16, 6, 'sp4_r_v_b_39')
// (16, 7, 'local_g1_2')
// (16, 7, 'lutff_2/in_1')
// (16, 7, 'sp4_r_v_b_26')
// (16, 8, 'local_g2_7')
// (16, 8, 'lutff_2/in_1')
// (16, 8, 'sp4_r_v_b_15')
// (16, 9, 'sp4_r_v_b_2')
// (16, 10, 'sp4_r_v_b_46')
// (16, 11, 'sp4_r_v_b_35')
// (16, 12, 'sp4_r_v_b_22')
// (16, 13, 'local_g2_0')
// (16, 13, 'lutff_6/in_0')
// (16, 13, 'sp4_h_l_45')
// (16, 13, 'sp4_h_r_11')
// (16, 13, 'sp4_h_r_24')
// (16, 13, 'sp4_h_r_40')
// (16, 13, 'sp4_r_v_b_11')
// (17, 5, 'sp4_v_t_39')
// (17, 6, 'sp4_r_v_b_38')
// (17, 6, 'sp4_v_b_39')
// (17, 7, 'sp4_r_v_b_27')
// (17, 7, 'sp4_v_b_26')
// (17, 8, 'sp4_r_v_b_14')
// (17, 8, 'sp4_v_b_15')
// (17, 9, 'local_g0_4')
// (17, 9, 'lutff_1/in_1')
// (17, 9, 'sp4_h_r_4')
// (17, 9, 'sp4_r_v_b_3')
// (17, 9, 'sp4_v_b_2')
// (17, 9, 'sp4_v_t_46')
// (17, 10, 'sp4_r_v_b_37')
// (17, 10, 'sp4_v_b_46')
// (17, 11, 'sp4_r_v_b_24')
// (17, 11, 'sp4_v_b_35')
// (17, 12, 'sp4_r_v_b_13')
// (17, 12, 'sp4_v_b_22')
// (17, 13, 'sp4_h_l_40')
// (17, 13, 'sp4_h_r_22')
// (17, 13, 'sp4_h_r_37')
// (17, 13, 'sp4_h_r_5')
// (17, 13, 'sp4_r_v_b_0')
// (17, 13, 'sp4_v_b_11')
// (18, 5, 'sp4_v_t_38')
// (18, 6, 'sp4_v_b_38')
// (18, 7, 'local_g2_3')
// (18, 7, 'lutff_5/in_0')
// (18, 7, 'sp4_v_b_27')
// (18, 8, 'local_g1_6')
// (18, 8, 'lutff_0/in_3')
// (18, 8, 'sp4_v_b_14')
// (18, 9, 'sp4_h_r_17')
// (18, 9, 'sp4_v_b_3')
// (18, 9, 'sp4_v_t_37')
// (18, 10, 'sp4_v_b_37')
// (18, 11, 'sp4_v_b_24')
// (18, 12, 'sp4_v_b_13')
// (18, 13, 'sp4_h_l_37')
// (18, 13, 'sp4_h_r_16')
// (18, 13, 'sp4_h_r_35')
// (18, 13, 'sp4_v_b_0')
// (19, 9, 'sp4_h_r_28')
// (19, 10, 'sp4_r_v_b_40')
// (19, 11, 'sp4_r_v_b_29')
// (19, 12, 'sp4_r_v_b_16')
// (19, 13, 'sp4_h_r_29')
// (19, 13, 'sp4_h_r_46')
// (19, 13, 'sp4_r_v_b_5')
// (20, 9, 'sp4_h_r_41')
// (20, 9, 'sp4_v_t_40')
// (20, 10, 'local_g3_0')
// (20, 10, 'lutff_7/in_0')
// (20, 10, 'sp4_r_v_b_40')
// (20, 10, 'sp4_v_b_40')
// (20, 11, 'sp4_r_v_b_29')
// (20, 11, 'sp4_v_b_29')
// (20, 12, 'sp4_r_v_b_16')
// (20, 12, 'sp4_v_b_16')
// (20, 13, 'sp4_h_l_46')
// (20, 13, 'sp4_h_r_40')
// (20, 13, 'sp4_r_v_b_5')
// (20, 13, 'sp4_v_b_5')
// (21, 9, 'sp4_h_l_41')
// (21, 9, 'sp4_v_t_40')
// (21, 10, 'sp4_v_b_40')
// (21, 11, 'local_g2_5')
// (21, 11, 'lutff_3/in_2')
// (21, 11, 'sp4_v_b_29')
// (21, 12, 'sp4_v_b_16')
// (21, 13, 'sp4_h_l_40')
// (21, 13, 'sp4_v_b_5')

reg n1790 = 0;
// (12, 13, 'sp4_r_v_b_40')
// (12, 14, 'sp4_r_v_b_29')
// (12, 15, 'sp4_r_v_b_16')
// (12, 16, 'sp4_r_v_b_5')
// (13, 12, 'sp4_v_t_40')
// (13, 13, 'local_g2_0')
// (13, 13, 'lutff_0/in_2')
// (13, 13, 'lutff_2/in_0')
// (13, 13, 'sp4_v_b_40')
// (13, 14, 'local_g2_5')
// (13, 14, 'lutff_2/in_3')
// (13, 14, 'sp4_v_b_29')
// (13, 15, 'sp4_v_b_16')
// (13, 16, 'sp4_h_r_0')
// (13, 16, 'sp4_v_b_5')
// (14, 13, 'sp4_r_v_b_45')
// (14, 14, 'sp4_r_v_b_32')
// (14, 15, 'neigh_op_tnr_4')
// (14, 15, 'sp4_r_v_b_21')
// (14, 16, 'neigh_op_rgt_4')
// (14, 16, 'sp4_h_r_13')
// (14, 16, 'sp4_r_v_b_8')
// (14, 17, 'neigh_op_bnr_4')
// (15, 12, 'sp4_v_t_45')
// (15, 13, 'sp4_r_v_b_44')
// (15, 13, 'sp4_v_b_45')
// (15, 14, 'local_g3_0')
// (15, 14, 'lutff_5/in_2')
// (15, 14, 'sp4_r_v_b_33')
// (15, 14, 'sp4_v_b_32')
// (15, 15, 'local_g0_4')
// (15, 15, 'local_g1_4')
// (15, 15, 'lutff_4/in_0')
// (15, 15, 'lutff_5/in_0')
// (15, 15, 'neigh_op_top_4')
// (15, 15, 'sp4_r_v_b_20')
// (15, 15, 'sp4_v_b_21')
// (15, 16, 'local_g1_4')
// (15, 16, 'local_g2_4')
// (15, 16, 'lutff_0/in_2')
// (15, 16, 'lutff_3/in_1')
// (15, 16, 'lutff_4/in_2')
// (15, 16, 'lutff_4/out')
// (15, 16, 'lutff_7/in_0')
// (15, 16, 'sp4_h_r_24')
// (15, 16, 'sp4_r_v_b_9')
// (15, 16, 'sp4_v_b_8')
// (15, 17, 'neigh_op_bot_4')
// (16, 12, 'local_g0_2')
// (16, 12, 'lutff_0/in_0')
// (16, 12, 'lutff_6/in_0')
// (16, 12, 'sp4_h_r_2')
// (16, 12, 'sp4_v_t_44')
// (16, 13, 'local_g2_4')
// (16, 13, 'lutff_7/in_3')
// (16, 13, 'sp4_v_b_44')
// (16, 14, 'local_g3_1')
// (16, 14, 'lutff_5/in_1')
// (16, 14, 'sp4_v_b_33')
// (16, 15, 'neigh_op_tnl_4')
// (16, 15, 'sp4_v_b_20')
// (16, 16, 'neigh_op_lft_4')
// (16, 16, 'sp4_h_r_37')
// (16, 16, 'sp4_v_b_9')
// (16, 17, 'neigh_op_bnl_4')
// (17, 12, 'sp4_h_r_15')
// (17, 16, 'sp4_h_l_37')
// (18, 12, 'sp4_h_r_26')
// (19, 12, 'sp4_h_r_39')
// (20, 12, 'sp4_h_l_39')

wire n1791;
// (12, 13, 'sp4_r_v_b_46')
// (12, 14, 'sp4_r_v_b_35')
// (12, 15, 'sp4_r_v_b_22')
// (12, 16, 'local_g2_3')
// (12, 16, 'lutff_0/in_1')
// (12, 16, 'sp4_r_v_b_11')
// (13, 12, 'sp4_v_t_46')
// (13, 13, 'sp4_v_b_46')
// (13, 14, 'sp4_v_b_35')
// (13, 15, 'sp4_v_b_22')
// (13, 16, 'sp4_h_r_6')
// (13, 16, 'sp4_v_b_11')
// (14, 16, 'sp4_h_r_19')
// (15, 16, 'sp4_h_r_30')
// (16, 16, 'sp4_h_r_43')
// (17, 16, 'sp4_h_l_43')
// (17, 16, 'sp4_h_r_10')
// (18, 15, 'neigh_op_tnr_1')
// (18, 16, 'neigh_op_rgt_1')
// (18, 16, 'sp4_h_r_23')
// (18, 17, 'neigh_op_bnr_1')
// (19, 15, 'neigh_op_top_1')
// (19, 16, 'ram/RDATA_6')
// (19, 16, 'sp4_h_r_34')
// (19, 17, 'neigh_op_bot_1')
// (20, 15, 'neigh_op_tnl_1')
// (20, 16, 'neigh_op_lft_1')
// (20, 16, 'sp4_h_r_47')
// (20, 17, 'neigh_op_bnl_1')
// (21, 16, 'sp4_h_l_47')

wire n1792;
// (12, 14, 'local_g2_3')
// (12, 14, 'lutff_5/in_2')
// (12, 14, 'neigh_op_tnr_3')
// (12, 15, 'neigh_op_rgt_3')
// (12, 16, 'neigh_op_bnr_3')
// (13, 14, 'neigh_op_top_3')
// (13, 15, 'lutff_3/out')
// (13, 15, 'sp4_h_r_6')
// (13, 16, 'neigh_op_bot_3')
// (14, 14, 'neigh_op_tnl_3')
// (14, 15, 'neigh_op_lft_3')
// (14, 15, 'sp4_h_r_19')
// (14, 16, 'neigh_op_bnl_3')
// (15, 15, 'sp4_h_r_30')
// (16, 15, 'sp4_h_r_43')
// (17, 15, 'sp4_h_l_43')
// (17, 15, 'sp4_h_r_9')
// (18, 15, 'sp4_h_r_20')
// (19, 15, 'local_g3_1')
// (19, 15, 'ram/RADDR_3')
// (19, 15, 'sp4_h_r_33')
// (20, 15, 'sp4_h_r_44')
// (21, 15, 'sp4_h_l_44')

wire n1793;
// (12, 14, 'lutff_1/cout')
// (12, 14, 'lutff_2/in_3')

wire n1794;
// (12, 14, 'lutff_2/cout')
// (12, 14, 'lutff_3/in_3')

wire n1795;
// (12, 14, 'neigh_op_tnr_1')
// (12, 15, 'neigh_op_rgt_1')
// (12, 16, 'neigh_op_bnr_1')
// (13, 14, 'neigh_op_top_1')
// (13, 15, 'lutff_1/out')
// (13, 15, 'sp4_h_r_2')
// (13, 16, 'neigh_op_bot_1')
// (14, 14, 'neigh_op_tnl_1')
// (14, 15, 'local_g1_1')
// (14, 15, 'lutff_2/in_2')
// (14, 15, 'neigh_op_lft_1')
// (14, 15, 'sp4_h_r_15')
// (14, 16, 'neigh_op_bnl_1')
// (15, 15, 'sp4_h_r_26')
// (16, 15, 'sp4_h_r_39')
// (17, 15, 'sp4_h_l_39')
// (17, 15, 'sp4_h_r_5')
// (18, 15, 'sp4_h_r_16')
// (19, 15, 'local_g3_5')
// (19, 15, 'ram/RADDR_1')
// (19, 15, 'sp4_h_r_29')
// (20, 15, 'sp4_h_r_40')
// (21, 15, 'sp4_h_l_40')

wire n1796;
// (12, 14, 'neigh_op_tnr_2')
// (12, 15, 'neigh_op_rgt_2')
// (12, 16, 'neigh_op_bnr_2')
// (13, 14, 'neigh_op_top_2')
// (13, 15, 'lutff_2/out')
// (13, 15, 'sp4_h_r_4')
// (13, 16, 'neigh_op_bot_2')
// (14, 14, 'neigh_op_tnl_2')
// (14, 15, 'local_g1_2')
// (14, 15, 'lutff_7/in_0')
// (14, 15, 'neigh_op_lft_2')
// (14, 15, 'sp4_h_r_17')
// (14, 16, 'neigh_op_bnl_2')
// (15, 15, 'sp4_h_r_28')
// (16, 15, 'sp4_h_r_41')
// (17, 15, 'sp4_h_l_41')
// (17, 15, 'sp4_h_r_4')
// (18, 15, 'sp4_h_r_17')
// (19, 15, 'local_g3_4')
// (19, 15, 'ram/RADDR_2')
// (19, 15, 'sp4_h_r_28')
// (20, 15, 'sp4_h_r_41')
// (21, 15, 'sp4_h_l_41')

wire n1797;
// (12, 14, 'neigh_op_tnr_4')
// (12, 15, 'neigh_op_rgt_4')
// (12, 16, 'neigh_op_bnr_4')
// (13, 14, 'neigh_op_top_4')
// (13, 15, 'lutff_4/out')
// (13, 15, 'sp12_h_r_0')
// (13, 16, 'neigh_op_bot_4')
// (14, 14, 'neigh_op_tnl_4')
// (14, 15, 'local_g0_4')
// (14, 15, 'lutff_6/in_0')
// (14, 15, 'neigh_op_lft_4')
// (14, 15, 'sp12_h_r_3')
// (14, 16, 'neigh_op_bnl_4')
// (15, 15, 'sp12_h_r_4')
// (16, 15, 'sp12_h_r_7')
// (17, 15, 'sp12_h_r_8')
// (18, 15, 'sp12_h_r_11')
// (19, 15, 'local_g1_4')
// (19, 15, 'ram/RADDR_4')
// (19, 15, 'sp12_h_r_12')
// (20, 15, 'sp12_h_r_15')
// (21, 15, 'sp12_h_r_16')
// (22, 15, 'sp12_h_r_19')
// (23, 15, 'sp12_h_r_20')
// (24, 15, 'sp12_h_r_23')
// (25, 15, 'sp12_h_l_23')

wire n1798;
// (12, 14, 'neigh_op_tnr_5')
// (12, 15, 'neigh_op_rgt_5')
// (12, 15, 'sp12_h_r_1')
// (12, 16, 'neigh_op_bnr_5')
// (13, 14, 'neigh_op_top_5')
// (13, 15, 'lutff_5/out')
// (13, 15, 'sp12_h_r_2')
// (13, 16, 'neigh_op_bot_5')
// (14, 14, 'neigh_op_tnl_5')
// (14, 15, 'local_g0_5')
// (14, 15, 'lutff_7/in_2')
// (14, 15, 'neigh_op_lft_5')
// (14, 15, 'sp12_h_r_5')
// (14, 16, 'neigh_op_bnl_5')
// (15, 15, 'sp12_h_r_6')
// (16, 15, 'sp12_h_r_9')
// (17, 15, 'sp12_h_r_10')
// (18, 15, 'sp12_h_r_13')
// (19, 15, 'local_g0_6')
// (19, 15, 'ram/RADDR_5')
// (19, 15, 'sp12_h_r_14')
// (20, 15, 'sp12_h_r_17')
// (21, 15, 'sp12_h_r_18')
// (22, 15, 'sp12_h_r_21')
// (23, 15, 'sp12_h_r_22')
// (24, 15, 'sp12_h_l_22')

reg n1799 = 0;
// (12, 14, 'neigh_op_tnr_6')
// (12, 15, 'neigh_op_rgt_6')
// (12, 16, 'local_g1_6')
// (12, 16, 'lutff_1/in_0')
// (12, 16, 'neigh_op_bnr_6')
// (13, 14, 'neigh_op_top_6')
// (13, 15, 'lutff_6/out')
// (13, 16, 'neigh_op_bot_6')
// (14, 14, 'neigh_op_tnl_6')
// (14, 15, 'neigh_op_lft_6')
// (14, 16, 'neigh_op_bnl_6')

reg n1800 = 0;
// (12, 14, 'neigh_op_tnr_7')
// (12, 15, 'neigh_op_rgt_7')
// (12, 16, 'local_g0_7')
// (12, 16, 'lutff_0/in_3')
// (12, 16, 'neigh_op_bnr_7')
// (13, 14, 'neigh_op_top_7')
// (13, 15, 'lutff_7/out')
// (13, 16, 'neigh_op_bot_7')
// (14, 14, 'neigh_op_tnl_7')
// (14, 15, 'neigh_op_lft_7')
// (14, 16, 'neigh_op_bnl_7')

wire n1801;
// (12, 14, 'sp4_r_v_b_38')
// (12, 15, 'neigh_op_tnr_7')
// (12, 15, 'sp4_r_v_b_27')
// (12, 16, 'neigh_op_rgt_7')
// (12, 16, 'sp4_r_v_b_14')
// (12, 17, 'neigh_op_bnr_7')
// (12, 17, 'sp4_r_v_b_3')
// (13, 13, 'sp4_v_t_38')
// (13, 14, 'sp4_v_b_38')
// (13, 15, 'local_g2_3')
// (13, 15, 'lutff_3/in_2')
// (13, 15, 'neigh_op_top_7')
// (13, 15, 'sp4_v_b_27')
// (13, 16, 'lutff_7/out')
// (13, 16, 'sp4_v_b_14')
// (13, 17, 'neigh_op_bot_7')
// (13, 17, 'sp4_v_b_3')
// (14, 15, 'neigh_op_tnl_7')
// (14, 16, 'neigh_op_lft_7')
// (14, 17, 'neigh_op_bnl_7')

wire n1802;
// (12, 15, 'neigh_op_tnr_0')
// (12, 16, 'neigh_op_rgt_0')
// (12, 17, 'neigh_op_bnr_0')
// (13, 15, 'local_g0_0')
// (13, 15, 'lutff_3/in_1')
// (13, 15, 'neigh_op_top_0')
// (13, 16, 'lutff_0/out')
// (13, 17, 'neigh_op_bot_0')
// (14, 15, 'neigh_op_tnl_0')
// (14, 16, 'neigh_op_lft_0')
// (14, 17, 'neigh_op_bnl_0')

wire n1803;
// (12, 15, 'neigh_op_tnr_1')
// (12, 16, 'neigh_op_rgt_1')
// (12, 17, 'neigh_op_bnr_1')
// (13, 15, 'local_g0_1')
// (13, 15, 'lutff_4/in_1')
// (13, 15, 'neigh_op_top_1')
// (13, 16, 'lutff_1/out')
// (13, 17, 'neigh_op_bot_1')
// (14, 15, 'neigh_op_tnl_1')
// (14, 16, 'neigh_op_lft_1')
// (14, 17, 'neigh_op_bnl_1')

wire n1804;
// (12, 15, 'neigh_op_tnr_3')
// (12, 16, 'neigh_op_rgt_3')
// (12, 17, 'neigh_op_bnr_3')
// (13, 15, 'local_g1_3')
// (13, 15, 'lutff_4/in_2')
// (13, 15, 'neigh_op_top_3')
// (13, 16, 'lutff_3/out')
// (13, 17, 'neigh_op_bot_3')
// (14, 15, 'neigh_op_tnl_3')
// (14, 16, 'neigh_op_lft_3')
// (14, 17, 'neigh_op_bnl_3')

wire n1805;
// (12, 15, 'neigh_op_tnr_5')
// (12, 16, 'neigh_op_rgt_5')
// (12, 17, 'neigh_op_bnr_5')
// (13, 15, 'local_g0_5')
// (13, 15, 'lutff_5/in_2')
// (13, 15, 'neigh_op_top_5')
// (13, 16, 'lutff_5/out')
// (13, 17, 'neigh_op_bot_5')
// (14, 15, 'neigh_op_tnl_5')
// (14, 16, 'neigh_op_lft_5')
// (14, 17, 'neigh_op_bnl_5')

wire n1806;
// (12, 15, 'neigh_op_tnr_6')
// (12, 16, 'neigh_op_rgt_6')
// (12, 17, 'neigh_op_bnr_6')
// (13, 15, 'local_g1_6')
// (13, 15, 'lutff_2/in_1')
// (13, 15, 'neigh_op_top_6')
// (13, 16, 'lutff_6/out')
// (13, 17, 'neigh_op_bot_6')
// (14, 15, 'neigh_op_tnl_6')
// (14, 16, 'neigh_op_lft_6')
// (14, 17, 'neigh_op_bnl_6')

reg n1807 = 0;
// (12, 15, 'sp4_r_v_b_42')
// (12, 16, 'sp4_r_v_b_31')
// (12, 17, 'local_g3_2')
// (12, 17, 'lutff_0/in_1')
// (12, 17, 'sp4_r_v_b_18')
// (12, 18, 'sp4_r_v_b_7')
// (13, 14, 'sp4_h_r_1')
// (13, 14, 'sp4_v_t_42')
// (13, 15, 'sp4_v_b_42')
// (13, 16, 'sp4_v_b_31')
// (13, 17, 'sp4_v_b_18')
// (13, 18, 'sp4_v_b_7')
// (14, 14, 'sp4_h_r_12')
// (15, 13, 'neigh_op_tnr_2')
// (15, 14, 'neigh_op_rgt_2')
// (15, 14, 'sp4_h_r_25')
// (15, 15, 'neigh_op_bnr_2')
// (16, 11, 'sp4_r_v_b_40')
// (16, 12, 'sp4_r_v_b_29')
// (16, 13, 'neigh_op_top_2')
// (16, 13, 'sp4_r_v_b_16')
// (16, 14, 'local_g1_2')
// (16, 14, 'lutff_1/in_2')
// (16, 14, 'lutff_2/out')
// (16, 14, 'sp4_h_r_36')
// (16, 14, 'sp4_r_v_b_37')
// (16, 14, 'sp4_r_v_b_5')
// (16, 15, 'neigh_op_bot_2')
// (16, 15, 'sp4_r_v_b_24')
// (16, 16, 'local_g2_5')
// (16, 16, 'lutff_3/in_0')
// (16, 16, 'sp4_r_v_b_13')
// (16, 17, 'sp4_r_v_b_0')
// (17, 10, 'sp4_v_t_40')
// (17, 11, 'sp4_v_b_40')
// (17, 12, 'local_g2_5')
// (17, 12, 'lutff_1/in_0')
// (17, 12, 'sp4_v_b_29')
// (17, 13, 'neigh_op_tnl_2')
// (17, 13, 'sp4_v_b_16')
// (17, 13, 'sp4_v_t_37')
// (17, 14, 'neigh_op_lft_2')
// (17, 14, 'sp4_h_l_36')
// (17, 14, 'sp4_v_b_37')
// (17, 14, 'sp4_v_b_5')
// (17, 15, 'neigh_op_bnl_2')
// (17, 15, 'sp4_v_b_24')
// (17, 16, 'sp4_v_b_13')
// (17, 17, 'sp4_v_b_0')

wire n1808;
// (12, 16, 'neigh_op_tnr_2')
// (12, 17, 'neigh_op_rgt_2')
// (12, 18, 'neigh_op_bnr_2')
// (13, 16, 'neigh_op_top_2')
// (13, 17, 'lutff_2/out')
// (13, 18, 'local_g1_2')
// (13, 18, 'lutff_2/in_1')
// (13, 18, 'neigh_op_bot_2')
// (14, 16, 'neigh_op_tnl_2')
// (14, 17, 'neigh_op_lft_2')
// (14, 18, 'neigh_op_bnl_2')

wire n1809;
// (12, 16, 'neigh_op_tnr_4')
// (12, 17, 'neigh_op_rgt_4')
// (12, 18, 'neigh_op_bnr_4')
// (13, 16, 'neigh_op_top_4')
// (13, 17, 'lutff_4/out')
// (13, 18, 'local_g1_4')
// (13, 18, 'lutff_6/in_1')
// (13, 18, 'neigh_op_bot_4')
// (14, 16, 'neigh_op_tnl_4')
// (14, 17, 'neigh_op_lft_4')
// (14, 18, 'neigh_op_bnl_4')

wire n1810;
// (12, 16, 'neigh_op_tnr_6')
// (12, 17, 'neigh_op_rgt_6')
// (12, 18, 'neigh_op_bnr_6')
// (13, 16, 'neigh_op_top_6')
// (13, 17, 'lutff_6/out')
// (13, 18, 'local_g1_6')
// (13, 18, 'lutff_7/in_2')
// (13, 18, 'neigh_op_bot_6')
// (14, 16, 'neigh_op_tnl_6')
// (14, 17, 'neigh_op_lft_6')
// (14, 18, 'neigh_op_bnl_6')

wire n1811;
// (12, 16, 'sp4_h_r_9')
// (13, 16, 'sp4_h_r_20')
// (14, 15, 'neigh_op_tnr_6')
// (14, 16, 'neigh_op_rgt_6')
// (14, 16, 'sp4_h_r_33')
// (14, 17, 'neigh_op_bnr_6')
// (15, 13, 'sp4_r_v_b_38')
// (15, 14, 'sp4_r_v_b_27')
// (15, 15, 'neigh_op_top_6')
// (15, 15, 'sp4_r_v_b_14')
// (15, 16, 'local_g1_3')
// (15, 16, 'lutff_6/out')
// (15, 16, 'lutff_global/cen')
// (15, 16, 'sp4_h_r_44')
// (15, 16, 'sp4_r_v_b_3')
// (15, 17, 'neigh_op_bot_6')
// (16, 12, 'sp4_v_t_38')
// (16, 13, 'sp4_v_b_38')
// (16, 14, 'sp4_v_b_27')
// (16, 15, 'neigh_op_tnl_6')
// (16, 15, 'sp4_v_b_14')
// (16, 16, 'neigh_op_lft_6')
// (16, 16, 'sp4_h_l_44')
// (16, 16, 'sp4_v_b_3')
// (16, 17, 'neigh_op_bnl_6')

reg n1812 = 0;
// (12, 17, 'neigh_op_tnr_2')
// (12, 18, 'neigh_op_rgt_2')
// (12, 18, 'sp4_h_r_9')
// (12, 19, 'neigh_op_bnr_2')
// (13, 15, 'sp4_r_v_b_40')
// (13, 16, 'sp4_r_v_b_29')
// (13, 17, 'local_g1_2')
// (13, 17, 'lutff_3/in_2')
// (13, 17, 'neigh_op_top_2')
// (13, 17, 'sp4_r_v_b_16')
// (13, 18, 'local_g3_2')
// (13, 18, 'lutff_2/in_3')
// (13, 18, 'lutff_2/out')
// (13, 18, 'sp4_h_r_20')
// (13, 18, 'sp4_r_v_b_5')
// (13, 19, 'neigh_op_bot_2')
// (14, 14, 'sp4_v_t_40')
// (14, 15, 'local_g2_0')
// (14, 15, 'lutff_7/in_1')
// (14, 15, 'sp4_v_b_40')
// (14, 16, 'sp4_v_b_29')
// (14, 17, 'neigh_op_tnl_2')
// (14, 17, 'sp4_v_b_16')
// (14, 18, 'neigh_op_lft_2')
// (14, 18, 'sp4_h_r_33')
// (14, 18, 'sp4_v_b_5')
// (14, 19, 'neigh_op_bnl_2')
// (15, 18, 'sp4_h_r_44')
// (16, 18, 'sp4_h_l_44')
// (16, 18, 'sp4_h_r_5')
// (17, 18, 'sp4_h_r_16')
// (18, 18, 'sp4_h_r_29')
// (19, 15, 'sp4_r_v_b_40')
// (19, 16, 'local_g0_5')
// (19, 16, 'ram/WADDR_2')
// (19, 16, 'sp4_r_v_b_29')
// (19, 17, 'sp4_r_v_b_16')
// (19, 18, 'sp4_h_r_40')
// (19, 18, 'sp4_r_v_b_5')
// (20, 14, 'sp4_v_t_40')
// (20, 15, 'sp4_v_b_40')
// (20, 16, 'sp4_v_b_29')
// (20, 17, 'sp4_v_b_16')
// (20, 18, 'sp4_h_l_40')
// (20, 18, 'sp4_v_b_5')

wire n1813;
// (12, 17, 'neigh_op_tnr_4')
// (12, 18, 'local_g3_4')
// (12, 18, 'lutff_7/in_0')
// (12, 18, 'neigh_op_rgt_4')
// (12, 19, 'neigh_op_bnr_4')
// (13, 17, 'neigh_op_top_4')
// (13, 18, 'lutff_4/out')
// (13, 19, 'neigh_op_bot_4')
// (14, 17, 'neigh_op_tnl_4')
// (14, 18, 'neigh_op_lft_4')
// (14, 19, 'local_g3_4')
// (14, 19, 'lutff_6/in_1')
// (14, 19, 'neigh_op_bnl_4')

wire n1814;
// (12, 17, 'neigh_op_tnr_5')
// (12, 18, 'neigh_op_rgt_5')
// (12, 19, 'neigh_op_bnr_5')
// (13, 17, 'neigh_op_top_5')
// (13, 18, 'local_g3_5')
// (13, 18, 'lutff_4/in_2')
// (13, 18, 'lutff_5/out')
// (13, 19, 'neigh_op_bot_5')
// (14, 17, 'neigh_op_tnl_5')
// (14, 18, 'neigh_op_lft_5')
// (14, 19, 'neigh_op_bnl_5')

wire n1815;
// (12, 17, 'sp4_r_v_b_43')
// (12, 18, 'sp4_r_v_b_30')
// (12, 19, 'local_g3_3')
// (12, 19, 'lutff_global/cen')
// (12, 19, 'sp4_r_v_b_19')
// (12, 20, 'sp4_r_v_b_6')
// (13, 16, 'sp4_v_t_43')
// (13, 17, 'sp4_v_b_43')
// (13, 18, 'sp4_v_b_30')
// (13, 19, 'local_g1_3')
// (13, 19, 'lutff_global/cen')
// (13, 19, 'sp4_v_b_19')
// (13, 20, 'sp4_h_r_6')
// (13, 20, 'sp4_v_b_6')
// (14, 18, 'sp4_r_v_b_38')
// (14, 19, 'neigh_op_tnr_7')
// (14, 19, 'sp4_r_v_b_27')
// (14, 20, 'neigh_op_rgt_7')
// (14, 20, 'sp4_h_r_19')
// (14, 20, 'sp4_h_r_3')
// (14, 20, 'sp4_h_r_6')
// (14, 20, 'sp4_r_v_b_14')
// (14, 21, 'neigh_op_bnr_7')
// (14, 21, 'sp4_r_v_b_3')
// (15, 17, 'local_g1_3')
// (15, 17, 'lutff_global/cen')
// (15, 17, 'sp4_h_r_3')
// (15, 17, 'sp4_v_t_38')
// (15, 18, 'sp4_v_b_38')
// (15, 19, 'neigh_op_top_7')
// (15, 19, 'sp4_v_b_27')
// (15, 20, 'local_g1_3')
// (15, 20, 'lutff_7/out')
// (15, 20, 'lutff_global/cen')
// (15, 20, 'sp4_h_r_14')
// (15, 20, 'sp4_h_r_19')
// (15, 20, 'sp4_h_r_30')
// (15, 20, 'sp4_v_b_14')
// (15, 21, 'neigh_op_bot_7')
// (15, 21, 'sp4_v_b_3')
// (16, 17, 'sp4_h_r_14')
// (16, 19, 'neigh_op_tnl_7')
// (16, 20, 'neigh_op_lft_7')
// (16, 20, 'sp4_h_r_27')
// (16, 20, 'sp4_h_r_30')
// (16, 20, 'sp4_h_r_43')
// (16, 21, 'neigh_op_bnl_7')
// (17, 17, 'sp4_h_r_27')
// (17, 20, 'sp4_h_l_43')
// (17, 20, 'sp4_h_r_38')
// (17, 20, 'sp4_h_r_43')
// (18, 17, 'sp4_h_r_38')
// (18, 20, 'sp4_h_l_38')
// (18, 20, 'sp4_h_l_43')
// (18, 20, 'sp4_h_r_3')
// (19, 17, 'sp4_h_l_38')
// (19, 20, 'sp4_h_r_14')
// (20, 20, 'sp4_h_r_27')
// (21, 20, 'sp4_h_r_38')
// (22, 20, 'sp4_h_l_38')

wire n1816;
// (12, 18, 'neigh_op_tnr_1')
// (12, 19, 'neigh_op_rgt_1')
// (12, 20, 'neigh_op_bnr_1')
// (13, 17, 'sp4_r_v_b_43')
// (13, 18, 'neigh_op_top_1')
// (13, 18, 'sp4_r_v_b_30')
// (13, 19, 'lutff_1/out')
// (13, 19, 'sp4_r_v_b_19')
// (13, 20, 'neigh_op_bot_1')
// (13, 20, 'sp4_r_v_b_6')
// (14, 16, 'sp4_v_t_43')
// (14, 17, 'sp4_v_b_43')
// (14, 18, 'neigh_op_tnl_1')
// (14, 18, 'sp4_v_b_30')
// (14, 19, 'neigh_op_lft_1')
// (14, 19, 'sp4_v_b_19')
// (14, 20, 'neigh_op_bnl_1')
// (14, 20, 'sp4_h_r_0')
// (14, 20, 'sp4_v_b_6')
// (15, 20, 'local_g1_5')
// (15, 20, 'lutff_2/in_2')
// (15, 20, 'sp4_h_r_13')
// (16, 20, 'sp4_h_r_24')
// (17, 20, 'sp4_h_r_37')
// (18, 20, 'sp4_h_l_37')

wire n1817;
// (12, 18, 'neigh_op_tnr_2')
// (12, 19, 'local_g3_2')
// (12, 19, 'lutff_1/in_0')
// (12, 19, 'neigh_op_rgt_2')
// (12, 20, 'neigh_op_bnr_2')
// (13, 18, 'neigh_op_top_2')
// (13, 19, 'lutff_2/out')
// (13, 20, 'neigh_op_bot_2')
// (14, 18, 'neigh_op_tnl_2')
// (14, 19, 'neigh_op_lft_2')
// (14, 20, 'neigh_op_bnl_2')

wire n1818;
// (12, 18, 'neigh_op_tnr_3')
// (12, 19, 'neigh_op_rgt_3')
// (12, 20, 'neigh_op_bnr_3')
// (13, 17, 'sp4_r_v_b_47')
// (13, 18, 'neigh_op_top_3')
// (13, 18, 'sp4_r_v_b_34')
// (13, 19, 'lutff_3/out')
// (13, 19, 'sp4_r_v_b_23')
// (13, 20, 'neigh_op_bot_3')
// (13, 20, 'sp4_r_v_b_10')
// (14, 16, 'sp4_v_t_47')
// (14, 17, 'sp4_v_b_47')
// (14, 18, 'neigh_op_tnl_3')
// (14, 18, 'sp4_v_b_34')
// (14, 19, 'neigh_op_lft_3')
// (14, 19, 'sp4_v_b_23')
// (14, 20, 'neigh_op_bnl_3')
// (14, 20, 'sp4_h_r_10')
// (14, 20, 'sp4_v_b_10')
// (15, 20, 'local_g0_7')
// (15, 20, 'lutff_6/in_3')
// (15, 20, 'sp4_h_r_23')
// (16, 20, 'sp4_h_r_34')
// (17, 20, 'sp4_h_r_47')
// (18, 20, 'sp4_h_l_47')

wire n1819;
// (12, 18, 'neigh_op_tnr_4')
// (12, 19, 'neigh_op_rgt_4')
// (12, 20, 'neigh_op_bnr_4')
// (13, 18, 'neigh_op_top_4')
// (13, 19, 'local_g3_4')
// (13, 19, 'lutff_4/out')
// (13, 19, 'lutff_7/in_0')
// (13, 20, 'neigh_op_bot_4')
// (14, 18, 'neigh_op_tnl_4')
// (14, 19, 'neigh_op_lft_4')
// (14, 20, 'neigh_op_bnl_4')

wire n1820;
// (12, 18, 'neigh_op_tnr_5')
// (12, 19, 'local_g2_5')
// (12, 19, 'lutff_7/in_2')
// (12, 19, 'neigh_op_rgt_5')
// (12, 20, 'neigh_op_bnr_5')
// (13, 18, 'neigh_op_top_5')
// (13, 19, 'lutff_5/out')
// (13, 20, 'neigh_op_bot_5')
// (14, 18, 'neigh_op_tnl_5')
// (14, 19, 'neigh_op_lft_5')
// (14, 20, 'neigh_op_bnl_5')

wire n1821;
// (12, 18, 'neigh_op_tnr_6')
// (12, 19, 'local_g3_6')
// (12, 19, 'lutff_3/in_0')
// (12, 19, 'neigh_op_rgt_6')
// (12, 20, 'neigh_op_bnr_6')
// (13, 18, 'neigh_op_top_6')
// (13, 19, 'lutff_6/out')
// (13, 20, 'neigh_op_bot_6')
// (14, 18, 'neigh_op_tnl_6')
// (14, 19, 'neigh_op_lft_6')
// (14, 20, 'neigh_op_bnl_6')

reg n1822 = 0;
// (12, 18, 'sp4_h_r_4')
// (12, 18, 'sp4_r_v_b_39')
// (12, 19, 'sp4_h_r_9')
// (12, 19, 'sp4_r_v_b_26')
// (12, 20, 'sp4_r_v_b_15')
// (12, 21, 'sp4_r_v_b_2')
// (13, 17, 'sp4_h_r_8')
// (13, 17, 'sp4_v_t_39')
// (13, 18, 'local_g0_1')
// (13, 18, 'lutff_4/in_1')
// (13, 18, 'sp4_h_r_17')
// (13, 18, 'sp4_v_b_39')
// (13, 19, 'local_g1_4')
// (13, 19, 'local_g2_2')
// (13, 19, 'lutff_0/in_1')
// (13, 19, 'lutff_1/in_3')
// (13, 19, 'sp4_h_r_20')
// (13, 19, 'sp4_v_b_26')
// (13, 20, 'local_g0_7')
// (13, 20, 'lutff_0/in_1')
// (13, 20, 'sp4_v_b_15')
// (13, 21, 'sp4_v_b_2')
// (14, 1, 'sp4_r_v_b_34')
// (14, 2, 'local_g3_7')
// (14, 2, 'lutff_7/in_1')
// (14, 2, 'sp4_r_v_b_23')
// (14, 3, 'sp4_r_v_b_10')
// (14, 4, 'sp4_r_v_b_47')
// (14, 5, 'sp4_r_v_b_34')
// (14, 6, 'sp4_r_v_b_23')
// (14, 7, 'sp4_r_v_b_10')
// (14, 16, 'neigh_op_tnr_0')
// (14, 17, 'neigh_op_rgt_0')
// (14, 17, 'sp4_h_r_21')
// (14, 18, 'neigh_op_bnr_0')
// (14, 18, 'sp4_h_r_28')
// (14, 19, 'sp4_h_r_33')
// (15, 0, 'span4_vert_34')
// (15, 1, 'sp4_v_b_34')
// (15, 2, 'sp4_v_b_23')
// (15, 3, 'sp4_v_b_10')
// (15, 3, 'sp4_v_t_47')
// (15, 4, 'sp4_v_b_47')
// (15, 5, 'sp12_v_t_23')
// (15, 5, 'sp4_v_b_34')
// (15, 6, 'sp12_v_b_23')
// (15, 6, 'sp4_v_b_23')
// (15, 7, 'sp12_v_b_20')
// (15, 7, 'sp4_v_b_10')
// (15, 8, 'sp12_v_b_19')
// (15, 9, 'sp12_v_b_16')
// (15, 10, 'sp12_v_b_15')
// (15, 11, 'sp12_v_b_12')
// (15, 12, 'sp12_v_b_11')
// (15, 13, 'sp12_v_b_8')
// (15, 14, 'sp12_v_b_7')
// (15, 14, 'sp4_r_v_b_36')
// (15, 15, 'sp12_v_b_4')
// (15, 15, 'sp4_r_v_b_25')
// (15, 15, 'sp4_r_v_b_41')
// (15, 16, 'neigh_op_top_0')
// (15, 16, 'sp12_v_b_3')
// (15, 16, 'sp4_r_v_b_12')
// (15, 16, 'sp4_r_v_b_28')
// (15, 16, 'sp4_r_v_b_44')
// (15, 17, 'local_g1_0')
// (15, 17, 'lutff_0/in_3')
// (15, 17, 'lutff_0/out')
// (15, 17, 'sp12_v_b_0')
// (15, 17, 'sp4_h_r_32')
// (15, 17, 'sp4_r_v_b_1')
// (15, 17, 'sp4_r_v_b_17')
// (15, 17, 'sp4_r_v_b_33')
// (15, 18, 'neigh_op_bot_0')
// (15, 18, 'sp4_h_r_41')
// (15, 18, 'sp4_r_v_b_20')
// (15, 18, 'sp4_r_v_b_36')
// (15, 18, 'sp4_r_v_b_4')
// (15, 19, 'sp4_h_r_44')
// (15, 19, 'sp4_r_v_b_25')
// (15, 19, 'sp4_r_v_b_9')
// (15, 20, 'local_g2_4')
// (15, 20, 'lutff_3/in_1')
// (15, 20, 'sp4_r_v_b_12')
// (15, 21, 'sp4_r_v_b_1')
// (16, 13, 'sp4_v_t_36')
// (16, 14, 'sp4_v_b_36')
// (16, 14, 'sp4_v_t_41')
// (16, 15, 'sp4_v_b_25')
// (16, 15, 'sp4_v_b_41')
// (16, 15, 'sp4_v_t_44')
// (16, 16, 'neigh_op_tnl_0')
// (16, 16, 'sp4_v_b_12')
// (16, 16, 'sp4_v_b_28')
// (16, 16, 'sp4_v_b_44')
// (16, 17, 'neigh_op_lft_0')
// (16, 17, 'sp4_h_r_45')
// (16, 17, 'sp4_v_b_1')
// (16, 17, 'sp4_v_b_17')
// (16, 17, 'sp4_v_b_33')
// (16, 17, 'sp4_v_t_36')
// (16, 18, 'neigh_op_bnl_0')
// (16, 18, 'sp4_h_l_41')
// (16, 18, 'sp4_v_b_20')
// (16, 18, 'sp4_v_b_36')
// (16, 18, 'sp4_v_b_4')
// (16, 19, 'sp4_h_l_44')
// (16, 19, 'sp4_v_b_25')
// (16, 19, 'sp4_v_b_9')
// (16, 20, 'sp4_v_b_12')
// (16, 21, 'sp4_v_b_1')
// (17, 17, 'sp4_h_l_45')

wire n1823;
// (12, 18, 'sp4_h_r_5')
// (13, 18, 'sp4_h_r_16')
// (14, 18, 'local_g3_5')
// (14, 18, 'lutff_0/in_0')
// (14, 18, 'lutff_1/in_1')
// (14, 18, 'lutff_3/in_1')
// (14, 18, 'sp4_h_r_29')
// (15, 15, 'neigh_op_tnr_4')
// (15, 15, 'sp4_r_v_b_37')
// (15, 16, 'neigh_op_rgt_4')
// (15, 16, 'sp4_r_v_b_24')
// (15, 16, 'sp4_r_v_b_40')
// (15, 17, 'neigh_op_bnr_4')
// (15, 17, 'sp4_r_v_b_13')
// (15, 17, 'sp4_r_v_b_29')
// (15, 18, 'sp4_h_r_40')
// (15, 18, 'sp4_r_v_b_0')
// (15, 18, 'sp4_r_v_b_16')
// (15, 19, 'sp4_r_v_b_5')
// (16, 14, 'sp4_v_t_37')
// (16, 15, 'neigh_op_top_4')
// (16, 15, 'sp4_v_b_37')
// (16, 15, 'sp4_v_t_40')
// (16, 16, 'lutff_4/out')
// (16, 16, 'sp4_v_b_24')
// (16, 16, 'sp4_v_b_40')
// (16, 17, 'local_g1_4')
// (16, 17, 'lutff_5/in_2')
// (16, 17, 'neigh_op_bot_4')
// (16, 17, 'sp4_v_b_13')
// (16, 17, 'sp4_v_b_29')
// (16, 18, 'local_g1_0')
// (16, 18, 'lutff_1/in_0')
// (16, 18, 'sp4_h_l_40')
// (16, 18, 'sp4_v_b_0')
// (16, 18, 'sp4_v_b_16')
// (16, 19, 'local_g0_5')
// (16, 19, 'lutff_4/in_1')
// (16, 19, 'lutff_6/in_1')
// (16, 19, 'lutff_7/in_0')
// (16, 19, 'sp4_v_b_5')
// (17, 15, 'neigh_op_tnl_4')
// (17, 16, 'neigh_op_lft_4')
// (17, 17, 'neigh_op_bnl_4')

wire n1824;
// (12, 19, 'local_g2_2')
// (12, 19, 'lutff_1/in_1')
// (12, 19, 'neigh_op_tnr_2')
// (12, 20, 'neigh_op_rgt_2')
// (12, 21, 'neigh_op_bnr_2')
// (13, 19, 'neigh_op_top_2')
// (13, 20, 'lutff_2/out')
// (13, 21, 'neigh_op_bot_2')
// (14, 19, 'neigh_op_tnl_2')
// (14, 20, 'neigh_op_lft_2')
// (14, 21, 'neigh_op_bnl_2')

wire n1825;
// (12, 19, 'local_g2_6')
// (12, 19, 'lutff_3/in_3')
// (12, 19, 'neigh_op_tnr_6')
// (12, 20, 'neigh_op_rgt_6')
// (12, 21, 'neigh_op_bnr_6')
// (13, 19, 'neigh_op_top_6')
// (13, 20, 'lutff_6/out')
// (13, 21, 'neigh_op_bot_6')
// (14, 19, 'neigh_op_tnl_6')
// (14, 20, 'neigh_op_lft_6')
// (14, 21, 'neigh_op_bnl_6')

wire n1826;
// (12, 19, 'local_g3_5')
// (12, 19, 'lutff_7/in_3')
// (12, 19, 'neigh_op_tnr_5')
// (12, 20, 'neigh_op_rgt_5')
// (12, 21, 'neigh_op_bnr_5')
// (13, 19, 'neigh_op_top_5')
// (13, 20, 'lutff_5/out')
// (13, 21, 'neigh_op_bot_5')
// (14, 19, 'neigh_op_tnl_5')
// (14, 20, 'neigh_op_lft_5')
// (14, 21, 'neigh_op_bnl_5')

wire n1827;
// (12, 19, 'neigh_op_tnr_3')
// (12, 20, 'neigh_op_rgt_3')
// (12, 20, 'sp4_h_r_11')
// (12, 21, 'neigh_op_bnr_3')
// (13, 19, 'neigh_op_top_3')
// (13, 20, 'lutff_3/out')
// (13, 20, 'sp4_h_r_22')
// (13, 21, 'neigh_op_bot_3')
// (14, 19, 'neigh_op_tnl_3')
// (14, 20, 'neigh_op_lft_3')
// (14, 20, 'sp4_h_r_35')
// (14, 21, 'neigh_op_bnl_3')
// (15, 20, 'local_g2_6')
// (15, 20, 'lutff_6/in_2')
// (15, 20, 'sp4_h_r_46')
// (16, 20, 'sp4_h_l_46')

wire n1828;
// (12, 19, 'neigh_op_tnr_4')
// (12, 20, 'neigh_op_rgt_4')
// (12, 21, 'neigh_op_bnr_4')
// (13, 19, 'local_g0_4')
// (13, 19, 'lutff_7/in_3')
// (13, 19, 'neigh_op_top_4')
// (13, 20, 'lutff_4/out')
// (13, 21, 'neigh_op_bot_4')
// (14, 19, 'neigh_op_tnl_4')
// (14, 20, 'neigh_op_lft_4')
// (14, 21, 'neigh_op_bnl_4')

reg n1829 = 0;
// (12, 19, 'neigh_op_tnr_7')
// (12, 20, 'neigh_op_rgt_7')
// (12, 21, 'neigh_op_bnr_7')
// (13, 19, 'neigh_op_top_7')
// (13, 19, 'sp4_r_v_b_42')
// (13, 20, 'lutff_7/out')
// (13, 20, 'sp4_r_v_b_31')
// (13, 21, 'neigh_op_bot_7')
// (13, 21, 'sp4_r_v_b_18')
// (13, 22, 'sp4_r_v_b_7')
// (14, 18, 'sp4_h_r_7')
// (14, 18, 'sp4_v_t_42')
// (14, 19, 'neigh_op_tnl_7')
// (14, 19, 'sp4_v_b_42')
// (14, 20, 'neigh_op_lft_7')
// (14, 20, 'sp4_v_b_31')
// (14, 21, 'neigh_op_bnl_7')
// (14, 21, 'sp4_v_b_18')
// (14, 22, 'sp4_v_b_7')
// (15, 18, 'sp4_h_r_18')
// (16, 18, 'sp4_h_r_31')
// (17, 18, 'local_g3_2')
// (17, 18, 'lutff_6/in_1')
// (17, 18, 'sp4_h_r_42')
// (18, 18, 'sp4_h_l_42')

wire n1830;
// (12, 20, 'neigh_op_tnr_0')
// (12, 21, 'neigh_op_rgt_0')
// (12, 22, 'neigh_op_bnr_0')
// (13, 20, 'neigh_op_top_0')
// (13, 20, 'sp4_r_v_b_44')
// (13, 21, 'local_g0_2')
// (13, 21, 'lutff_0/out')
// (13, 21, 'lutff_global/cen')
// (13, 21, 'sp4_r_v_b_33')
// (13, 22, 'neigh_op_bot_0')
// (13, 22, 'sp4_r_v_b_20')
// (13, 23, 'sp4_r_v_b_9')
// (14, 19, 'sp4_v_t_44')
// (14, 20, 'neigh_op_tnl_0')
// (14, 20, 'sp4_v_b_44')
// (14, 21, 'neigh_op_lft_0')
// (14, 21, 'sp4_v_b_33')
// (14, 22, 'neigh_op_bnl_0')
// (14, 22, 'sp4_v_b_20')
// (14, 23, 'sp4_v_b_9')

reg n1831 = 0;
// (12, 20, 'neigh_op_tnr_1')
// (12, 21, 'local_g3_1')
// (12, 21, 'lutff_1/in_1')
// (12, 21, 'neigh_op_rgt_1')
// (12, 22, 'neigh_op_bnr_1')
// (13, 20, 'neigh_op_top_1')
// (13, 21, 'lutff_1/out')
// (13, 22, 'neigh_op_bot_1')
// (14, 20, 'local_g2_1')
// (14, 20, 'lutff_4/in_1')
// (14, 20, 'neigh_op_tnl_1')
// (14, 21, 'neigh_op_lft_1')
// (14, 22, 'neigh_op_bnl_1')

reg n1832 = 0;
// (12, 20, 'neigh_op_tnr_2')
// (12, 21, 'local_g2_2')
// (12, 21, 'lutff_3/in_1')
// (12, 21, 'neigh_op_rgt_2')
// (12, 22, 'neigh_op_bnr_2')
// (13, 20, 'neigh_op_top_2')
// (13, 21, 'lutff_2/out')
// (13, 22, 'neigh_op_bot_2')
// (14, 20, 'local_g3_2')
// (14, 20, 'lutff_3/in_2')
// (14, 20, 'neigh_op_tnl_2')
// (14, 21, 'neigh_op_lft_2')
// (14, 22, 'neigh_op_bnl_2')

reg n1833 = 0;
// (12, 20, 'neigh_op_tnr_3')
// (12, 21, 'local_g3_3')
// (12, 21, 'lutff_0/in_2')
// (12, 21, 'lutff_1/in_3')
// (12, 21, 'neigh_op_rgt_3')
// (12, 22, 'neigh_op_bnr_3')
// (13, 20, 'neigh_op_top_3')
// (13, 21, 'local_g2_3')
// (13, 21, 'lutff_3/in_0')
// (13, 21, 'lutff_3/out')
// (13, 22, 'neigh_op_bot_3')
// (14, 20, 'local_g3_3')
// (14, 20, 'lutff_2/in_0')
// (14, 20, 'neigh_op_tnl_3')
// (14, 21, 'neigh_op_lft_3')
// (14, 22, 'neigh_op_bnl_3')

reg n1834 = 0;
// (12, 20, 'neigh_op_tnr_6')
// (12, 21, 'local_g3_6')
// (12, 21, 'lutff_2/in_1')
// (12, 21, 'neigh_op_rgt_6')
// (12, 22, 'neigh_op_bnr_6')
// (13, 20, 'neigh_op_top_6')
// (13, 21, 'lutff_6/out')
// (13, 22, 'neigh_op_bot_6')
// (14, 20, 'local_g2_6')
// (14, 20, 'lutff_0/in_0')
// (14, 20, 'neigh_op_tnl_6')
// (14, 21, 'neigh_op_lft_6')
// (14, 22, 'neigh_op_bnl_6')

wire n1835;
// (12, 20, 'neigh_op_tnr_7')
// (12, 21, 'neigh_op_rgt_7')
// (12, 21, 'sp4_r_v_b_46')
// (12, 22, 'local_g1_7')
// (12, 22, 'lutff_7/in_3')
// (12, 22, 'neigh_op_bnr_7')
// (12, 22, 'sp4_r_v_b_35')
// (12, 23, 'local_g3_6')
// (12, 23, 'lutff_4/in_1')
// (12, 23, 'sp4_r_v_b_22')
// (12, 24, 'sp4_r_v_b_11')
// (13, 20, 'neigh_op_top_7')
// (13, 20, 'sp4_v_t_46')
// (13, 21, 'lutff_7/out')
// (13, 21, 'sp4_r_v_b_47')
// (13, 21, 'sp4_v_b_46')
// (13, 22, 'local_g1_7')
// (13, 22, 'lutff_0/in_0')
// (13, 22, 'lutff_2/in_0')
// (13, 22, 'lutff_3/in_1')
// (13, 22, 'lutff_4/in_2')
// (13, 22, 'lutff_6/in_2')
// (13, 22, 'neigh_op_bot_7')
// (13, 22, 'sp4_r_v_b_34')
// (13, 22, 'sp4_v_b_35')
// (13, 23, 'local_g3_7')
// (13, 23, 'lutff_7/in_1')
// (13, 23, 'sp4_r_v_b_23')
// (13, 23, 'sp4_v_b_22')
// (13, 24, 'sp4_r_v_b_10')
// (13, 24, 'sp4_v_b_11')
// (14, 20, 'neigh_op_tnl_7')
// (14, 20, 'sp4_v_t_47')
// (14, 21, 'neigh_op_lft_7')
// (14, 21, 'sp4_v_b_47')
// (14, 22, 'neigh_op_bnl_7')
// (14, 22, 'sp4_v_b_34')
// (14, 23, 'sp4_v_b_23')
// (14, 24, 'sp4_v_b_10')

reg n1836 = 0;
// (12, 20, 'sp4_h_r_1')
// (13, 17, 'sp4_r_v_b_39')
// (13, 17, 'sp4_r_v_b_44')
// (13, 18, 'local_g0_2')
// (13, 18, 'lutff_4/in_0')
// (13, 18, 'sp4_r_v_b_26')
// (13, 18, 'sp4_r_v_b_33')
// (13, 19, 'local_g2_7')
// (13, 19, 'lutff_1/in_2')
// (13, 19, 'sp4_r_v_b_15')
// (13, 19, 'sp4_r_v_b_20')
// (13, 20, 'local_g0_4')
// (13, 20, 'lutff_1/in_1')
// (13, 20, 'sp4_h_r_12')
// (13, 20, 'sp4_r_v_b_2')
// (13, 20, 'sp4_r_v_b_9')
// (14, 16, 'sp4_v_t_39')
// (14, 16, 'sp4_v_t_44')
// (14, 17, 'sp4_v_b_39')
// (14, 17, 'sp4_v_b_44')
// (14, 18, 'sp4_v_b_26')
// (14, 18, 'sp4_v_b_33')
// (14, 19, 'neigh_op_tnr_2')
// (14, 19, 'sp4_v_b_15')
// (14, 19, 'sp4_v_b_20')
// (14, 20, 'neigh_op_rgt_2')
// (14, 20, 'sp4_h_r_25')
// (14, 20, 'sp4_h_r_9')
// (14, 20, 'sp4_v_b_2')
// (14, 20, 'sp4_v_b_9')
// (14, 21, 'neigh_op_bnr_2')
// (15, 0, 'span12_vert_19')
// (15, 1, 'sp12_v_b_19')
// (15, 2, 'sp12_v_b_16')
// (15, 3, 'sp12_v_b_15')
// (15, 4, 'local_g3_4')
// (15, 4, 'lutff_5/in_2')
// (15, 4, 'sp12_v_b_12')
// (15, 5, 'sp12_v_b_11')
// (15, 6, 'sp12_v_b_8')
// (15, 7, 'sp12_v_b_7')
// (15, 8, 'sp12_v_b_4')
// (15, 9, 'sp12_v_b_3')
// (15, 10, 'sp12_v_b_0')
// (15, 10, 'sp12_v_t_23')
// (15, 11, 'sp12_v_b_23')
// (15, 12, 'sp12_v_b_20')
// (15, 13, 'sp12_v_b_19')
// (15, 14, 'sp12_v_b_16')
// (15, 15, 'sp12_v_b_15')
// (15, 16, 'sp12_v_b_12')
// (15, 17, 'sp12_v_b_11')
// (15, 18, 'sp12_v_b_8')
// (15, 19, 'neigh_op_top_2')
// (15, 19, 'sp12_v_b_7')
// (15, 20, 'local_g3_2')
// (15, 20, 'lutff_2/out')
// (15, 20, 'lutff_3/in_0')
// (15, 20, 'sp12_v_b_4')
// (15, 20, 'sp4_h_r_20')
// (15, 20, 'sp4_h_r_36')
// (15, 21, 'neigh_op_bot_2')
// (15, 21, 'sp12_v_b_3')
// (15, 22, 'sp12_v_b_0')
// (16, 19, 'neigh_op_tnl_2')
// (16, 20, 'neigh_op_lft_2')
// (16, 20, 'sp4_h_l_36')
// (16, 20, 'sp4_h_r_33')
// (16, 21, 'neigh_op_bnl_2')
// (17, 20, 'sp4_h_r_44')
// (18, 20, 'sp4_h_l_44')

wire n1837;
// (12, 20, 'sp4_h_r_6')
// (13, 20, 'sp4_h_r_19')
// (14, 20, 'sp4_h_r_30')
// (15, 20, 'sp4_h_r_43')
// (16, 20, 'sp4_h_l_43')
// (16, 20, 'sp4_h_r_2')
// (16, 20, 'sp4_h_r_6')
// (17, 19, 'neigh_op_tnr_7')
// (17, 20, 'neigh_op_rgt_7')
// (17, 20, 'sp4_h_r_15')
// (17, 20, 'sp4_h_r_19')
// (17, 21, 'neigh_op_bnr_7')
// (18, 19, 'neigh_op_top_7')
// (18, 20, 'local_g2_2')
// (18, 20, 'lutff_7/out')
// (18, 20, 'lutff_global/cen')
// (18, 20, 'sp4_h_r_26')
// (18, 20, 'sp4_h_r_30')
// (18, 21, 'neigh_op_bot_7')
// (19, 19, 'neigh_op_tnl_7')
// (19, 20, 'neigh_op_lft_7')
// (19, 20, 'sp4_h_r_39')
// (19, 20, 'sp4_h_r_43')
// (19, 21, 'neigh_op_bnl_7')
// (20, 20, 'sp4_h_l_39')
// (20, 20, 'sp4_h_l_43')

wire n1838;
// (12, 20, 'sp4_h_r_7')
// (13, 20, 'local_g0_2')
// (13, 20, 'lutff_global/cen')
// (13, 20, 'sp4_h_r_1')
// (13, 20, 'sp4_h_r_18')
// (13, 20, 'sp4_h_r_7')
// (14, 20, 'local_g0_2')
// (14, 20, 'lutff_global/cen')
// (14, 20, 'sp4_h_r_12')
// (14, 20, 'sp4_h_r_18')
// (14, 20, 'sp4_h_r_31')
// (15, 19, 'neigh_op_tnr_2')
// (15, 20, 'neigh_op_rgt_2')
// (15, 20, 'sp4_h_r_25')
// (15, 20, 'sp4_h_r_31')
// (15, 20, 'sp4_h_r_42')
// (15, 21, 'neigh_op_bnr_2')
// (16, 19, 'neigh_op_top_2')
// (16, 20, 'lutff_2/out')
// (16, 20, 'sp4_h_l_42')
// (16, 20, 'sp4_h_r_36')
// (16, 20, 'sp4_h_r_4')
// (16, 20, 'sp4_h_r_42')
// (16, 21, 'neigh_op_bot_2')
// (17, 19, 'neigh_op_tnl_2')
// (17, 20, 'neigh_op_lft_2')
// (17, 20, 'sp4_h_l_36')
// (17, 20, 'sp4_h_l_42')
// (17, 20, 'sp4_h_r_17')
// (17, 20, 'sp4_h_r_4')
// (17, 21, 'neigh_op_bnl_2')
// (18, 20, 'sp4_h_r_17')
// (18, 20, 'sp4_h_r_28')
// (19, 20, 'sp4_h_r_28')
// (19, 20, 'sp4_h_r_41')
// (20, 20, 'sp4_h_l_41')
// (20, 20, 'sp4_h_r_41')
// (21, 20, 'sp4_h_l_41')

wire n1839;
// (12, 21, 'lutff_1/cout')
// (12, 21, 'lutff_2/in_3')

wire n1840;
// (12, 21, 'lutff_2/cout')
// (12, 21, 'lutff_3/in_3')

wire n1841;
// (12, 21, 'neigh_op_tnr_0')
// (12, 22, 'neigh_op_rgt_0')
// (12, 23, 'neigh_op_bnr_0')
// (13, 21, 'neigh_op_top_0')
// (13, 22, 'local_g2_0')
// (13, 22, 'lutff_0/out')
// (13, 22, 'lutff_5/in_1')
// (13, 23, 'neigh_op_bot_0')
// (14, 21, 'neigh_op_tnl_0')
// (14, 22, 'neigh_op_lft_0')
// (14, 23, 'neigh_op_bnl_0')

wire n1842;
// (12, 21, 'neigh_op_tnr_1')
// (12, 22, 'neigh_op_rgt_1')
// (12, 23, 'neigh_op_bnr_1')
// (13, 21, 'neigh_op_top_1')
// (13, 22, 'local_g2_1')
// (13, 22, 'lutff_0/in_3')
// (13, 22, 'lutff_1/out')
// (13, 22, 'lutff_7/in_0')
// (13, 23, 'local_g0_1')
// (13, 23, 'local_g1_1')
// (13, 23, 'lutff_1/in_0')
// (13, 23, 'lutff_2/in_0')
// (13, 23, 'lutff_3/in_0')
// (13, 23, 'lutff_4/in_0')
// (13, 23, 'lutff_5/in_0')
// (13, 23, 'lutff_6/in_0')
// (13, 23, 'neigh_op_bot_1')
// (14, 21, 'neigh_op_tnl_1')
// (14, 22, 'neigh_op_lft_1')
// (14, 23, 'neigh_op_bnl_1')

reg n1843 = 0;
// (12, 21, 'neigh_op_tnr_2')
// (12, 22, 'local_g2_2')
// (12, 22, 'lutff_2/in_2')
// (12, 22, 'neigh_op_rgt_2')
// (12, 23, 'neigh_op_bnr_2')
// (13, 21, 'neigh_op_top_2')
// (13, 22, 'lutff_2/out')
// (13, 23, 'neigh_op_bot_2')
// (14, 21, 'neigh_op_tnl_2')
// (14, 22, 'local_g1_2')
// (14, 22, 'lutff_1/in_2')
// (14, 22, 'neigh_op_lft_2')
// (14, 23, 'local_g3_2')
// (14, 23, 'lutff_2/in_1')
// (14, 23, 'neigh_op_bnl_2')

wire n1844;
// (12, 21, 'neigh_op_tnr_3')
// (12, 22, 'neigh_op_rgt_3')
// (12, 23, 'neigh_op_bnr_3')
// (13, 21, 'neigh_op_top_3')
// (13, 22, 'local_g3_3')
// (13, 22, 'lutff_3/out')
// (13, 22, 'lutff_7/in_3')
// (13, 23, 'neigh_op_bot_3')
// (14, 21, 'neigh_op_tnl_3')
// (14, 22, 'neigh_op_lft_3')
// (14, 23, 'neigh_op_bnl_3')

reg n1845 = 0;
// (12, 21, 'neigh_op_tnr_4')
// (12, 22, 'local_g3_4')
// (12, 22, 'lutff_3/in_2')
// (12, 22, 'neigh_op_rgt_4')
// (12, 23, 'neigh_op_bnr_4')
// (13, 21, 'neigh_op_top_4')
// (13, 22, 'lutff_4/out')
// (13, 23, 'neigh_op_bot_4')
// (14, 21, 'neigh_op_tnl_4')
// (14, 22, 'local_g1_4')
// (14, 22, 'lutff_1/in_0')
// (14, 22, 'neigh_op_lft_4')
// (14, 23, 'local_g2_4')
// (14, 23, 'lutff_3/in_1')
// (14, 23, 'neigh_op_bnl_4')

reg n1846 = 0;
// (12, 21, 'neigh_op_tnr_5')
// (12, 22, 'local_g2_5')
// (12, 22, 'local_g3_5')
// (12, 22, 'lutff_0/in_1')
// (12, 22, 'lutff_1/in_3')
// (12, 22, 'neigh_op_rgt_5')
// (12, 23, 'neigh_op_bnr_5')
// (13, 21, 'neigh_op_top_5')
// (13, 22, 'local_g3_5')
// (13, 22, 'lutff_0/in_2')
// (13, 22, 'lutff_5/out')
// (13, 23, 'neigh_op_bot_5')
// (14, 21, 'neigh_op_tnl_5')
// (14, 22, 'local_g1_5')
// (14, 22, 'lutff_5/in_3')
// (14, 22, 'lutff_6/in_2')
// (14, 22, 'neigh_op_lft_5')
// (14, 23, 'local_g2_5')
// (14, 23, 'lutff_0/in_1')
// (14, 23, 'neigh_op_bnl_5')

reg n1847 = 0;
// (12, 21, 'neigh_op_tnr_6')
// (12, 22, 'local_g2_6')
// (12, 22, 'lutff_5/in_1')
// (12, 22, 'neigh_op_rgt_6')
// (12, 23, 'neigh_op_bnr_6')
// (13, 21, 'neigh_op_top_6')
// (13, 22, 'lutff_6/out')
// (13, 23, 'neigh_op_bot_6')
// (14, 21, 'neigh_op_tnl_6')
// (14, 22, 'local_g0_6')
// (14, 22, 'lutff_1/in_1')
// (14, 22, 'neigh_op_lft_6')
// (14, 23, 'local_g3_6')
// (14, 23, 'lutff_5/in_2')
// (14, 23, 'neigh_op_bnl_6')

reg n1848 = 0;
// (12, 22, 'local_g2_7')
// (12, 22, 'lutff_4/in_1')
// (12, 22, 'neigh_op_tnr_7')
// (12, 23, 'neigh_op_rgt_7')
// (12, 24, 'neigh_op_bnr_7')
// (13, 22, 'neigh_op_top_7')
// (13, 23, 'lutff_7/out')
// (13, 24, 'neigh_op_bot_7')
// (14, 22, 'local_g3_7')
// (14, 22, 'lutff_1/in_3')
// (14, 22, 'neigh_op_tnl_7')
// (14, 23, 'local_g0_7')
// (14, 23, 'lutff_4/in_1')
// (14, 23, 'neigh_op_lft_7')
// (14, 24, 'neigh_op_bnl_7')

wire n1849;
// (12, 22, 'local_g3_6')
// (12, 22, 'lutff_7/in_0')
// (12, 22, 'neigh_op_tnr_6')
// (12, 23, 'neigh_op_rgt_6')
// (12, 24, 'neigh_op_bnr_6')
// (13, 22, 'neigh_op_top_6')
// (13, 23, 'lutff_6/out')
// (13, 24, 'neigh_op_bot_6')
// (14, 22, 'neigh_op_tnl_6')
// (14, 23, 'neigh_op_lft_6')
// (14, 24, 'neigh_op_bnl_6')

wire n1850;
// (12, 22, 'lutff_1/cout')
// (12, 22, 'lutff_2/in_3')

wire n1851;
// (12, 22, 'lutff_2/cout')
// (12, 22, 'lutff_3/in_3')

wire n1852;
// (12, 22, 'lutff_3/cout')
// (12, 22, 'lutff_4/in_3')

wire n1853;
// (12, 22, 'lutff_4/cout')
// (12, 22, 'lutff_5/in_3')

wire n1854;
// (12, 22, 'lutff_5/cout')
// (12, 22, 'lutff_6/in_3')

wire n1855;
// (12, 22, 'neigh_op_tnr_1')
// (12, 23, 'local_g2_1')
// (12, 23, 'lutff_4/in_3')
// (12, 23, 'neigh_op_rgt_1')
// (12, 24, 'neigh_op_bnr_1')
// (13, 22, 'neigh_op_top_1')
// (13, 23, 'lutff_1/out')
// (13, 24, 'neigh_op_bot_1')
// (14, 22, 'neigh_op_tnl_1')
// (14, 23, 'neigh_op_lft_1')
// (14, 24, 'neigh_op_bnl_1')

wire n1856;
// (12, 22, 'neigh_op_tnr_2')
// (12, 23, 'neigh_op_rgt_2')
// (12, 24, 'neigh_op_bnr_2')
// (13, 22, 'local_g1_2')
// (13, 22, 'lutff_2/in_3')
// (13, 22, 'neigh_op_top_2')
// (13, 23, 'lutff_2/out')
// (13, 24, 'neigh_op_bot_2')
// (14, 22, 'neigh_op_tnl_2')
// (14, 23, 'neigh_op_lft_2')
// (14, 24, 'neigh_op_bnl_2')

wire n1857;
// (12, 22, 'neigh_op_tnr_3')
// (12, 23, 'neigh_op_rgt_3')
// (12, 24, 'neigh_op_bnr_3')
// (13, 22, 'local_g0_3')
// (13, 22, 'lutff_4/in_3')
// (13, 22, 'neigh_op_top_3')
// (13, 23, 'lutff_3/out')
// (13, 24, 'neigh_op_bot_3')
// (14, 22, 'neigh_op_tnl_3')
// (14, 23, 'neigh_op_lft_3')
// (14, 24, 'neigh_op_bnl_3')

wire n1858;
// (12, 22, 'neigh_op_tnr_4')
// (12, 23, 'neigh_op_rgt_4')
// (12, 24, 'neigh_op_bnr_4')
// (13, 22, 'neigh_op_top_4')
// (13, 23, 'local_g1_4')
// (13, 23, 'lutff_4/out')
// (13, 23, 'lutff_7/in_0')
// (13, 24, 'neigh_op_bot_4')
// (14, 22, 'neigh_op_tnl_4')
// (14, 23, 'neigh_op_lft_4')
// (14, 24, 'neigh_op_bnl_4')

wire n1859;
// (12, 22, 'neigh_op_tnr_5')
// (12, 23, 'neigh_op_rgt_5')
// (12, 24, 'neigh_op_bnr_5')
// (13, 22, 'local_g0_5')
// (13, 22, 'lutff_6/in_3')
// (13, 22, 'neigh_op_top_5')
// (13, 23, 'lutff_5/out')
// (13, 24, 'neigh_op_bot_5')
// (14, 22, 'neigh_op_tnl_5')
// (14, 23, 'neigh_op_lft_5')
// (14, 24, 'neigh_op_bnl_5')

wire n1860;
// (13, 0, 'logic_op_tnr_0')
// (13, 1, 'neigh_op_rgt_0')
// (13, 1, 'sp4_r_v_b_0')
// (13, 2, 'neigh_op_bnr_0')
// (13, 2, 'sp4_r_v_b_38')
// (13, 3, 'sp4_r_v_b_27')
// (13, 4, 'sp4_r_v_b_14')
// (13, 5, 'sp4_r_v_b_3')
// (13, 6, 'sp4_r_v_b_43')
// (13, 7, 'sp4_r_v_b_30')
// (13, 8, 'local_g3_3')
// (13, 8, 'lutff_global/cen')
// (13, 8, 'sp4_r_v_b_19')
// (13, 9, 'sp4_r_v_b_6')
// (14, 0, 'logic_op_top_0')
// (14, 0, 'span4_vert_0')
// (14, 1, 'local_g0_2')
// (14, 1, 'lutff_0/out')
// (14, 1, 'lutff_global/cen')
// (14, 1, 'sp4_r_v_b_33')
// (14, 1, 'sp4_v_b_0')
// (14, 1, 'sp4_v_t_38')
// (14, 2, 'neigh_op_bot_0')
// (14, 2, 'sp4_r_v_b_20')
// (14, 2, 'sp4_v_b_38')
// (14, 3, 'sp4_r_v_b_9')
// (14, 3, 'sp4_v_b_27')
// (14, 4, 'sp4_v_b_14')
// (14, 5, 'sp4_v_b_3')
// (14, 5, 'sp4_v_t_43')
// (14, 6, 'sp4_v_b_43')
// (14, 7, 'sp4_v_b_30')
// (14, 8, 'sp4_v_b_19')
// (14, 9, 'sp4_v_b_6')
// (15, 0, 'logic_op_tnl_0')
// (15, 0, 'span4_vert_33')
// (15, 1, 'neigh_op_lft_0')
// (15, 1, 'sp4_v_b_33')
// (15, 2, 'neigh_op_bnl_0')
// (15, 2, 'sp4_v_b_20')
// (15, 3, 'sp4_v_b_9')

reg n1861 = 0;
// (13, 0, 'logic_op_tnr_2')
// (13, 1, 'neigh_op_rgt_2')
// (13, 2, 'neigh_op_bnr_2')
// (14, 0, 'logic_op_top_2')
// (14, 1, 'lutff_2/out')
// (14, 2, 'local_g0_2')
// (14, 2, 'lutff_1/in_3')
// (14, 2, 'neigh_op_bot_2')
// (15, 0, 'logic_op_tnl_2')
// (15, 1, 'neigh_op_lft_2')
// (15, 2, 'neigh_op_bnl_2')

wire n1862;
// (13, 1, 'lutff_7/cout')
// (13, 2, 'carry_in')
// (13, 2, 'carry_in_mux')
// (13, 2, 'lutff_0/in_3')

wire n1863;
// (13, 1, 'neigh_op_tnr_2')
// (13, 2, 'neigh_op_rgt_2')
// (13, 2, 'sp4_r_v_b_36')
// (13, 3, 'local_g0_2')
// (13, 3, 'lutff_0/in_2')
// (13, 3, 'lutff_6/in_0')
// (13, 3, 'neigh_op_bnr_2')
// (13, 3, 'sp4_r_v_b_25')
// (13, 4, 'sp4_r_v_b_12')
// (13, 5, 'sp4_r_v_b_1')
// (14, 1, 'neigh_op_top_2')
// (14, 1, 'sp4_v_t_36')
// (14, 2, 'local_g2_2')
// (14, 2, 'lutff_2/out')
// (14, 2, 'lutff_5/in_3')
// (14, 2, 'sp4_v_b_36')
// (14, 3, 'local_g0_2')
// (14, 3, 'lutff_0/in_2')
// (14, 3, 'neigh_op_bot_2')
// (14, 3, 'sp4_v_b_25')
// (14, 4, 'local_g1_4')
// (14, 4, 'lutff_7/in_2')
// (14, 4, 'sp4_v_b_12')
// (14, 5, 'sp4_v_b_1')
// (15, 1, 'neigh_op_tnl_2')
// (15, 2, 'local_g1_2')
// (15, 2, 'lutff_1/in_0')
// (15, 2, 'lutff_3/in_0')
// (15, 2, 'lutff_7/in_2')
// (15, 2, 'neigh_op_lft_2')
// (15, 3, 'neigh_op_bnl_2')

reg n1864 = 0;
// (13, 1, 'neigh_op_tnr_3')
// (13, 2, 'neigh_op_rgt_3')
// (13, 3, 'neigh_op_bnr_3')
// (14, 1, 'neigh_op_top_3')
// (14, 2, 'local_g0_3')
// (14, 2, 'lutff_3/out')
// (14, 2, 'lutff_6/in_1')
// (14, 3, 'neigh_op_bot_3')
// (15, 1, 'neigh_op_tnl_3')
// (15, 2, 'neigh_op_lft_3')
// (15, 3, 'neigh_op_bnl_3')

wire n1865;
// (13, 1, 'neigh_op_tnr_4')
// (13, 1, 'sp4_r_v_b_37')
// (13, 2, 'neigh_op_rgt_4')
// (13, 2, 'sp4_r_v_b_24')
// (13, 3, 'neigh_op_bnr_4')
// (13, 3, 'sp4_r_v_b_13')
// (13, 4, 'sp4_r_v_b_0')
// (14, 0, 'span4_vert_37')
// (14, 1, 'neigh_op_top_4')
// (14, 1, 'sp4_v_b_37')
// (14, 2, 'lutff_4/out')
// (14, 2, 'sp4_v_b_24')
// (14, 3, 'neigh_op_bot_4')
// (14, 3, 'sp4_v_b_13')
// (14, 4, 'local_g1_0')
// (14, 4, 'lutff_3/in_0')
// (14, 4, 'sp4_v_b_0')
// (15, 1, 'neigh_op_tnl_4')
// (15, 2, 'neigh_op_lft_4')
// (15, 3, 'neigh_op_bnl_4')

wire n1866;
// (13, 1, 'neigh_op_tnr_5')
// (13, 2, 'neigh_op_rgt_5')
// (13, 3, 'local_g1_5')
// (13, 3, 'lutff_4/in_0')
// (13, 3, 'neigh_op_bnr_5')
// (14, 1, 'neigh_op_top_5')
// (14, 2, 'lutff_5/out')
// (14, 3, 'neigh_op_bot_5')
// (15, 1, 'neigh_op_tnl_5')
// (15, 2, 'neigh_op_lft_5')
// (15, 3, 'neigh_op_bnl_5')

wire n1867;
// (13, 1, 'neigh_op_tnr_7')
// (13, 2, 'neigh_op_rgt_7')
// (13, 3, 'neigh_op_bnr_7')
// (14, 1, 'neigh_op_top_7')
// (14, 2, 'local_g0_7')
// (14, 2, 'lutff_4/in_1')
// (14, 2, 'lutff_7/out')
// (14, 3, 'neigh_op_bot_7')
// (15, 1, 'neigh_op_tnl_7')
// (15, 2, 'neigh_op_lft_7')
// (15, 3, 'neigh_op_bnl_7')

reg n1868 = 0;
// (13, 1, 'sp4_r_v_b_34')
// (13, 2, 'local_g3_7')
// (13, 2, 'lutff_1/in_1')
// (13, 2, 'sp4_r_v_b_23')
// (13, 3, 'sp12_h_r_1')
// (13, 3, 'sp12_v_t_22')
// (13, 3, 'sp4_r_v_b_10')
// (13, 4, 'sp12_v_b_22')
// (13, 5, 'sp12_v_b_21')
// (13, 6, 'sp12_v_b_18')
// (13, 7, 'sp12_v_b_17')
// (13, 8, 'sp12_v_b_14')
// (13, 9, 'sp12_v_b_13')
// (13, 10, 'sp12_v_b_10')
// (13, 11, 'sp12_v_b_9')
// (13, 12, 'sp12_v_b_6')
// (13, 13, 'sp12_v_b_5')
// (13, 14, 'sp12_v_b_2')
// (13, 15, 'local_g3_1')
// (13, 15, 'lutff_5/in_1')
// (13, 15, 'sp12_v_b_1')
// (14, 0, 'span4_vert_34')
// (14, 1, 'sp4_v_b_34')
// (14, 2, 'sp4_v_b_23')
// (14, 3, 'sp12_h_r_2')
// (14, 3, 'sp4_h_r_5')
// (14, 3, 'sp4_v_b_10')
// (15, 3, 'sp12_h_r_5')
// (15, 3, 'sp4_h_r_16')
// (15, 5, 'sp4_h_r_11')
// (16, 3, 'sp12_h_r_6')
// (16, 3, 'sp4_h_r_29')
// (16, 4, 'sp4_r_v_b_42')
// (16, 5, 'local_g0_6')
// (16, 5, 'lutff_4/in_0')
// (16, 5, 'sp4_h_r_22')
// (16, 5, 'sp4_r_v_b_31')
// (16, 6, 'sp4_r_v_b_18')
// (16, 7, 'sp4_r_v_b_7')
// (17, 2, 'neigh_op_tnr_1')
// (17, 3, 'neigh_op_rgt_1')
// (17, 3, 'sp12_h_r_9')
// (17, 3, 'sp4_h_r_40')
// (17, 3, 'sp4_h_r_7')
// (17, 3, 'sp4_v_t_42')
// (17, 4, 'neigh_op_bnr_1')
// (17, 4, 'sp4_v_b_42')
// (17, 5, 'sp4_h_r_35')
// (17, 5, 'sp4_v_b_31')
// (17, 6, 'sp4_v_b_18')
// (17, 7, 'local_g0_7')
// (17, 7, 'lutff_2/in_1')
// (17, 7, 'sp4_v_b_7')
// (18, 2, 'neigh_op_top_1')
// (18, 2, 'sp4_r_v_b_46')
// (18, 3, 'local_g1_1')
// (18, 3, 'lutff_1/in_1')
// (18, 3, 'lutff_1/out')
// (18, 3, 'sp12_h_r_10')
// (18, 3, 'sp4_h_l_40')
// (18, 3, 'sp4_h_r_18')
// (18, 3, 'sp4_h_r_2')
// (18, 3, 'sp4_r_v_b_35')
// (18, 4, 'neigh_op_bot_1')
// (18, 4, 'sp4_r_v_b_22')
// (18, 5, 'sp4_h_r_46')
// (18, 5, 'sp4_r_v_b_11')
// (19, 1, 'sp4_v_t_46')
// (19, 2, 'neigh_op_tnl_1')
// (19, 2, 'sp4_v_b_46')
// (19, 3, 'neigh_op_lft_1')
// (19, 3, 'sp12_h_r_13')
// (19, 3, 'sp4_h_r_15')
// (19, 3, 'sp4_h_r_31')
// (19, 3, 'sp4_v_b_35')
// (19, 4, 'neigh_op_bnl_1')
// (19, 4, 'sp4_v_b_22')
// (19, 5, 'sp4_h_l_46')
// (19, 5, 'sp4_v_b_11')
// (20, 3, 'sp12_h_r_14')
// (20, 3, 'sp4_h_r_26')
// (20, 3, 'sp4_h_r_42')
// (21, 3, 'sp12_h_r_17')
// (21, 3, 'sp4_h_l_42')
// (21, 3, 'sp4_h_r_39')
// (22, 3, 'sp12_h_r_18')
// (22, 3, 'sp4_h_l_39')
// (23, 3, 'sp12_h_r_21')
// (24, 3, 'sp12_h_r_22')
// (25, 3, 'sp12_h_l_22')

wire n1869;
// (13, 1, 'sp4_r_v_b_47')
// (13, 2, 'sp4_r_v_b_34')
// (13, 3, 'sp4_r_v_b_23')
// (13, 4, 'sp4_r_v_b_10')
// (14, 0, 'span4_vert_47')
// (14, 1, 'sp4_v_b_47')
// (14, 2, 'sp4_v_b_34')
// (14, 3, 'neigh_op_tnr_0')
// (14, 3, 'sp4_v_b_23')
// (14, 4, 'local_g0_2')
// (14, 4, 'lutff_global/cen')
// (14, 4, 'neigh_op_rgt_0')
// (14, 4, 'sp4_h_r_5')
// (14, 4, 'sp4_v_b_10')
// (14, 5, 'neigh_op_bnr_0')
// (14, 5, 'sp4_r_v_b_43')
// (14, 6, 'sp4_r_v_b_30')
// (14, 7, 'sp4_r_v_b_19')
// (14, 8, 'sp4_r_v_b_6')
// (15, 2, 'sp4_r_v_b_41')
// (15, 3, 'neigh_op_top_0')
// (15, 3, 'sp4_r_v_b_28')
// (15, 4, 'lutff_0/out')
// (15, 4, 'sp4_h_r_0')
// (15, 4, 'sp4_h_r_16')
// (15, 4, 'sp4_r_v_b_17')
// (15, 4, 'sp4_v_t_43')
// (15, 5, 'local_g3_3')
// (15, 5, 'lutff_global/cen')
// (15, 5, 'neigh_op_bot_0')
// (15, 5, 'sp4_r_v_b_4')
// (15, 5, 'sp4_v_b_43')
// (15, 6, 'sp4_v_b_30')
// (15, 7, 'sp4_v_b_19')
// (15, 8, 'sp4_v_b_6')
// (16, 1, 'sp4_v_t_41')
// (16, 2, 'sp4_v_b_41')
// (16, 3, 'neigh_op_tnl_0')
// (16, 3, 'sp4_v_b_28')
// (16, 4, 'neigh_op_lft_0')
// (16, 4, 'sp4_h_r_13')
// (16, 4, 'sp4_h_r_29')
// (16, 4, 'sp4_v_b_17')
// (16, 5, 'local_g0_2')
// (16, 5, 'lutff_global/cen')
// (16, 5, 'neigh_op_bnl_0')
// (16, 5, 'sp4_h_r_10')
// (16, 5, 'sp4_v_b_4')
// (17, 4, 'sp4_h_r_24')
// (17, 4, 'sp4_h_r_40')
// (17, 5, 'sp4_h_r_23')
// (18, 4, 'sp4_h_l_40')
// (18, 4, 'sp4_h_r_37')
// (18, 5, 'sp4_h_r_34')
// (19, 4, 'sp4_h_l_37')
// (19, 5, 'sp4_h_r_47')
// (20, 5, 'sp4_h_l_47')

wire n1870;
// (13, 2, 'neigh_op_tnr_0')
// (13, 3, 'neigh_op_rgt_0')
// (13, 4, 'neigh_op_bnr_0')
// (14, 2, 'neigh_op_top_0')
// (14, 3, 'local_g1_0')
// (14, 3, 'lutff_0/out')
// (14, 3, 'lutff_4/in_3')
// (14, 4, 'neigh_op_bot_0')
// (15, 2, 'neigh_op_tnl_0')
// (15, 3, 'neigh_op_lft_0')
// (15, 4, 'neigh_op_bnl_0')

reg n1871 = 0;
// (13, 2, 'neigh_op_tnr_2')
// (13, 3, 'neigh_op_rgt_2')
// (13, 3, 'sp4_r_v_b_36')
// (13, 4, 'neigh_op_bnr_2')
// (13, 4, 'sp4_r_v_b_25')
// (13, 5, 'sp4_r_v_b_12')
// (13, 6, 'local_g1_1')
// (13, 6, 'lutff_3/in_3')
// (13, 6, 'lutff_5/in_3')
// (13, 6, 'sp4_r_v_b_1')
// (14, 2, 'neigh_op_top_2')
// (14, 2, 'sp4_v_t_36')
// (14, 3, 'lutff_2/out')
// (14, 3, 'sp4_v_b_36')
// (14, 4, 'local_g1_2')
// (14, 4, 'lutff_4/in_3')
// (14, 4, 'neigh_op_bot_2')
// (14, 4, 'sp4_v_b_25')
// (14, 5, 'sp4_v_b_12')
// (14, 6, 'sp4_v_b_1')
// (15, 2, 'neigh_op_tnl_2')
// (15, 3, 'neigh_op_lft_2')
// (15, 4, 'neigh_op_bnl_2')

wire n1872;
// (13, 2, 'neigh_op_tnr_4')
// (13, 3, 'neigh_op_rgt_4')
// (13, 4, 'local_g0_4')
// (13, 4, 'lutff_4/in_2')
// (13, 4, 'neigh_op_bnr_4')
// (14, 2, 'neigh_op_top_4')
// (14, 3, 'lutff_4/out')
// (14, 4, 'neigh_op_bot_4')
// (15, 2, 'neigh_op_tnl_4')
// (15, 3, 'neigh_op_lft_4')
// (15, 4, 'neigh_op_bnl_4')

wire n1873;
// (13, 2, 'neigh_op_tnr_5')
// (13, 3, 'neigh_op_rgt_5')
// (13, 4, 'neigh_op_bnr_5')
// (14, 2, 'neigh_op_top_5')
// (14, 3, 'lutff_5/out')
// (14, 4, 'local_g0_5')
// (14, 4, 'lutff_6/in_1')
// (14, 4, 'neigh_op_bot_5')
// (15, 2, 'neigh_op_tnl_5')
// (15, 3, 'neigh_op_lft_5')
// (15, 4, 'neigh_op_bnl_5')

wire n1874;
// (13, 2, 'neigh_op_tnr_7')
// (13, 3, 'local_g3_7')
// (13, 3, 'lutff_1/in_1')
// (13, 3, 'lutff_2/in_2')
// (13, 3, 'neigh_op_rgt_7')
// (13, 4, 'local_g1_7')
// (13, 4, 'lutff_0/in_0')
// (13, 4, 'neigh_op_bnr_7')
// (14, 2, 'local_g1_7')
// (14, 2, 'lutff_7/in_3')
// (14, 2, 'neigh_op_top_7')
// (14, 3, 'lutff_7/out')
// (14, 4, 'local_g0_7')
// (14, 4, 'lutff_4/in_1')
// (14, 4, 'neigh_op_bot_7')
// (15, 2, 'local_g3_7')
// (15, 2, 'lutff_1/in_1')
// (15, 2, 'neigh_op_tnl_7')
// (15, 3, 'neigh_op_lft_7')
// (15, 4, 'local_g3_7')
// (15, 4, 'lutff_5/in_1')
// (15, 4, 'neigh_op_bnl_7')

wire n1875;
// (13, 2, 'sp4_r_v_b_40')
// (13, 3, 'local_g3_0')
// (13, 3, 'lutff_6/in_1')
// (13, 3, 'lutff_7/in_0')
// (13, 3, 'neigh_op_tnr_0')
// (13, 3, 'sp4_r_v_b_29')
// (13, 4, 'neigh_op_rgt_0')
// (13, 4, 'sp4_r_v_b_16')
// (13, 5, 'neigh_op_bnr_0')
// (13, 5, 'sp4_r_v_b_5')
// (14, 1, 'sp4_v_t_40')
// (14, 2, 'local_g2_0')
// (14, 2, 'lutff_4/in_0')
// (14, 2, 'sp4_r_v_b_41')
// (14, 2, 'sp4_v_b_40')
// (14, 3, 'local_g0_0')
// (14, 3, 'lutff_4/in_0')
// (14, 3, 'neigh_op_top_0')
// (14, 3, 'sp4_r_v_b_28')
// (14, 3, 'sp4_v_b_29')
// (14, 4, 'local_g0_0')
// (14, 4, 'lutff_0/out')
// (14, 4, 'lutff_4/in_2')
// (14, 4, 'sp4_r_v_b_17')
// (14, 4, 'sp4_v_b_16')
// (14, 5, 'neigh_op_bot_0')
// (14, 5, 'sp4_r_v_b_4')
// (14, 5, 'sp4_v_b_5')
// (15, 1, 'local_g0_4')
// (15, 1, 'lutff_4/in_2')
// (15, 1, 'sp4_h_r_4')
// (15, 1, 'sp4_v_t_41')
// (15, 2, 'local_g2_1')
// (15, 2, 'lutff_5/in_2')
// (15, 2, 'sp4_v_b_41')
// (15, 3, 'local_g3_0')
// (15, 3, 'lutff_6/in_1')
// (15, 3, 'neigh_op_tnl_0')
// (15, 3, 'sp4_v_b_28')
// (15, 4, 'local_g0_0')
// (15, 4, 'lutff_4/in_2')
// (15, 4, 'neigh_op_lft_0')
// (15, 4, 'sp4_v_b_17')
// (15, 5, 'neigh_op_bnl_0')
// (15, 5, 'sp4_v_b_4')
// (16, 1, 'sp4_h_r_17')
// (17, 1, 'sp4_h_r_28')
// (18, 1, 'sp4_h_r_41')
// (19, 1, 'sp4_h_l_41')

reg n1876 = 0;
// (13, 2, 'sp4_r_v_b_42')
// (13, 3, 'neigh_op_tnr_1')
// (13, 3, 'sp4_r_v_b_31')
// (13, 4, 'local_g3_1')
// (13, 4, 'lutff_2/in_0')
// (13, 4, 'neigh_op_rgt_1')
// (13, 4, 'sp4_r_v_b_18')
// (13, 5, 'neigh_op_bnr_1')
// (13, 5, 'sp4_r_v_b_7')
// (13, 6, 'sp4_r_v_b_38')
// (13, 7, 'local_g1_3')
// (13, 7, 'lutff_5/in_3')
// (13, 7, 'lutff_7/in_1')
// (13, 7, 'sp4_r_v_b_27')
// (13, 8, 'sp4_r_v_b_14')
// (13, 9, 'sp4_r_v_b_3')
// (14, 1, 'sp4_r_v_b_38')
// (14, 1, 'sp4_v_t_42')
// (14, 2, 'sp4_r_v_b_27')
// (14, 2, 'sp4_v_b_42')
// (14, 3, 'neigh_op_top_1')
// (14, 3, 'sp4_r_v_b_14')
// (14, 3, 'sp4_v_b_31')
// (14, 4, 'lutff_1/out')
// (14, 4, 'sp4_r_v_b_3')
// (14, 4, 'sp4_v_b_18')
// (14, 5, 'neigh_op_bot_1')
// (14, 5, 'sp4_r_v_b_38')
// (14, 5, 'sp4_v_b_7')
// (14, 5, 'sp4_v_t_38')
// (14, 6, 'sp4_r_v_b_27')
// (14, 6, 'sp4_v_b_38')
// (14, 7, 'sp4_r_v_b_14')
// (14, 7, 'sp4_v_b_27')
// (14, 8, 'sp4_r_v_b_3')
// (14, 8, 'sp4_v_b_14')
// (14, 9, 'sp4_v_b_3')
// (15, 0, 'span4_vert_38')
// (15, 1, 'sp4_v_b_38')
// (15, 2, 'sp4_v_b_27')
// (15, 3, 'neigh_op_tnl_1')
// (15, 3, 'sp4_v_b_14')
// (15, 4, 'neigh_op_lft_1')
// (15, 4, 'sp4_v_b_3')
// (15, 4, 'sp4_v_t_38')
// (15, 5, 'local_g2_1')
// (15, 5, 'lutff_2/in_1')
// (15, 5, 'neigh_op_bnl_1')
// (15, 5, 'sp4_v_b_38')
// (15, 6, 'sp4_v_b_27')
// (15, 7, 'local_g0_6')
// (15, 7, 'lutff_4/in_2')
// (15, 7, 'sp4_v_b_14')
// (15, 8, 'sp4_v_b_3')

reg n1877 = 0;
// (13, 2, 'sp4_r_v_b_46')
// (13, 3, 'sp4_r_v_b_35')
// (13, 4, 'local_g3_6')
// (13, 4, 'lutff_3/in_2')
// (13, 4, 'sp4_r_v_b_22')
// (13, 5, 'sp4_r_v_b_11')
// (13, 6, 'local_g3_6')
// (13, 6, 'lutff_1/in_0')
// (13, 6, 'sp4_r_v_b_46')
// (13, 7, 'sp4_r_v_b_35')
// (13, 8, 'sp4_r_v_b_22')
// (13, 9, 'sp4_r_v_b_11')
// (14, 1, 'sp4_v_t_46')
// (14, 2, 'sp4_v_b_46')
// (14, 3, 'sp4_v_b_35')
// (14, 4, 'neigh_op_tnr_3')
// (14, 4, 'sp4_v_b_22')
// (14, 5, 'neigh_op_rgt_3')
// (14, 5, 'sp4_h_r_11')
// (14, 5, 'sp4_v_b_11')
// (14, 5, 'sp4_v_t_46')
// (14, 6, 'local_g1_3')
// (14, 6, 'lutff_1/in_3')
// (14, 6, 'neigh_op_bnr_3')
// (14, 6, 'sp4_v_b_46')
// (14, 7, 'sp4_v_b_35')
// (14, 8, 'sp4_v_b_22')
// (14, 9, 'sp4_v_b_11')
// (15, 4, 'neigh_op_top_3')
// (15, 5, 'lutff_3/out')
// (15, 5, 'sp4_h_r_22')
// (15, 5, 'sp4_r_v_b_39')
// (15, 6, 'neigh_op_bot_3')
// (15, 6, 'sp4_r_v_b_26')
// (15, 7, 'sp4_r_v_b_15')
// (15, 8, 'sp4_r_v_b_2')
// (16, 4, 'neigh_op_tnl_3')
// (16, 4, 'sp4_v_t_39')
// (16, 5, 'neigh_op_lft_3')
// (16, 5, 'sp4_h_r_35')
// (16, 5, 'sp4_v_b_39')
// (16, 6, 'neigh_op_bnl_3')
// (16, 6, 'sp4_v_b_26')
// (16, 7, 'local_g1_7')
// (16, 7, 'lutff_0/in_2')
// (16, 7, 'sp4_v_b_15')
// (16, 8, 'sp4_v_b_2')
// (17, 5, 'sp4_h_r_46')
// (18, 5, 'sp4_h_l_46')

wire n1878;
// (13, 3, 'neigh_op_tnr_2')
// (13, 4, 'neigh_op_rgt_2')
// (13, 5, 'neigh_op_bnr_2')
// (14, 3, 'neigh_op_top_2')
// (14, 4, 'local_g3_2')
// (14, 4, 'lutff_2/out')
// (14, 4, 'lutff_6/in_3')
// (14, 5, 'neigh_op_bot_2')
// (15, 3, 'neigh_op_tnl_2')
// (15, 4, 'neigh_op_lft_2')
// (15, 5, 'neigh_op_bnl_2')

wire n1879;
// (13, 3, 'neigh_op_tnr_3')
// (13, 4, 'neigh_op_rgt_3')
// (13, 5, 'neigh_op_bnr_3')
// (14, 3, 'neigh_op_top_3')
// (14, 4, 'lutff_3/out')
// (14, 5, 'local_g1_3')
// (14, 5, 'lutff_4/in_0')
// (14, 5, 'neigh_op_bot_3')
// (15, 3, 'neigh_op_tnl_3')
// (15, 4, 'neigh_op_lft_3')
// (15, 5, 'neigh_op_bnl_3')

wire n1880;
// (13, 3, 'neigh_op_tnr_4')
// (13, 4, 'local_g3_4')
// (13, 4, 'lutff_6/in_3')
// (13, 4, 'neigh_op_rgt_4')
// (13, 5, 'neigh_op_bnr_4')
// (14, 3, 'neigh_op_top_4')
// (14, 4, 'lutff_4/out')
// (14, 5, 'neigh_op_bot_4')
// (15, 3, 'neigh_op_tnl_4')
// (15, 4, 'neigh_op_lft_4')
// (15, 5, 'neigh_op_bnl_4')

wire n1881;
// (13, 3, 'neigh_op_tnr_7')
// (13, 4, 'local_g2_7')
// (13, 4, 'lutff_6/in_1')
// (13, 4, 'neigh_op_rgt_7')
// (13, 5, 'neigh_op_bnr_7')
// (14, 3, 'neigh_op_top_7')
// (14, 4, 'lutff_7/out')
// (14, 5, 'neigh_op_bot_7')
// (15, 3, 'neigh_op_tnl_7')
// (15, 4, 'neigh_op_lft_7')
// (15, 5, 'neigh_op_bnl_7')

reg n1882 = 0;
// (13, 3, 'sp4_r_v_b_38')
// (13, 4, 'sp4_r_v_b_27')
// (13, 5, 'sp4_r_v_b_14')
// (13, 6, 'sp4_r_v_b_3')
// (13, 7, 'sp4_r_v_b_38')
// (13, 8, 'sp4_r_v_b_27')
// (13, 9, 'sp4_r_v_b_14')
// (13, 10, 'sp4_r_v_b_3')
// (14, 1, 'neigh_op_tnr_2')
// (14, 2, 'neigh_op_rgt_2')
// (14, 2, 'sp4_h_r_9')
// (14, 2, 'sp4_v_t_38')
// (14, 3, 'local_g1_2')
// (14, 3, 'lutff_0/in_1')
// (14, 3, 'neigh_op_bnr_2')
// (14, 3, 'sp4_v_b_38')
// (14, 4, 'sp4_v_b_27')
// (14, 5, 'sp4_v_b_14')
// (14, 6, 'local_g0_3')
// (14, 6, 'lutff_4/in_3')
// (14, 6, 'sp4_v_b_3')
// (14, 6, 'sp4_v_t_38')
// (14, 7, 'sp4_v_b_38')
// (14, 8, 'sp4_v_b_27')
// (14, 9, 'sp4_v_b_14')
// (14, 10, 'local_g1_3')
// (14, 10, 'lutff_7/in_3')
// (14, 10, 'sp4_v_b_3')
// (15, 0, 'span12_vert_23')
// (15, 1, 'neigh_op_top_2')
// (15, 1, 'sp12_v_b_23')
// (15, 2, 'lutff_2/out')
// (15, 2, 'sp12_v_b_20')
// (15, 2, 'sp4_h_r_20')
// (15, 3, 'neigh_op_bot_2')
// (15, 3, 'sp12_v_b_19')
// (15, 4, 'sp12_v_b_16')
// (15, 5, 'sp12_v_b_15')
// (15, 6, 'sp12_v_b_12')
// (15, 7, 'sp12_v_b_11')
// (15, 8, 'sp12_v_b_8')
// (15, 9, 'local_g3_7')
// (15, 9, 'lutff_1/in_3')
// (15, 9, 'sp12_v_b_7')
// (15, 10, 'local_g3_4')
// (15, 10, 'lutff_7/in_2')
// (15, 10, 'sp12_v_b_4')
// (15, 11, 'sp12_v_b_3')
// (15, 12, 'sp12_v_b_0')
// (16, 1, 'neigh_op_tnl_2')
// (16, 2, 'neigh_op_lft_2')
// (16, 2, 'sp4_h_r_33')
// (16, 3, 'neigh_op_bnl_2')
// (17, 2, 'sp4_h_r_44')
// (18, 2, 'sp4_h_l_44')

reg n1883 = 0;
// (13, 3, 'sp4_r_v_b_40')
// (13, 4, 'sp4_r_v_b_29')
// (13, 5, 'sp4_r_v_b_16')
// (13, 6, 'sp4_r_v_b_5')
// (14, 1, 'neigh_op_tnr_0')
// (14, 2, 'local_g3_0')
// (14, 2, 'lutff_5/in_2')
// (14, 2, 'neigh_op_rgt_0')
// (14, 2, 'sp4_h_r_5')
// (14, 2, 'sp4_v_t_40')
// (14, 3, 'neigh_op_bnr_0')
// (14, 3, 'sp4_v_b_40')
// (14, 4, 'sp4_v_b_29')
// (14, 5, 'sp4_v_b_16')
// (14, 6, 'local_g1_5')
// (14, 6, 'lutff_0/in_0')
// (14, 6, 'lutff_6/in_2')
// (14, 6, 'sp4_v_b_5')
// (15, 1, 'neigh_op_top_0')
// (15, 1, 'sp4_r_v_b_28')
// (15, 2, 'lutff_0/out')
// (15, 2, 'sp4_h_r_16')
// (15, 2, 'sp4_r_v_b_17')
// (15, 3, 'neigh_op_bot_0')
// (15, 3, 'sp4_r_v_b_4')
// (15, 4, 'sp4_r_v_b_41')
// (15, 5, 'sp4_r_v_b_28')
// (15, 6, 'sp4_r_v_b_17')
// (15, 7, 'sp4_r_v_b_4')
// (16, 0, 'span4_vert_28')
// (16, 1, 'neigh_op_tnl_0')
// (16, 1, 'sp4_v_b_28')
// (16, 2, 'neigh_op_lft_0')
// (16, 2, 'sp4_h_r_29')
// (16, 2, 'sp4_v_b_17')
// (16, 3, 'neigh_op_bnl_0')
// (16, 3, 'sp4_v_b_4')
// (16, 3, 'sp4_v_t_41')
// (16, 4, 'sp4_v_b_41')
// (16, 5, 'sp4_v_b_28')
// (16, 6, 'local_g0_1')
// (16, 6, 'lutff_7/in_0')
// (16, 6, 'sp4_v_b_17')
// (16, 7, 'local_g0_4')
// (16, 7, 'lutff_4/in_0')
// (16, 7, 'sp4_v_b_4')
// (17, 2, 'sp4_h_r_40')
// (18, 2, 'sp4_h_l_40')

reg n1884 = 0;
// (13, 3, 'sp4_r_v_b_47')
// (13, 4, 'sp4_h_r_4')
// (13, 4, 'sp4_r_v_b_34')
// (13, 5, 'sp4_r_v_b_23')
// (13, 6, 'sp4_r_v_b_10')
// (14, 2, 'sp4_h_r_10')
// (14, 2, 'sp4_v_t_47')
// (14, 3, 'sp4_v_b_47')
// (14, 4, 'local_g0_1')
// (14, 4, 'lutff_7/in_0')
// (14, 4, 'sp4_h_r_17')
// (14, 4, 'sp4_v_b_34')
// (14, 5, 'sp4_v_b_23')
// (14, 6, 'local_g1_2')
// (14, 6, 'lutff_3/in_2')
// (14, 6, 'sp4_v_b_10')
// (15, 1, 'neigh_op_tnr_1')
// (15, 2, 'neigh_op_rgt_1')
// (15, 2, 'sp4_h_r_23')
// (15, 3, 'neigh_op_bnr_1')
// (15, 3, 'sp4_r_v_b_45')
// (15, 4, 'sp4_h_r_28')
// (15, 4, 'sp4_r_v_b_32')
// (15, 5, 'sp4_r_v_b_21')
// (15, 6, 'sp4_r_v_b_8')
// (16, 1, 'neigh_op_top_1')
// (16, 1, 'sp4_r_v_b_46')
// (16, 2, 'lutff_1/out')
// (16, 2, 'sp4_h_r_2')
// (16, 2, 'sp4_h_r_34')
// (16, 2, 'sp4_r_v_b_35')
// (16, 2, 'sp4_v_t_45')
// (16, 3, 'neigh_op_bot_1')
// (16, 3, 'sp4_r_v_b_22')
// (16, 3, 'sp4_v_b_45')
// (16, 4, 'sp4_h_r_41')
// (16, 4, 'sp4_r_v_b_11')
// (16, 4, 'sp4_v_b_32')
// (16, 5, 'local_g1_5')
// (16, 5, 'lutff_6/in_2')
// (16, 5, 'sp4_r_v_b_46')
// (16, 5, 'sp4_v_b_21')
// (16, 6, 'local_g1_0')
// (16, 6, 'lutff_0/in_3')
// (16, 6, 'sp4_r_v_b_35')
// (16, 6, 'sp4_v_b_8')
// (16, 7, 'local_g3_6')
// (16, 7, 'lutff_5/in_2')
// (16, 7, 'sp4_r_v_b_22')
// (16, 8, 'sp4_r_v_b_11')
// (17, 0, 'span4_vert_46')
// (17, 1, 'neigh_op_tnl_1')
// (17, 1, 'sp4_v_b_46')
// (17, 2, 'neigh_op_lft_1')
// (17, 2, 'sp4_h_r_15')
// (17, 2, 'sp4_h_r_47')
// (17, 2, 'sp4_v_b_35')
// (17, 3, 'neigh_op_bnl_1')
// (17, 3, 'sp4_v_b_22')
// (17, 4, 'sp4_h_l_41')
// (17, 4, 'sp4_v_b_11')
// (17, 4, 'sp4_v_t_46')
// (17, 5, 'sp4_v_b_46')
// (17, 6, 'sp4_v_b_35')
// (17, 7, 'sp4_v_b_22')
// (17, 8, 'sp4_v_b_11')
// (18, 2, 'sp4_h_l_47')
// (18, 2, 'sp4_h_r_26')
// (19, 2, 'sp4_h_r_39')
// (20, 2, 'sp4_h_l_39')

reg n1885 = 0;
// (13, 4, 'neigh_op_tnr_0')
// (13, 4, 'sp4_r_v_b_45')
// (13, 5, 'local_g3_0')
// (13, 5, 'lutff_4/in_1')
// (13, 5, 'neigh_op_rgt_0')
// (13, 5, 'sp4_r_v_b_32')
// (13, 6, 'neigh_op_bnr_0')
// (13, 6, 'sp4_r_v_b_21')
// (13, 7, 'local_g2_0')
// (13, 7, 'lutff_2/in_2')
// (13, 7, 'sp4_r_v_b_8')
// (13, 8, 'sp4_r_v_b_41')
// (13, 9, 'local_g0_4')
// (13, 9, 'lutff_6/in_0')
// (13, 9, 'sp4_r_v_b_28')
// (13, 10, 'sp4_r_v_b_17')
// (13, 11, 'sp4_r_v_b_4')
// (14, 3, 'sp4_v_t_45')
// (14, 4, 'neigh_op_top_0')
// (14, 4, 'sp4_r_v_b_44')
// (14, 4, 'sp4_v_b_45')
// (14, 5, 'lutff_0/out')
// (14, 5, 'sp4_r_v_b_33')
// (14, 5, 'sp4_v_b_32')
// (14, 6, 'neigh_op_bot_0')
// (14, 6, 'sp4_r_v_b_20')
// (14, 6, 'sp4_v_b_21')
// (14, 7, 'sp4_h_r_8')
// (14, 7, 'sp4_r_v_b_9')
// (14, 7, 'sp4_v_b_8')
// (14, 7, 'sp4_v_t_41')
// (14, 8, 'sp4_r_v_b_40')
// (14, 8, 'sp4_v_b_41')
// (14, 9, 'sp4_r_v_b_29')
// (14, 9, 'sp4_v_b_28')
// (14, 10, 'sp4_r_v_b_16')
// (14, 10, 'sp4_v_b_17')
// (14, 11, 'sp4_r_v_b_5')
// (14, 11, 'sp4_v_b_4')
// (15, 3, 'sp4_v_t_44')
// (15, 4, 'neigh_op_tnl_0')
// (15, 4, 'sp4_v_b_44')
// (15, 5, 'neigh_op_lft_0')
// (15, 5, 'sp4_v_b_33')
// (15, 6, 'neigh_op_bnl_0')
// (15, 6, 'sp4_v_b_20')
// (15, 7, 'local_g1_5')
// (15, 7, 'lutff_3/in_1')
// (15, 7, 'sp4_h_r_21')
// (15, 7, 'sp4_v_b_9')
// (15, 7, 'sp4_v_t_40')
// (15, 8, 'sp4_v_b_40')
// (15, 9, 'local_g2_5')
// (15, 9, 'lutff_0/in_1')
// (15, 9, 'sp4_v_b_29')
// (15, 10, 'sp4_v_b_16')
// (15, 11, 'sp4_v_b_5')
// (16, 7, 'sp4_h_r_32')
// (17, 7, 'sp4_h_r_45')
// (18, 7, 'sp4_h_l_45')

wire n1886;
// (13, 4, 'neigh_op_tnr_1')
// (13, 5, 'local_g2_1')
// (13, 5, 'lutff_3/in_2')
// (13, 5, 'neigh_op_rgt_1')
// (13, 6, 'neigh_op_bnr_1')
// (14, 4, 'neigh_op_top_1')
// (14, 5, 'lutff_1/out')
// (14, 6, 'neigh_op_bot_1')
// (15, 4, 'neigh_op_tnl_1')
// (15, 5, 'neigh_op_lft_1')
// (15, 6, 'neigh_op_bnl_1')

reg n1887 = 0;
// (13, 4, 'neigh_op_tnr_3')
// (13, 5, 'local_g3_3')
// (13, 5, 'lutff_2/in_2')
// (13, 5, 'neigh_op_rgt_3')
// (13, 5, 'sp4_r_v_b_38')
// (13, 6, 'neigh_op_bnr_3')
// (13, 6, 'sp4_r_v_b_27')
// (13, 7, 'local_g2_6')
// (13, 7, 'lutff_0/in_2')
// (13, 7, 'sp4_r_v_b_14')
// (13, 8, 'local_g1_3')
// (13, 8, 'lutff_6/in_0')
// (13, 8, 'sp4_r_v_b_3')
// (14, 4, 'neigh_op_top_3')
// (14, 4, 'sp4_v_t_38')
// (14, 5, 'lutff_3/out')
// (14, 5, 'sp4_v_b_38')
// (14, 6, 'neigh_op_bot_3')
// (14, 6, 'sp4_v_b_27')
// (14, 7, 'sp4_v_b_14')
// (14, 8, 'sp4_h_r_9')
// (14, 8, 'sp4_v_b_3')
// (15, 4, 'neigh_op_tnl_3')
// (15, 5, 'neigh_op_lft_3')
// (15, 6, 'local_g3_3')
// (15, 6, 'lutff_6/in_0')
// (15, 6, 'neigh_op_bnl_3')
// (15, 8, 'local_g0_4')
// (15, 8, 'lutff_7/in_1')
// (15, 8, 'sp4_h_r_20')
// (16, 8, 'sp4_h_r_33')
// (17, 8, 'sp4_h_r_44')
// (18, 8, 'sp4_h_l_44')

reg n1888 = 0;
// (13, 4, 'neigh_op_tnr_6')
// (13, 5, 'neigh_op_rgt_6')
// (13, 6, 'neigh_op_bnr_6')
// (14, 0, 'span12_vert_20')
// (14, 1, 'sp12_v_b_20')
// (14, 2, 'sp12_v_b_19')
// (14, 3, 'sp12_v_b_16')
// (14, 4, 'neigh_op_top_6')
// (14, 4, 'sp12_v_b_15')
// (14, 5, 'local_g3_6')
// (14, 5, 'lutff_1/in_2')
// (14, 5, 'lutff_6/out')
// (14, 5, 'sp12_v_b_12')
// (14, 5, 'sp4_r_v_b_45')
// (14, 6, 'neigh_op_bot_6')
// (14, 6, 'sp12_v_b_11')
// (14, 6, 'sp4_r_v_b_32')
// (14, 7, 'sp12_v_b_8')
// (14, 7, 'sp4_r_v_b_21')
// (14, 8, 'local_g2_0')
// (14, 8, 'lutff_2/in_2')
// (14, 8, 'sp12_v_b_7')
// (14, 8, 'sp4_r_v_b_8')
// (14, 9, 'sp12_v_b_4')
// (14, 9, 'sp4_r_v_b_45')
// (14, 10, 'local_g2_3')
// (14, 10, 'lutff_5/in_0')
// (14, 10, 'sp12_v_b_3')
// (14, 10, 'sp4_r_v_b_32')
// (14, 11, 'sp12_v_b_0')
// (14, 11, 'sp4_r_v_b_21')
// (14, 12, 'sp4_r_v_b_8')
// (15, 4, 'neigh_op_tnl_6')
// (15, 4, 'sp4_v_t_45')
// (15, 5, 'neigh_op_lft_6')
// (15, 5, 'sp4_v_b_45')
// (15, 6, 'local_g2_6')
// (15, 6, 'lutff_2/in_2')
// (15, 6, 'neigh_op_bnl_6')
// (15, 6, 'sp4_v_b_32')
// (15, 7, 'sp4_v_b_21')
// (15, 8, 'sp4_v_b_8')
// (15, 8, 'sp4_v_t_45')
// (15, 9, 'sp4_v_b_45')
// (15, 10, 'local_g2_0')
// (15, 10, 'lutff_1/in_3')
// (15, 10, 'sp4_v_b_32')
// (15, 11, 'sp4_v_b_21')
// (15, 12, 'sp4_v_b_8')

reg n1889 = 0;
// (13, 4, 'neigh_op_tnr_7')
// (13, 5, 'neigh_op_rgt_7')
// (13, 6, 'neigh_op_bnr_7')
// (14, 4, 'neigh_op_top_7')
// (14, 5, 'lutff_7/out')
// (14, 5, 'sp4_r_v_b_47')
// (14, 6, 'neigh_op_bot_7')
// (14, 6, 'sp4_r_v_b_34')
// (14, 7, 'local_g3_7')
// (14, 7, 'lutff_2/in_2')
// (14, 7, 'lutff_5/in_1')
// (14, 7, 'sp4_r_v_b_23')
// (14, 8, 'local_g2_2')
// (14, 8, 'lutff_3/in_3')
// (14, 8, 'sp4_r_v_b_10')
// (15, 4, 'neigh_op_tnl_7')
// (15, 4, 'sp4_v_t_47')
// (15, 5, 'neigh_op_lft_7')
// (15, 5, 'sp4_v_b_47')
// (15, 6, 'local_g3_7')
// (15, 6, 'lutff_1/in_1')
// (15, 6, 'neigh_op_bnl_7')
// (15, 6, 'sp4_v_b_34')
// (15, 7, 'sp4_v_b_23')
// (15, 8, 'local_g1_2')
// (15, 8, 'lutff_0/in_3')
// (15, 8, 'sp4_v_b_10')

reg n1890 = 0;
// (13, 4, 'sp4_r_v_b_38')
// (13, 5, 'sp4_r_v_b_27')
// (13, 6, 'sp4_r_v_b_14')
// (13, 7, 'sp4_r_v_b_3')
// (13, 8, 'sp4_r_v_b_46')
// (13, 9, 'local_g2_3')
// (13, 9, 'lutff_1/in_2')
// (13, 9, 'sp4_r_v_b_35')
// (13, 10, 'sp4_r_v_b_22')
// (13, 11, 'sp4_r_v_b_11')
// (14, 2, 'neigh_op_tnr_2')
// (14, 3, 'neigh_op_rgt_2')
// (14, 3, 'sp4_h_r_9')
// (14, 3, 'sp4_v_t_38')
// (14, 4, 'neigh_op_bnr_2')
// (14, 4, 'sp4_v_b_38')
// (14, 5, 'sp4_v_b_27')
// (14, 6, 'sp4_v_b_14')
// (14, 7, 'sp4_v_b_3')
// (14, 7, 'sp4_v_t_46')
// (14, 8, 'sp4_v_b_46')
// (14, 9, 'sp4_v_b_35')
// (14, 10, 'sp4_v_b_22')
// (14, 11, 'sp4_v_b_11')
// (15, 1, 'sp12_v_t_23')
// (15, 2, 'local_g0_2')
// (15, 2, 'lutff_3/in_1')
// (15, 2, 'neigh_op_top_2')
// (15, 2, 'sp12_v_b_23')
// (15, 3, 'lutff_2/out')
// (15, 3, 'sp12_v_b_20')
// (15, 3, 'sp4_h_r_20')
// (15, 3, 'sp4_r_v_b_37')
// (15, 4, 'neigh_op_bot_2')
// (15, 4, 'sp12_v_b_19')
// (15, 4, 'sp4_r_v_b_24')
// (15, 5, 'sp12_v_b_16')
// (15, 5, 'sp4_r_v_b_13')
// (15, 6, 'sp12_v_b_15')
// (15, 6, 'sp4_r_v_b_0')
// (15, 7, 'sp12_v_b_12')
// (15, 8, 'sp12_v_b_11')
// (15, 9, 'local_g3_0')
// (15, 9, 'lutff_5/in_0')
// (15, 9, 'sp12_v_b_8')
// (15, 10, 'sp12_v_b_7')
// (15, 11, 'sp12_v_b_4')
// (15, 12, 'sp12_v_b_3')
// (15, 13, 'sp12_v_b_0')
// (16, 2, 'neigh_op_tnl_2')
// (16, 2, 'sp4_v_t_37')
// (16, 3, 'neigh_op_lft_2')
// (16, 3, 'sp4_h_r_33')
// (16, 3, 'sp4_v_b_37')
// (16, 4, 'neigh_op_bnl_2')
// (16, 4, 'sp4_v_b_24')
// (16, 5, 'sp4_v_b_13')
// (16, 6, 'local_g0_0')
// (16, 6, 'lutff_2/in_0')
// (16, 6, 'lutff_6/in_2')
// (16, 6, 'sp4_v_b_0')
// (17, 3, 'sp4_h_r_44')
// (18, 3, 'sp4_h_l_44')

reg n1891 = 0;
// (13, 4, 'sp4_r_v_b_39')
// (13, 5, 'sp4_r_v_b_26')
// (13, 6, 'local_g2_7')
// (13, 6, 'lutff_1/in_2')
// (13, 6, 'lutff_5/in_0')
// (13, 6, 'sp4_r_v_b_15')
// (13, 7, 'sp4_r_v_b_2')
// (13, 8, 'sp4_r_v_b_43')
// (13, 9, 'sp4_r_v_b_30')
// (13, 10, 'neigh_op_tnr_3')
// (13, 10, 'sp4_r_v_b_19')
// (13, 11, 'local_g2_3')
// (13, 11, 'lutff_5/in_2')
// (13, 11, 'neigh_op_rgt_3')
// (13, 11, 'sp4_h_r_11')
// (13, 11, 'sp4_r_v_b_6')
// (13, 12, 'neigh_op_bnr_3')
// (14, 3, 'sp4_v_t_39')
// (14, 4, 'sp4_v_b_39')
// (14, 5, 'sp4_v_b_26')
// (14, 6, 'sp4_v_b_15')
// (14, 7, 'sp4_v_b_2')
// (14, 7, 'sp4_v_t_43')
// (14, 8, 'sp4_v_b_43')
// (14, 9, 'sp4_r_v_b_47')
// (14, 9, 'sp4_v_b_30')
// (14, 10, 'neigh_op_top_3')
// (14, 10, 'sp4_r_v_b_34')
// (14, 10, 'sp4_v_b_19')
// (14, 11, 'lutff_3/out')
// (14, 11, 'sp4_h_r_22')
// (14, 11, 'sp4_r_v_b_23')
// (14, 11, 'sp4_v_b_6')
// (14, 12, 'neigh_op_bot_3')
// (14, 12, 'sp4_r_v_b_10')
// (15, 8, 'sp4_v_t_47')
// (15, 9, 'sp4_v_b_47')
// (15, 10, 'neigh_op_tnl_3')
// (15, 10, 'sp4_v_b_34')
// (15, 11, 'neigh_op_lft_3')
// (15, 11, 'sp4_h_r_35')
// (15, 11, 'sp4_v_b_23')
// (15, 12, 'local_g3_3')
// (15, 12, 'lutff_2/in_2')
// (15, 12, 'neigh_op_bnl_3')
// (15, 12, 'sp4_h_r_10')
// (15, 12, 'sp4_v_b_10')
// (16, 4, 'sp4_r_v_b_45')
// (16, 5, 'sp4_r_v_b_32')
// (16, 6, 'local_g3_5')
// (16, 6, 'lutff_0/in_2')
// (16, 6, 'sp4_r_v_b_21')
// (16, 7, 'sp4_r_v_b_8')
// (16, 8, 'sp4_r_v_b_40')
// (16, 9, 'sp4_r_v_b_29')
// (16, 10, 'sp4_r_v_b_16')
// (16, 11, 'sp4_h_r_46')
// (16, 11, 'sp4_r_v_b_5')
// (16, 12, 'local_g1_7')
// (16, 12, 'lutff_3/in_3')
// (16, 12, 'sp4_h_r_23')
// (17, 3, 'sp4_v_t_45')
// (17, 4, 'sp4_v_b_45')
// (17, 5, 'sp4_v_b_32')
// (17, 6, 'sp4_v_b_21')
// (17, 7, 'sp4_v_b_8')
// (17, 7, 'sp4_v_t_40')
// (17, 8, 'sp4_v_b_40')
// (17, 9, 'sp4_v_b_29')
// (17, 10, 'sp4_v_b_16')
// (17, 11, 'sp4_h_l_46')
// (17, 11, 'sp4_v_b_5')
// (17, 12, 'sp4_h_r_34')
// (18, 12, 'sp4_h_r_47')
// (19, 12, 'sp4_h_l_47')

reg n1892 = 0;
// (13, 4, 'sp4_r_v_b_42')
// (13, 5, 'sp4_r_v_b_31')
// (13, 6, 'local_g3_2')
// (13, 6, 'lutff_2/in_1')
// (13, 6, 'sp4_r_v_b_18')
// (13, 7, 'sp4_r_v_b_7')
// (13, 8, 'sp4_r_v_b_42')
// (13, 9, 'neigh_op_tnr_1')
// (13, 9, 'sp4_r_v_b_31')
// (13, 10, 'neigh_op_rgt_1')
// (13, 10, 'sp4_h_r_7')
// (13, 10, 'sp4_r_v_b_18')
// (13, 11, 'neigh_op_bnr_1')
// (13, 11, 'sp4_r_v_b_7')
// (14, 3, 'sp4_r_v_b_38')
// (14, 3, 'sp4_v_t_42')
// (14, 4, 'sp4_r_v_b_27')
// (14, 4, 'sp4_v_b_42')
// (14, 5, 'sp4_r_v_b_14')
// (14, 5, 'sp4_v_b_31')
// (14, 6, 'sp4_r_v_b_3')
// (14, 6, 'sp4_v_b_18')
// (14, 7, 'sp4_r_v_b_38')
// (14, 7, 'sp4_v_b_7')
// (14, 7, 'sp4_v_t_42')
// (14, 8, 'sp4_r_v_b_27')
// (14, 8, 'sp4_r_v_b_43')
// (14, 8, 'sp4_v_b_42')
// (14, 9, 'neigh_op_top_1')
// (14, 9, 'sp4_r_v_b_14')
// (14, 9, 'sp4_r_v_b_30')
// (14, 9, 'sp4_v_b_31')
// (14, 10, 'lutff_1/out')
// (14, 10, 'sp4_h_r_18')
// (14, 10, 'sp4_r_v_b_19')
// (14, 10, 'sp4_r_v_b_3')
// (14, 10, 'sp4_v_b_18')
// (14, 11, 'local_g1_1')
// (14, 11, 'lutff_3/in_1')
// (14, 11, 'neigh_op_bot_1')
// (14, 11, 'sp4_r_v_b_6')
// (14, 11, 'sp4_v_b_7')
// (14, 12, 'sp4_r_v_b_44')
// (14, 13, 'sp4_r_v_b_33')
// (14, 14, 'sp4_r_v_b_20')
// (14, 15, 'sp4_r_v_b_9')
// (15, 2, 'sp4_v_t_38')
// (15, 3, 'sp4_v_b_38')
// (15, 4, 'sp4_v_b_27')
// (15, 5, 'local_g0_6')
// (15, 5, 'lutff_2/in_0')
// (15, 5, 'sp4_v_b_14')
// (15, 6, 'sp4_v_b_3')
// (15, 6, 'sp4_v_t_38')
// (15, 7, 'sp4_v_b_38')
// (15, 7, 'sp4_v_t_43')
// (15, 8, 'sp4_v_b_27')
// (15, 8, 'sp4_v_b_43')
// (15, 9, 'neigh_op_tnl_1')
// (15, 9, 'sp4_v_b_14')
// (15, 9, 'sp4_v_b_30')
// (15, 10, 'neigh_op_lft_1')
// (15, 10, 'sp4_h_r_31')
// (15, 10, 'sp4_v_b_19')
// (15, 10, 'sp4_v_b_3')
// (15, 11, 'local_g3_1')
// (15, 11, 'lutff_1/in_3')
// (15, 11, 'neigh_op_bnl_1')
// (15, 11, 'sp4_v_b_6')
// (15, 11, 'sp4_v_t_44')
// (15, 12, 'sp4_v_b_44')
// (15, 13, 'local_g2_1')
// (15, 13, 'lutff_0/in_1')
// (15, 13, 'sp4_v_b_33')
// (15, 14, 'sp4_v_b_20')
// (15, 15, 'sp4_v_b_9')
// (16, 3, 'sp4_r_v_b_47')
// (16, 4, 'sp4_r_v_b_34')
// (16, 5, 'local_g3_7')
// (16, 5, 'lutff_7/in_1')
// (16, 5, 'sp4_r_v_b_23')
// (16, 6, 'sp4_r_v_b_10')
// (16, 7, 'sp4_r_v_b_42')
// (16, 8, 'sp4_r_v_b_31')
// (16, 9, 'sp4_r_v_b_18')
// (16, 10, 'sp4_h_r_42')
// (16, 10, 'sp4_r_v_b_7')
// (17, 2, 'sp4_v_t_47')
// (17, 3, 'sp4_v_b_47')
// (17, 4, 'sp4_v_b_34')
// (17, 5, 'sp4_v_b_23')
// (17, 6, 'sp4_v_b_10')
// (17, 6, 'sp4_v_t_42')
// (17, 7, 'sp4_v_b_42')
// (17, 8, 'sp4_v_b_31')
// (17, 9, 'sp4_v_b_18')
// (17, 10, 'sp4_h_l_42')
// (17, 10, 'sp4_v_b_7')

reg n1893 = 0;
// (13, 5, 'local_g1_0')
// (13, 5, 'lutff_6/in_3')
// (13, 5, 'sp4_h_r_8')
// (14, 4, 'neigh_op_tnr_0')
// (14, 5, 'neigh_op_rgt_0')
// (14, 5, 'sp4_h_r_21')
// (14, 6, 'local_g1_0')
// (14, 6, 'lutff_0/in_3')
// (14, 6, 'lutff_6/in_1')
// (14, 6, 'neigh_op_bnr_0')
// (15, 4, 'neigh_op_top_0')
// (15, 4, 'sp4_r_v_b_44')
// (15, 5, 'lutff_0/out')
// (15, 5, 'sp4_h_r_32')
// (15, 5, 'sp4_r_v_b_33')
// (15, 6, 'neigh_op_bot_0')
// (15, 6, 'sp4_r_v_b_20')
// (15, 7, 'sp4_r_v_b_9')
// (16, 3, 'sp4_v_t_44')
// (16, 4, 'neigh_op_tnl_0')
// (16, 4, 'sp4_v_b_44')
// (16, 5, 'neigh_op_lft_0')
// (16, 5, 'sp4_h_r_45')
// (16, 5, 'sp4_v_b_33')
// (16, 6, 'local_g3_0')
// (16, 6, 'lutff_7/in_2')
// (16, 6, 'neigh_op_bnl_0')
// (16, 6, 'sp4_v_b_20')
// (16, 7, 'local_g0_1')
// (16, 7, 'lutff_4/in_1')
// (16, 7, 'sp4_v_b_9')
// (17, 5, 'sp4_h_l_45')

wire n1894;
// (13, 5, 'neigh_op_tnr_0')
// (13, 6, 'neigh_op_rgt_0')
// (13, 7, 'neigh_op_bnr_0')
// (14, 5, 'neigh_op_top_0')
// (14, 6, 'local_g3_0')
// (14, 6, 'lutff_0/out')
// (14, 6, 'lutff_5/in_2')
// (14, 7, 'neigh_op_bot_0')
// (15, 5, 'neigh_op_tnl_0')
// (15, 6, 'neigh_op_lft_0')
// (15, 7, 'neigh_op_bnl_0')

wire n1895;
// (13, 5, 'neigh_op_tnr_1')
// (13, 6, 'neigh_op_rgt_1')
// (13, 7, 'neigh_op_bnr_1')
// (14, 5, 'neigh_op_top_1')
// (14, 6, 'local_g3_1')
// (14, 6, 'lutff_1/out')
// (14, 6, 'lutff_5/in_3')
// (14, 7, 'neigh_op_bot_1')
// (15, 5, 'neigh_op_tnl_1')
// (15, 6, 'neigh_op_lft_1')
// (15, 7, 'neigh_op_bnl_1')

wire n1896;
// (13, 5, 'neigh_op_tnr_2')
// (13, 6, 'neigh_op_rgt_2')
// (13, 7, 'local_g0_2')
// (13, 7, 'lutff_3/in_3')
// (13, 7, 'neigh_op_bnr_2')
// (14, 5, 'neigh_op_top_2')
// (14, 6, 'lutff_2/out')
// (14, 7, 'neigh_op_bot_2')
// (15, 5, 'neigh_op_tnl_2')
// (15, 6, 'neigh_op_lft_2')
// (15, 7, 'neigh_op_bnl_2')

wire n1897;
// (13, 5, 'neigh_op_tnr_3')
// (13, 6, 'neigh_op_rgt_3')
// (13, 7, 'neigh_op_bnr_3')
// (14, 5, 'neigh_op_top_3')
// (14, 6, 'local_g3_3')
// (14, 6, 'lutff_3/out')
// (14, 6, 'lutff_5/in_1')
// (14, 7, 'neigh_op_bot_3')
// (15, 5, 'neigh_op_tnl_3')
// (15, 6, 'neigh_op_lft_3')
// (15, 7, 'neigh_op_bnl_3')

wire n1898;
// (13, 5, 'neigh_op_tnr_4')
// (13, 6, 'neigh_op_rgt_4')
// (13, 7, 'neigh_op_bnr_4')
// (14, 5, 'neigh_op_top_4')
// (14, 6, 'local_g3_4')
// (14, 6, 'lutff_4/out')
// (14, 6, 'lutff_5/in_0')
// (14, 7, 'neigh_op_bot_4')
// (15, 5, 'neigh_op_tnl_4')
// (15, 6, 'neigh_op_lft_4')
// (15, 7, 'neigh_op_bnl_4')

wire n1899;
// (13, 5, 'neigh_op_tnr_5')
// (13, 6, 'neigh_op_rgt_5')
// (13, 6, 'sp4_r_v_b_42')
// (13, 7, 'neigh_op_bnr_5')
// (13, 7, 'sp4_r_v_b_31')
// (13, 8, 'sp4_r_v_b_18')
// (13, 9, 'sp4_r_v_b_7')
// (14, 5, 'neigh_op_top_5')
// (14, 5, 'sp4_v_t_42')
// (14, 6, 'lutff_5/out')
// (14, 6, 'sp4_v_b_42')
// (14, 7, 'neigh_op_bot_5')
// (14, 7, 'sp4_v_b_31')
// (14, 8, 'local_g0_2')
// (14, 8, 'lutff_0/in_0')
// (14, 8, 'sp4_v_b_18')
// (14, 9, 'sp4_v_b_7')
// (15, 5, 'neigh_op_tnl_5')
// (15, 6, 'neigh_op_lft_5')
// (15, 7, 'neigh_op_bnl_5')

wire n1900;
// (13, 5, 'neigh_op_tnr_6')
// (13, 6, 'neigh_op_rgt_6')
// (13, 7, 'neigh_op_bnr_6')
// (14, 5, 'neigh_op_top_6')
// (14, 6, 'lutff_6/out')
// (14, 7, 'local_g1_6')
// (14, 7, 'lutff_6/in_3')
// (14, 7, 'neigh_op_bot_6')
// (15, 5, 'neigh_op_tnl_6')
// (15, 6, 'neigh_op_lft_6')
// (15, 7, 'neigh_op_bnl_6')

reg n1901 = 0;
// (13, 5, 'neigh_op_tnr_7')
// (13, 6, 'neigh_op_rgt_7')
// (13, 7, 'neigh_op_bnr_7')
// (14, 5, 'local_g1_7')
// (14, 5, 'lutff_1/in_1')
// (14, 5, 'neigh_op_top_7')
// (14, 6, 'local_g3_7')
// (14, 6, 'lutff_2/in_2')
// (14, 6, 'lutff_7/out')
// (14, 7, 'neigh_op_bot_7')
// (15, 5, 'neigh_op_tnl_7')
// (15, 6, 'local_g1_7')
// (15, 6, 'lutff_7/in_3')
// (15, 6, 'neigh_op_lft_7')
// (15, 7, 'neigh_op_bnl_7')

wire n1902;
// (13, 5, 'sp4_h_r_10')
// (14, 4, 'neigh_op_tnr_1')
// (14, 5, 'neigh_op_rgt_1')
// (14, 5, 'sp4_h_r_23')
// (14, 6, 'neigh_op_bnr_1')
// (15, 4, 'neigh_op_top_1')
// (15, 5, 'lutff_1/out')
// (15, 5, 'sp4_h_r_34')
// (15, 6, 'neigh_op_bot_1')
// (16, 4, 'neigh_op_tnl_1')
// (16, 5, 'local_g2_7')
// (16, 5, 'lutff_1/in_0')
// (16, 5, 'neigh_op_lft_1')
// (16, 5, 'sp4_h_r_47')
// (16, 6, 'neigh_op_bnl_1')
// (17, 5, 'sp4_h_l_47')

reg n1903 = 0;
// (13, 5, 'sp4_r_v_b_40')
// (13, 5, 'sp4_r_v_b_46')
// (13, 6, 'sp4_r_v_b_29')
// (13, 6, 'sp4_r_v_b_35')
// (13, 7, 'sp4_r_v_b_16')
// (13, 7, 'sp4_r_v_b_22')
// (13, 8, 'sp4_r_v_b_11')
// (13, 8, 'sp4_r_v_b_5')
// (14, 2, 'sp4_r_v_b_46')
// (14, 3, 'neigh_op_tnr_3')
// (14, 3, 'sp4_r_v_b_35')
// (14, 4, 'neigh_op_rgt_3')
// (14, 4, 'sp4_h_r_11')
// (14, 4, 'sp4_r_v_b_22')
// (14, 4, 'sp4_v_t_40')
// (14, 4, 'sp4_v_t_46')
// (14, 5, 'neigh_op_bnr_3')
// (14, 5, 'sp4_r_v_b_11')
// (14, 5, 'sp4_v_b_40')
// (14, 5, 'sp4_v_b_46')
// (14, 6, 'sp4_r_v_b_39')
// (14, 6, 'sp4_v_b_29')
// (14, 6, 'sp4_v_b_35')
// (14, 7, 'local_g0_6')
// (14, 7, 'lutff_2/in_0')
// (14, 7, 'sp4_r_v_b_26')
// (14, 7, 'sp4_v_b_16')
// (14, 7, 'sp4_v_b_22')
// (14, 8, 'local_g0_5')
// (14, 8, 'lutff_3/in_0')
// (14, 8, 'sp4_r_v_b_15')
// (14, 8, 'sp4_v_b_11')
// (14, 8, 'sp4_v_b_5')
// (14, 9, 'sp4_r_v_b_2')
// (15, 1, 'sp4_v_t_46')
// (15, 2, 'sp4_v_b_46')
// (15, 3, 'neigh_op_top_3')
// (15, 3, 'sp4_v_b_35')
// (15, 4, 'local_g1_3')
// (15, 4, 'lutff_3/out')
// (15, 4, 'lutff_5/in_3')
// (15, 4, 'sp4_h_r_22')
// (15, 4, 'sp4_r_v_b_39')
// (15, 4, 'sp4_v_b_22')
// (15, 5, 'neigh_op_bot_3')
// (15, 5, 'sp4_r_v_b_26')
// (15, 5, 'sp4_v_b_11')
// (15, 5, 'sp4_v_t_39')
// (15, 6, 'local_g2_7')
// (15, 6, 'lutff_1/in_2')
// (15, 6, 'sp4_r_v_b_15')
// (15, 6, 'sp4_v_b_39')
// (15, 7, 'sp4_r_v_b_2')
// (15, 7, 'sp4_v_b_26')
// (15, 8, 'local_g1_7')
// (15, 8, 'lutff_0/in_0')
// (15, 8, 'sp4_v_b_15')
// (15, 9, 'sp4_v_b_2')
// (16, 3, 'neigh_op_tnl_3')
// (16, 3, 'sp4_v_t_39')
// (16, 4, 'neigh_op_lft_3')
// (16, 4, 'sp4_h_r_35')
// (16, 4, 'sp4_v_b_39')
// (16, 5, 'neigh_op_bnl_3')
// (16, 5, 'sp4_v_b_26')
// (16, 6, 'sp4_v_b_15')
// (16, 7, 'sp4_v_b_2')
// (17, 4, 'sp4_h_r_46')
// (18, 4, 'sp4_h_l_46')

reg n1904 = 0;
// (13, 5, 'sp4_r_v_b_42')
// (13, 6, 'sp4_r_v_b_31')
// (13, 7, 'sp4_r_v_b_18')
// (13, 8, 'sp4_r_v_b_7')
// (14, 3, 'neigh_op_tnr_1')
// (14, 4, 'local_g3_1')
// (14, 4, 'lutff_7/in_1')
// (14, 4, 'neigh_op_rgt_1')
// (14, 4, 'sp4_h_r_7')
// (14, 4, 'sp4_v_t_42')
// (14, 5, 'neigh_op_bnr_1')
// (14, 5, 'sp4_v_b_42')
// (14, 6, 'sp4_v_b_31')
// (14, 7, 'local_g0_2')
// (14, 7, 'lutff_0/in_0')
// (14, 7, 'lutff_1/in_1')
// (14, 7, 'sp4_v_b_18')
// (14, 8, 'sp4_v_b_7')
// (15, 1, 'sp4_r_v_b_38')
// (15, 2, 'sp4_r_v_b_27')
// (15, 3, 'neigh_op_top_1')
// (15, 3, 'sp4_r_v_b_14')
// (15, 4, 'lutff_1/out')
// (15, 4, 'sp4_h_r_18')
// (15, 4, 'sp4_r_v_b_3')
// (15, 5, 'neigh_op_bot_1')
// (15, 5, 'sp4_r_v_b_43')
// (15, 5, 'sp4_r_v_b_46')
// (15, 6, 'sp4_r_v_b_30')
// (15, 6, 'sp4_r_v_b_35')
// (15, 7, 'local_g3_6')
// (15, 7, 'lutff_6/in_1')
// (15, 7, 'sp4_r_v_b_19')
// (15, 7, 'sp4_r_v_b_22')
// (15, 8, 'sp4_r_v_b_11')
// (15, 8, 'sp4_r_v_b_6')
// (16, 0, 'span4_vert_38')
// (16, 1, 'sp4_v_b_38')
// (16, 2, 'sp4_v_b_27')
// (16, 3, 'neigh_op_tnl_1')
// (16, 3, 'sp4_v_b_14')
// (16, 4, 'neigh_op_lft_1')
// (16, 4, 'sp4_h_r_31')
// (16, 4, 'sp4_v_b_3')
// (16, 4, 'sp4_v_t_43')
// (16, 4, 'sp4_v_t_46')
// (16, 5, 'neigh_op_bnl_1')
// (16, 5, 'sp4_v_b_43')
// (16, 5, 'sp4_v_b_46')
// (16, 6, 'sp4_v_b_30')
// (16, 6, 'sp4_v_b_35')
// (16, 7, 'local_g1_3')
// (16, 7, 'lutff_7/in_1')
// (16, 7, 'sp4_v_b_19')
// (16, 7, 'sp4_v_b_22')
// (16, 8, 'sp4_v_b_11')
// (16, 8, 'sp4_v_b_6')
// (17, 4, 'sp4_h_r_42')
// (18, 4, 'sp4_h_l_42')

wire n1905;
// (13, 6, 'neigh_op_tnr_0')
// (13, 7, 'neigh_op_rgt_0')
// (13, 8, 'neigh_op_bnr_0')
// (14, 6, 'neigh_op_top_0')
// (14, 7, 'local_g0_0')
// (14, 7, 'lutff_0/out')
// (14, 7, 'lutff_6/in_0')
// (14, 8, 'neigh_op_bot_0')
// (15, 6, 'neigh_op_tnl_0')
// (15, 7, 'neigh_op_lft_0')
// (15, 8, 'neigh_op_bnl_0')

wire n1906;
// (13, 6, 'neigh_op_tnr_1')
// (13, 7, 'neigh_op_rgt_1')
// (13, 8, 'neigh_op_bnr_1')
// (14, 6, 'neigh_op_top_1')
// (14, 7, 'lutff_1/out')
// (14, 8, 'local_g1_1')
// (14, 8, 'lutff_4/in_2')
// (14, 8, 'neigh_op_bot_1')
// (15, 6, 'neigh_op_tnl_1')
// (15, 7, 'neigh_op_lft_1')
// (15, 8, 'neigh_op_bnl_1')

wire n1907;
// (13, 6, 'neigh_op_tnr_2')
// (13, 7, 'neigh_op_rgt_2')
// (13, 8, 'neigh_op_bnr_2')
// (14, 6, 'neigh_op_top_2')
// (14, 7, 'local_g3_2')
// (14, 7, 'lutff_2/out')
// (14, 7, 'lutff_6/in_1')
// (14, 8, 'neigh_op_bot_2')
// (15, 6, 'neigh_op_tnl_2')
// (15, 7, 'neigh_op_lft_2')
// (15, 8, 'neigh_op_bnl_2')

wire n1908;
// (13, 6, 'neigh_op_tnr_3')
// (13, 7, 'local_g3_3')
// (13, 7, 'lutff_3/in_1')
// (13, 7, 'neigh_op_rgt_3')
// (13, 8, 'neigh_op_bnr_3')
// (14, 6, 'neigh_op_top_3')
// (14, 7, 'lutff_3/out')
// (14, 8, 'neigh_op_bot_3')
// (15, 6, 'neigh_op_tnl_3')
// (15, 7, 'neigh_op_lft_3')
// (15, 8, 'neigh_op_bnl_3')

reg n1909 = 0;
// (13, 6, 'neigh_op_tnr_4')
// (13, 7, 'neigh_op_rgt_4')
// (13, 8, 'neigh_op_bnr_4')
// (14, 6, 'neigh_op_top_4')
// (14, 7, 'local_g2_4')
// (14, 7, 'lutff_4/out')
// (14, 7, 'lutff_5/in_3')
// (14, 8, 'local_g0_4')
// (14, 8, 'lutff_6/in_2')
// (14, 8, 'neigh_op_bot_4')
// (15, 6, 'neigh_op_tnl_4')
// (15, 7, 'neigh_op_lft_4')
// (15, 8, 'local_g2_4')
// (15, 8, 'lutff_5/in_3')
// (15, 8, 'neigh_op_bnl_4')

wire n1910;
// (13, 6, 'neigh_op_tnr_5')
// (13, 7, 'local_g3_5')
// (13, 7, 'lutff_1/in_3')
// (13, 7, 'neigh_op_rgt_5')
// (13, 8, 'neigh_op_bnr_5')
// (14, 6, 'neigh_op_top_5')
// (14, 7, 'lutff_5/out')
// (14, 8, 'neigh_op_bot_5')
// (15, 6, 'neigh_op_tnl_5')
// (15, 7, 'neigh_op_lft_5')
// (15, 8, 'neigh_op_bnl_5')

wire n1911;
// (13, 6, 'neigh_op_tnr_6')
// (13, 7, 'neigh_op_rgt_6')
// (13, 8, 'neigh_op_bnr_6')
// (14, 6, 'neigh_op_top_6')
// (14, 7, 'local_g2_6')
// (14, 7, 'lutff_6/out')
// (14, 7, 'lutff_7/in_3')
// (14, 8, 'neigh_op_bot_6')
// (15, 6, 'neigh_op_tnl_6')
// (15, 7, 'neigh_op_lft_6')
// (15, 8, 'neigh_op_bnl_6')

wire n1912;
// (13, 6, 'neigh_op_tnr_7')
// (13, 7, 'local_g3_7')
// (13, 7, 'lutff_6/in_2')
// (13, 7, 'neigh_op_rgt_7')
// (13, 8, 'neigh_op_bnr_7')
// (14, 6, 'neigh_op_top_7')
// (14, 7, 'lutff_7/out')
// (14, 8, 'neigh_op_bot_7')
// (15, 6, 'neigh_op_tnl_7')
// (15, 7, 'neigh_op_lft_7')
// (15, 8, 'neigh_op_bnl_7')

wire n1913;
// (13, 6, 'sp4_r_v_b_37')
// (13, 7, 'sp4_r_v_b_24')
// (13, 8, 'neigh_op_tnr_0')
// (13, 8, 'sp4_r_v_b_13')
// (13, 9, 'neigh_op_rgt_0')
// (13, 9, 'sp4_r_v_b_0')
// (13, 10, 'neigh_op_bnr_0')
// (14, 5, 'sp4_v_t_37')
// (14, 6, 'sp4_v_b_37')
// (14, 7, 'local_g2_0')
// (14, 7, 'lutff_6/in_2')
// (14, 7, 'sp4_v_b_24')
// (14, 8, 'neigh_op_top_0')
// (14, 8, 'sp4_v_b_13')
// (14, 9, 'lutff_0/out')
// (14, 9, 'sp4_v_b_0')
// (14, 10, 'neigh_op_bot_0')
// (15, 8, 'neigh_op_tnl_0')
// (15, 9, 'neigh_op_lft_0')
// (15, 10, 'neigh_op_bnl_0')

reg n1914 = 0;
// (13, 6, 'sp4_r_v_b_45')
// (13, 7, 'sp4_r_v_b_32')
// (13, 8, 'sp4_r_v_b_21')
// (13, 9, 'sp4_r_v_b_8')
// (14, 5, 'local_g1_0')
// (14, 5, 'lutff_4/in_3')
// (14, 5, 'sp4_h_r_8')
// (14, 5, 'sp4_v_t_45')
// (14, 6, 'sp4_v_b_45')
// (14, 7, 'sp4_v_b_32')
// (14, 8, 'local_g1_5')
// (14, 8, 'lutff_1/in_1')
// (14, 8, 'sp4_v_b_21')
// (14, 9, 'sp4_v_b_8')
// (15, 2, 'sp4_r_v_b_37')
// (15, 3, 'sp4_r_v_b_24')
// (15, 4, 'neigh_op_tnr_0')
// (15, 4, 'sp4_r_v_b_13')
// (15, 5, 'neigh_op_rgt_0')
// (15, 5, 'sp4_h_r_21')
// (15, 5, 'sp4_r_v_b_0')
// (15, 6, 'neigh_op_bnr_0')
// (15, 6, 'sp4_r_v_b_45')
// (15, 7, 'sp4_r_v_b_32')
// (15, 8, 'sp4_r_v_b_21')
// (15, 9, 'sp4_r_v_b_8')
// (16, 1, 'sp4_v_t_37')
// (16, 2, 'sp4_v_b_37')
// (16, 3, 'sp4_v_b_24')
// (16, 4, 'neigh_op_top_0')
// (16, 4, 'sp4_v_b_13')
// (16, 5, 'lutff_0/out')
// (16, 5, 'sp4_h_r_32')
// (16, 5, 'sp4_v_b_0')
// (16, 5, 'sp4_v_t_45')
// (16, 6, 'neigh_op_bot_0')
// (16, 6, 'sp4_v_b_45')
// (16, 7, 'sp4_v_b_32')
// (16, 8, 'local_g1_5')
// (16, 8, 'lutff_0/in_2')
// (16, 8, 'lutff_4/in_0')
// (16, 8, 'sp4_v_b_21')
// (16, 9, 'sp4_v_b_8')
// (17, 4, 'neigh_op_tnl_0')
// (17, 5, 'neigh_op_lft_0')
// (17, 5, 'sp4_h_r_45')
// (17, 6, 'neigh_op_bnl_0')
// (18, 5, 'sp4_h_l_45')

wire n1915;
// (13, 7, 'local_g0_0')
// (13, 7, 'lutff_6/in_0')
// (13, 7, 'sp4_h_r_8')
// (14, 6, 'neigh_op_tnr_0')
// (14, 7, 'neigh_op_rgt_0')
// (14, 7, 'sp4_h_r_21')
// (14, 8, 'neigh_op_bnr_0')
// (15, 6, 'neigh_op_top_0')
// (15, 7, 'lutff_0/out')
// (15, 7, 'sp4_h_r_32')
// (15, 8, 'neigh_op_bot_0')
// (16, 6, 'neigh_op_tnl_0')
// (16, 7, 'neigh_op_lft_0')
// (16, 7, 'sp4_h_r_45')
// (16, 8, 'neigh_op_bnl_0')
// (17, 7, 'sp4_h_l_45')

wire n1916;
// (13, 7, 'local_g3_6')
// (13, 7, 'lutff_3/in_2')
// (13, 7, 'neigh_op_tnr_6')
// (13, 8, 'neigh_op_rgt_6')
// (13, 9, 'neigh_op_bnr_6')
// (14, 7, 'neigh_op_top_6')
// (14, 8, 'lutff_6/out')
// (14, 9, 'neigh_op_bot_6')
// (15, 7, 'neigh_op_tnl_6')
// (15, 8, 'neigh_op_lft_6')
// (15, 9, 'neigh_op_bnl_6')

wire n1917;
// (13, 7, 'neigh_op_tnr_0')
// (13, 8, 'local_g2_0')
// (13, 8, 'lutff_5/in_1')
// (13, 8, 'neigh_op_rgt_0')
// (13, 9, 'neigh_op_bnr_0')
// (14, 7, 'neigh_op_top_0')
// (14, 8, 'lutff_0/out')
// (14, 9, 'neigh_op_bot_0')
// (15, 7, 'neigh_op_tnl_0')
// (15, 8, 'neigh_op_lft_0')
// (15, 9, 'neigh_op_bnl_0')

wire n1918;
// (13, 7, 'neigh_op_tnr_1')
// (13, 8, 'neigh_op_rgt_1')
// (13, 9, 'neigh_op_bnr_1')
// (14, 7, 'neigh_op_top_1')
// (14, 8, 'local_g2_1')
// (14, 8, 'lutff_1/out')
// (14, 8, 'lutff_4/in_3')
// (14, 9, 'neigh_op_bot_1')
// (15, 7, 'neigh_op_tnl_1')
// (15, 8, 'neigh_op_lft_1')
// (15, 9, 'neigh_op_bnl_1')

wire n1919;
// (13, 7, 'neigh_op_tnr_2')
// (13, 8, 'neigh_op_rgt_2')
// (13, 9, 'neigh_op_bnr_2')
// (14, 7, 'neigh_op_top_2')
// (14, 8, 'local_g1_2')
// (14, 8, 'lutff_2/out')
// (14, 8, 'lutff_4/in_1')
// (14, 9, 'neigh_op_bot_2')
// (15, 7, 'neigh_op_tnl_2')
// (15, 8, 'neigh_op_lft_2')
// (15, 9, 'neigh_op_bnl_2')

wire n1920;
// (13, 7, 'neigh_op_tnr_3')
// (13, 8, 'neigh_op_rgt_3')
// (13, 9, 'neigh_op_bnr_3')
// (14, 7, 'neigh_op_top_3')
// (14, 8, 'local_g2_3')
// (14, 8, 'lutff_0/in_3')
// (14, 8, 'lutff_3/out')
// (14, 9, 'neigh_op_bot_3')
// (15, 7, 'neigh_op_tnl_3')
// (15, 8, 'neigh_op_lft_3')
// (15, 9, 'neigh_op_bnl_3')

wire n1921;
// (13, 7, 'neigh_op_tnr_4')
// (13, 8, 'neigh_op_rgt_4')
// (13, 9, 'neigh_op_bnr_4')
// (14, 7, 'neigh_op_top_4')
// (14, 8, 'local_g1_4')
// (14, 8, 'lutff_0/in_1')
// (14, 8, 'lutff_4/out')
// (14, 9, 'neigh_op_bot_4')
// (15, 7, 'neigh_op_tnl_4')
// (15, 8, 'neigh_op_lft_4')
// (15, 9, 'neigh_op_bnl_4')

wire n1922;
// (13, 7, 'neigh_op_tnr_7')
// (13, 8, 'neigh_op_rgt_7')
// (13, 9, 'neigh_op_bnr_7')
// (14, 7, 'neigh_op_top_7')
// (14, 8, 'local_g3_7')
// (14, 8, 'lutff_4/in_0')
// (14, 8, 'lutff_7/out')
// (14, 9, 'neigh_op_bot_7')
// (15, 7, 'neigh_op_tnl_7')
// (15, 8, 'neigh_op_lft_7')
// (15, 9, 'neigh_op_bnl_7')

reg n1923 = 0;
// (13, 7, 'sp4_h_r_2')
// (14, 6, 'neigh_op_tnr_5')
// (14, 7, 'neigh_op_rgt_5')
// (14, 7, 'sp4_h_r_15')
// (14, 8, 'neigh_op_bnr_5')
// (15, 6, 'local_g1_5')
// (15, 6, 'lutff_7/in_1')
// (15, 6, 'neigh_op_top_5')
// (15, 7, 'lutff_5/out')
// (15, 7, 'sp4_h_r_26')
// (15, 8, 'neigh_op_bot_5')
// (16, 6, 'neigh_op_tnl_5')
// (16, 7, 'local_g0_5')
// (16, 7, 'lutff_7/in_2')
// (16, 7, 'neigh_op_lft_5')
// (16, 7, 'sp4_h_r_39')
// (16, 8, 'neigh_op_bnl_5')
// (16, 8, 'sp4_r_v_b_42')
// (16, 9, 'sp4_r_v_b_31')
// (16, 10, 'sp4_r_v_b_18')
// (16, 11, 'sp4_r_v_b_7')
// (17, 7, 'sp4_h_l_39')
// (17, 7, 'sp4_v_t_42')
// (17, 8, 'local_g3_2')
// (17, 8, 'lutff_2/in_1')
// (17, 8, 'sp4_v_b_42')
// (17, 9, 'sp4_v_b_31')
// (17, 10, 'sp4_v_b_18')
// (17, 11, 'sp4_v_b_7')

wire n1924;
// (13, 7, 'sp4_h_r_4')
// (14, 7, 'local_g1_1')
// (14, 7, 'lutff_7/in_1')
// (14, 7, 'sp4_h_r_17')
// (15, 4, 'neigh_op_tnr_1')
// (15, 5, 'neigh_op_rgt_1')
// (15, 6, 'neigh_op_bnr_1')
// (15, 7, 'sp4_h_r_28')
// (16, 4, 'neigh_op_top_1')
// (16, 4, 'sp4_r_v_b_46')
// (16, 5, 'lutff_1/out')
// (16, 5, 'sp4_r_v_b_35')
// (16, 6, 'neigh_op_bot_1')
// (16, 6, 'sp4_r_v_b_22')
// (16, 7, 'sp4_h_r_41')
// (16, 7, 'sp4_r_v_b_11')
// (17, 3, 'sp4_v_t_46')
// (17, 4, 'neigh_op_tnl_1')
// (17, 4, 'sp4_v_b_46')
// (17, 5, 'neigh_op_lft_1')
// (17, 5, 'sp4_v_b_35')
// (17, 6, 'neigh_op_bnl_1')
// (17, 6, 'sp4_v_b_22')
// (17, 7, 'sp4_h_l_41')
// (17, 7, 'sp4_v_b_11')

reg n1925 = 0;
// (13, 7, 'sp4_r_v_b_41')
// (13, 8, 'sp4_r_v_b_28')
// (13, 9, 'neigh_op_tnr_2')
// (13, 9, 'sp4_r_v_b_17')
// (13, 10, 'neigh_op_rgt_2')
// (13, 10, 'sp4_r_v_b_36')
// (13, 10, 'sp4_r_v_b_4')
// (13, 11, 'neigh_op_bnr_2')
// (13, 11, 'sp4_r_v_b_25')
// (13, 12, 'sp4_r_v_b_12')
// (13, 13, 'sp4_r_v_b_1')
// (14, 6, 'sp4_v_t_41')
// (14, 7, 'sp4_v_b_41')
// (14, 8, 'local_g3_4')
// (14, 8, 'lutff_6/in_1')
// (14, 8, 'sp4_r_v_b_45')
// (14, 8, 'sp4_v_b_28')
// (14, 9, 'neigh_op_top_2')
// (14, 9, 'sp4_r_v_b_32')
// (14, 9, 'sp4_v_b_17')
// (14, 9, 'sp4_v_t_36')
// (14, 10, 'local_g2_2')
// (14, 10, 'lutff_0/in_0')
// (14, 10, 'lutff_2/out')
// (14, 10, 'sp4_r_v_b_21')
// (14, 10, 'sp4_v_b_36')
// (14, 10, 'sp4_v_b_4')
// (14, 11, 'neigh_op_bot_2')
// (14, 11, 'sp4_r_v_b_8')
// (14, 11, 'sp4_v_b_25')
// (14, 12, 'local_g0_4')
// (14, 12, 'lutff_3/in_1')
// (14, 12, 'sp4_v_b_12')
// (14, 13, 'sp4_v_b_1')
// (15, 7, 'sp4_v_t_45')
// (15, 8, 'local_g2_5')
// (15, 8, 'lutff_2/in_3')
// (15, 8, 'sp4_v_b_45')
// (15, 9, 'neigh_op_tnl_2')
// (15, 9, 'sp4_v_b_32')
// (15, 10, 'neigh_op_lft_2')
// (15, 10, 'sp4_v_b_21')
// (15, 11, 'neigh_op_bnl_2')
// (15, 11, 'sp4_v_b_8')

reg n1926 = 0;
// (13, 7, 'sp4_r_v_b_45')
// (13, 8, 'sp4_r_v_b_32')
// (13, 9, 'neigh_op_tnr_4')
// (13, 9, 'sp4_r_v_b_21')
// (13, 10, 'neigh_op_rgt_4')
// (13, 10, 'sp4_r_v_b_8')
// (13, 11, 'neigh_op_bnr_4')
// (13, 11, 'sp4_r_v_b_46')
// (13, 12, 'sp4_r_v_b_35')
// (13, 13, 'sp4_r_v_b_22')
// (13, 14, 'sp4_r_v_b_11')
// (14, 6, 'sp4_v_t_45')
// (14, 7, 'local_g3_5')
// (14, 7, 'lutff_3/in_1')
// (14, 7, 'sp4_v_b_45')
// (14, 8, 'local_g3_0')
// (14, 8, 'lutff_1/in_2')
// (14, 8, 'sp4_v_b_32')
// (14, 9, 'neigh_op_top_4')
// (14, 9, 'sp4_v_b_21')
// (14, 10, 'local_g2_4')
// (14, 10, 'lutff_2/in_2')
// (14, 10, 'lutff_4/out')
// (14, 10, 'sp4_v_b_8')
// (14, 10, 'sp4_v_t_46')
// (14, 11, 'neigh_op_bot_4')
// (14, 11, 'sp4_v_b_46')
// (14, 12, 'sp4_v_b_35')
// (14, 13, 'sp4_v_b_22')
// (14, 14, 'local_g1_3')
// (14, 14, 'lutff_1/in_1')
// (14, 14, 'sp4_v_b_11')
// (15, 9, 'neigh_op_tnl_4')
// (15, 10, 'neigh_op_lft_4')
// (15, 11, 'neigh_op_bnl_4')

reg n1927 = 0;
// (13, 8, 'neigh_op_tnr_1')
// (13, 9, 'neigh_op_rgt_1')
// (13, 9, 'sp4_h_r_7')
// (13, 10, 'neigh_op_bnr_1')
// (14, 8, 'neigh_op_top_1')
// (14, 9, 'lutff_1/out')
// (14, 9, 'sp4_h_r_18')
// (14, 9, 'sp4_h_r_2')
// (14, 10, 'neigh_op_bot_1')
// (15, 8, 'neigh_op_tnl_1')
// (15, 9, 'local_g1_1')
// (15, 9, 'lutff_7/in_3')
// (15, 9, 'neigh_op_lft_1')
// (15, 9, 'sp4_h_r_15')
// (15, 9, 'sp4_h_r_31')
// (15, 10, 'neigh_op_bnl_1')
// (16, 6, 'sp4_r_v_b_42')
// (16, 7, 'sp4_r_v_b_31')
// (16, 8, 'local_g3_2')
// (16, 8, 'lutff_6/in_1')
// (16, 8, 'sp4_r_v_b_18')
// (16, 9, 'local_g3_2')
// (16, 9, 'lutff_0/in_1')
// (16, 9, 'sp4_h_r_26')
// (16, 9, 'sp4_h_r_42')
// (16, 9, 'sp4_r_v_b_7')
// (17, 5, 'sp4_v_t_42')
// (17, 6, 'sp4_v_b_42')
// (17, 7, 'sp4_v_b_31')
// (17, 8, 'sp4_v_b_18')
// (17, 9, 'sp4_h_l_42')
// (17, 9, 'sp4_h_r_39')
// (17, 9, 'sp4_v_b_7')
// (18, 9, 'sp4_h_l_39')

reg n1928 = 0;
// (13, 8, 'neigh_op_tnr_2')
// (13, 9, 'neigh_op_rgt_2')
// (13, 9, 'sp4_h_r_9')
// (13, 10, 'neigh_op_bnr_2')
// (14, 8, 'neigh_op_top_2')
// (14, 9, 'lutff_2/out')
// (14, 9, 'sp4_h_r_20')
// (14, 9, 'sp4_h_r_4')
// (14, 10, 'neigh_op_bot_2')
// (15, 8, 'neigh_op_tnl_2')
// (15, 9, 'local_g0_2')
// (15, 9, 'lutff_5/in_3')
// (15, 9, 'neigh_op_lft_2')
// (15, 9, 'sp4_h_r_17')
// (15, 9, 'sp4_h_r_33')
// (15, 10, 'neigh_op_bnl_2')
// (16, 6, 'sp4_r_v_b_44')
// (16, 7, 'sp4_r_v_b_33')
// (16, 8, 'local_g3_4')
// (16, 8, 'lutff_4/in_1')
// (16, 8, 'sp4_r_v_b_20')
// (16, 9, 'sp4_h_r_28')
// (16, 9, 'sp4_h_r_44')
// (16, 9, 'sp4_r_v_b_9')
// (17, 5, 'sp4_v_t_44')
// (17, 6, 'sp4_v_b_44')
// (17, 7, 'sp4_v_b_33')
// (17, 8, 'sp4_v_b_20')
// (17, 9, 'local_g3_1')
// (17, 9, 'lutff_7/in_3')
// (17, 9, 'sp4_h_l_44')
// (17, 9, 'sp4_h_r_41')
// (17, 9, 'sp4_v_b_9')
// (18, 9, 'sp4_h_l_41')

reg n1929 = 0;
// (13, 8, 'neigh_op_tnr_3')
// (13, 9, 'neigh_op_rgt_3')
// (13, 10, 'neigh_op_bnr_3')
// (14, 7, 'sp4_r_v_b_47')
// (14, 8, 'neigh_op_top_3')
// (14, 8, 'sp4_r_v_b_34')
// (14, 9, 'lutff_3/out')
// (14, 9, 'sp4_r_v_b_23')
// (14, 10, 'neigh_op_bot_3')
// (14, 10, 'sp4_r_v_b_10')
// (15, 6, 'sp4_v_t_47')
// (15, 7, 'sp4_v_b_47')
// (15, 8, 'local_g2_3')
// (15, 8, 'local_g3_3')
// (15, 8, 'lutff_5/in_1')
// (15, 8, 'lutff_7/in_0')
// (15, 8, 'neigh_op_tnl_3')
// (15, 8, 'sp4_v_b_34')
// (15, 9, 'neigh_op_lft_3')
// (15, 9, 'sp4_v_b_23')
// (15, 10, 'neigh_op_bnl_3')
// (15, 10, 'sp4_h_r_10')
// (15, 10, 'sp4_v_b_10')
// (16, 10, 'local_g1_7')
// (16, 10, 'lutff_7/in_3')
// (16, 10, 'sp4_h_r_23')
// (17, 10, 'sp4_h_r_34')
// (18, 10, 'sp4_h_r_47')
// (19, 10, 'sp4_h_l_47')

reg n1930 = 0;
// (13, 8, 'neigh_op_tnr_6')
// (13, 9, 'neigh_op_rgt_6')
// (13, 9, 'sp4_h_r_1')
// (13, 10, 'neigh_op_bnr_6')
// (14, 8, 'neigh_op_top_6')
// (14, 9, 'lutff_6/out')
// (14, 9, 'sp4_h_r_12')
// (14, 10, 'neigh_op_bot_6')
// (15, 8, 'local_g2_6')
// (15, 8, 'lutff_3/in_1')
// (15, 8, 'neigh_op_tnl_6')
// (15, 9, 'local_g0_6')
// (15, 9, 'lutff_2/in_0')
// (15, 9, 'neigh_op_lft_6')
// (15, 9, 'sp4_h_r_25')
// (15, 10, 'neigh_op_bnl_6')
// (16, 9, 'local_g2_4')
// (16, 9, 'lutff_5/in_1')
// (16, 9, 'sp4_h_r_36')
// (17, 9, 'sp4_h_l_36')

reg n1931 = 0;
// (13, 8, 'sp4_h_r_10')
// (14, 8, 'local_g0_7')
// (14, 8, 'lutff_7/in_0')
// (14, 8, 'sp4_h_r_23')
// (15, 1, 'neigh_op_tnr_6')
// (15, 2, 'local_g3_6')
// (15, 2, 'lutff_1/in_2')
// (15, 2, 'neigh_op_rgt_6')
// (15, 2, 'sp4_r_v_b_44')
// (15, 3, 'neigh_op_bnr_6')
// (15, 3, 'sp4_r_v_b_33')
// (15, 4, 'sp4_r_v_b_20')
// (15, 5, 'sp4_r_v_b_9')
// (15, 6, 'sp4_r_v_b_37')
// (15, 7, 'sp4_r_v_b_24')
// (15, 8, 'sp4_h_r_34')
// (15, 8, 'sp4_r_v_b_13')
// (15, 9, 'local_g1_0')
// (15, 9, 'lutff_7/in_2')
// (15, 9, 'sp4_r_v_b_0')
// (16, 1, 'neigh_op_top_6')
// (16, 1, 'sp4_r_v_b_40')
// (16, 1, 'sp4_v_t_44')
// (16, 2, 'lutff_6/out')
// (16, 2, 'sp4_r_v_b_29')
// (16, 2, 'sp4_v_b_44')
// (16, 3, 'neigh_op_bot_6')
// (16, 3, 'sp4_r_v_b_16')
// (16, 3, 'sp4_v_b_33')
// (16, 4, 'sp4_r_v_b_5')
// (16, 4, 'sp4_v_b_20')
// (16, 5, 'local_g1_1')
// (16, 5, 'lutff_7/in_3')
// (16, 5, 'sp4_r_v_b_40')
// (16, 5, 'sp4_v_b_9')
// (16, 5, 'sp4_v_t_37')
// (16, 6, 'sp4_r_v_b_29')
// (16, 6, 'sp4_v_b_37')
// (16, 7, 'sp4_r_v_b_16')
// (16, 7, 'sp4_v_b_24')
// (16, 8, 'local_g0_5')
// (16, 8, 'lutff_1/in_2')
// (16, 8, 'sp4_h_r_47')
// (16, 8, 'sp4_r_v_b_5')
// (16, 8, 'sp4_v_b_13')
// (16, 9, 'sp4_v_b_0')
// (17, 0, 'span4_vert_40')
// (17, 1, 'neigh_op_tnl_6')
// (17, 1, 'sp4_v_b_40')
// (17, 2, 'neigh_op_lft_6')
// (17, 2, 'sp4_v_b_29')
// (17, 3, 'neigh_op_bnl_6')
// (17, 3, 'sp4_v_b_16')
// (17, 4, 'sp4_v_b_5')
// (17, 4, 'sp4_v_t_40')
// (17, 5, 'sp4_v_b_40')
// (17, 6, 'sp4_v_b_29')
// (17, 7, 'sp4_v_b_16')
// (17, 8, 'sp4_h_l_47')
// (17, 8, 'sp4_v_b_5')

reg n1932 = 0;
// (13, 8, 'sp4_h_r_3')
// (14, 8, 'local_g1_6')
// (14, 8, 'lutff_6/in_3')
// (14, 8, 'sp4_h_r_14')
// (15, 1, 'sp4_r_v_b_36')
// (15, 2, 'neigh_op_tnr_6')
// (15, 2, 'sp4_r_v_b_25')
// (15, 3, 'neigh_op_rgt_6')
// (15, 3, 'sp4_r_v_b_12')
// (15, 4, 'local_g1_6')
// (15, 4, 'lutff_4/in_3')
// (15, 4, 'neigh_op_bnr_6')
// (15, 4, 'sp4_r_v_b_1')
// (15, 5, 'sp4_r_v_b_41')
// (15, 6, 'sp4_r_v_b_28')
// (15, 7, 'sp4_r_v_b_17')
// (15, 8, 'local_g1_4')
// (15, 8, 'lutff_5/in_2')
// (15, 8, 'sp4_h_r_27')
// (15, 8, 'sp4_r_v_b_4')
// (16, 0, 'span4_vert_36')
// (16, 1, 'sp4_r_v_b_37')
// (16, 1, 'sp4_v_b_36')
// (16, 2, 'neigh_op_top_6')
// (16, 2, 'sp4_r_v_b_24')
// (16, 2, 'sp4_v_b_25')
// (16, 3, 'lutff_6/out')
// (16, 3, 'sp4_r_v_b_13')
// (16, 3, 'sp4_v_b_12')
// (16, 4, 'neigh_op_bot_6')
// (16, 4, 'sp4_r_v_b_0')
// (16, 4, 'sp4_v_b_1')
// (16, 4, 'sp4_v_t_41')
// (16, 5, 'sp4_r_v_b_38')
// (16, 5, 'sp4_v_b_41')
// (16, 6, 'sp4_r_v_b_27')
// (16, 6, 'sp4_v_b_28')
// (16, 7, 'sp4_r_v_b_14')
// (16, 7, 'sp4_v_b_17')
// (16, 8, 'sp4_h_r_38')
// (16, 8, 'sp4_r_v_b_3')
// (16, 8, 'sp4_v_b_4')
// (17, 0, 'span4_vert_37')
// (17, 1, 'sp4_v_b_37')
// (17, 2, 'neigh_op_tnl_6')
// (17, 2, 'sp4_v_b_24')
// (17, 3, 'neigh_op_lft_6')
// (17, 3, 'sp4_v_b_13')
// (17, 4, 'neigh_op_bnl_6')
// (17, 4, 'sp4_v_b_0')
// (17, 4, 'sp4_v_t_38')
// (17, 5, 'sp4_v_b_38')
// (17, 6, 'sp4_v_b_27')
// (17, 7, 'sp4_v_b_14')
// (17, 8, 'sp4_h_l_38')
// (17, 8, 'sp4_v_b_3')

reg n1933 = 0;
// (13, 8, 'sp4_r_v_b_45')
// (13, 9, 'sp4_r_v_b_32')
// (13, 10, 'neigh_op_tnr_4')
// (13, 10, 'sp4_r_v_b_21')
// (13, 11, 'neigh_op_rgt_4')
// (13, 11, 'sp4_r_v_b_8')
// (13, 12, 'neigh_op_bnr_4')
// (14, 7, 'local_g0_1')
// (14, 7, 'lutff_0/in_1')
// (14, 7, 'sp4_h_r_1')
// (14, 7, 'sp4_v_t_45')
// (14, 8, 'sp4_v_b_45')
// (14, 9, 'sp4_v_b_32')
// (14, 10, 'local_g0_4')
// (14, 10, 'lutff_6/in_0')
// (14, 10, 'neigh_op_top_4')
// (14, 10, 'sp4_v_b_21')
// (14, 11, 'lutff_4/out')
// (14, 11, 'sp4_v_b_8')
// (14, 12, 'local_g1_4')
// (14, 12, 'lutff_1/in_0')
// (14, 12, 'neigh_op_bot_4')
// (15, 7, 'sp4_h_r_12')
// (15, 10, 'neigh_op_tnl_4')
// (15, 11, 'neigh_op_lft_4')
// (15, 12, 'neigh_op_bnl_4')
// (16, 7, 'sp4_h_r_25')
// (17, 7, 'sp4_h_r_36')
// (18, 7, 'sp4_h_l_36')

reg n1934 = 0;
// (13, 9, 'neigh_op_tnr_0')
// (13, 9, 'sp4_r_v_b_45')
// (13, 10, 'neigh_op_rgt_0')
// (13, 10, 'sp4_r_v_b_32')
// (13, 11, 'neigh_op_bnr_0')
// (13, 11, 'sp4_r_v_b_21')
// (13, 12, 'sp4_r_v_b_8')
// (14, 0, 'span12_vert_19')
// (14, 1, 'sp12_v_b_19')
// (14, 2, 'sp12_v_b_16')
// (14, 3, 'sp12_v_b_15')
// (14, 4, 'sp12_v_b_12')
// (14, 5, 'sp12_v_b_11')
// (14, 6, 'local_g2_0')
// (14, 6, 'lutff_2/in_0')
// (14, 6, 'lutff_4/in_0')
// (14, 6, 'sp12_v_b_8')
// (14, 7, 'sp12_v_b_7')
// (14, 8, 'sp12_v_b_4')
// (14, 8, 'sp4_v_t_45')
// (14, 9, 'neigh_op_top_0')
// (14, 9, 'sp12_v_b_3')
// (14, 9, 'sp4_v_b_45')
// (14, 10, 'lutff_0/out')
// (14, 10, 'sp12_v_b_0')
// (14, 10, 'sp4_v_b_32')
// (14, 11, 'local_g1_0')
// (14, 11, 'lutff_1/in_2')
// (14, 11, 'neigh_op_bot_0')
// (14, 11, 'sp4_v_b_21')
// (14, 12, 'local_g0_0')
// (14, 12, 'lutff_6/in_2')
// (14, 12, 'sp4_v_b_8')
// (15, 9, 'neigh_op_tnl_0')
// (15, 10, 'neigh_op_lft_0')
// (15, 11, 'neigh_op_bnl_0')

wire n1935;
// (13, 9, 'neigh_op_tnr_5')
// (13, 10, 'neigh_op_rgt_5')
// (13, 11, 'neigh_op_bnr_5')
// (14, 9, 'neigh_op_top_5')
// (14, 10, 'local_g0_5')
// (14, 10, 'lutff_5/out')
// (14, 10, 'lutff_7/in_2')
// (14, 11, 'neigh_op_bot_5')
// (15, 9, 'neigh_op_tnl_5')
// (15, 10, 'neigh_op_lft_5')
// (15, 11, 'neigh_op_bnl_5')

reg n1936 = 0;
// (13, 9, 'neigh_op_tnr_6')
// (13, 10, 'neigh_op_rgt_6')
// (13, 10, 'sp4_r_v_b_44')
// (13, 11, 'neigh_op_bnr_6')
// (13, 11, 'sp4_r_v_b_33')
// (13, 12, 'sp4_r_v_b_20')
// (13, 13, 'sp4_r_v_b_9')
// (14, 9, 'local_g1_6')
// (14, 9, 'lutff_0/in_3')
// (14, 9, 'neigh_op_top_6')
// (14, 9, 'sp4_v_t_44')
// (14, 10, 'local_g3_6')
// (14, 10, 'lutff_4/in_3')
// (14, 10, 'lutff_6/out')
// (14, 10, 'sp4_v_b_44')
// (14, 11, 'neigh_op_bot_6')
// (14, 11, 'sp4_v_b_33')
// (14, 12, 'sp4_v_b_20')
// (14, 13, 'local_g1_1')
// (14, 13, 'lutff_3/in_3')
// (14, 13, 'sp4_v_b_9')
// (15, 9, 'neigh_op_tnl_6')
// (15, 10, 'neigh_op_lft_6')
// (15, 11, 'neigh_op_bnl_6')

wire n1937;
// (13, 9, 'neigh_op_tnr_7')
// (13, 10, 'neigh_op_rgt_7')
// (13, 11, 'neigh_op_bnr_7')
// (14, 4, 'sp4_r_v_b_39')
// (14, 5, 'sp4_r_v_b_26')
// (14, 6, 'sp4_r_v_b_15')
// (14, 7, 'local_g1_2')
// (14, 7, 'lutff_7/in_2')
// (14, 7, 'sp4_r_v_b_2')
// (14, 8, 'sp4_r_v_b_39')
// (14, 9, 'neigh_op_top_7')
// (14, 9, 'sp4_r_v_b_26')
// (14, 10, 'lutff_7/out')
// (14, 10, 'sp4_r_v_b_15')
// (14, 11, 'neigh_op_bot_7')
// (14, 11, 'sp4_r_v_b_2')
// (15, 3, 'sp4_v_t_39')
// (15, 4, 'sp4_v_b_39')
// (15, 5, 'sp4_v_b_26')
// (15, 6, 'sp4_v_b_15')
// (15, 7, 'sp4_v_b_2')
// (15, 7, 'sp4_v_t_39')
// (15, 8, 'sp4_v_b_39')
// (15, 9, 'neigh_op_tnl_7')
// (15, 9, 'sp4_v_b_26')
// (15, 10, 'neigh_op_lft_7')
// (15, 10, 'sp4_v_b_15')
// (15, 11, 'neigh_op_bnl_7')
// (15, 11, 'sp4_v_b_2')

reg n1938 = 0;
// (13, 9, 'sp4_h_r_3')
// (14, 9, 'local_g0_6')
// (14, 9, 'lutff_3/in_3')
// (14, 9, 'sp4_h_r_14')
// (15, 6, 'sp4_r_v_b_46')
// (15, 7, 'sp4_r_v_b_35')
// (15, 8, 'sp4_r_v_b_22')
// (15, 9, 'sp4_h_r_27')
// (15, 9, 'sp4_r_v_b_11')
// (15, 10, 'local_g3_5')
// (15, 10, 'lutff_3/in_1')
// (15, 10, 'sp4_r_v_b_45')
// (15, 11, 'local_g2_0')
// (15, 11, 'lutff_5/in_3')
// (15, 11, 'sp4_r_v_b_32')
// (15, 12, 'neigh_op_tnr_4')
// (15, 12, 'sp4_r_v_b_21')
// (15, 13, 'neigh_op_rgt_4')
// (15, 13, 'sp4_r_v_b_8')
// (15, 14, 'neigh_op_bnr_4')
// (16, 5, 'sp4_v_t_46')
// (16, 6, 'sp4_v_b_46')
// (16, 7, 'sp4_v_b_35')
// (16, 8, 'local_g1_6')
// (16, 8, 'lutff_7/in_0')
// (16, 8, 'sp4_v_b_22')
// (16, 9, 'sp4_h_r_38')
// (16, 9, 'sp4_v_b_11')
// (16, 9, 'sp4_v_t_45')
// (16, 10, 'sp4_r_v_b_44')
// (16, 10, 'sp4_v_b_45')
// (16, 11, 'local_g3_0')
// (16, 11, 'lutff_7/in_0')
// (16, 11, 'sp4_r_v_b_33')
// (16, 11, 'sp4_v_b_32')
// (16, 12, 'local_g0_4')
// (16, 12, 'lutff_7/in_3')
// (16, 12, 'neigh_op_top_4')
// (16, 12, 'sp4_r_v_b_20')
// (16, 12, 'sp4_r_v_b_36')
// (16, 12, 'sp4_v_b_21')
// (16, 13, 'local_g1_4')
// (16, 13, 'lutff_4/out')
// (16, 13, 'lutff_5/in_2')
// (16, 13, 'sp4_r_v_b_25')
// (16, 13, 'sp4_r_v_b_9')
// (16, 13, 'sp4_v_b_8')
// (16, 14, 'neigh_op_bot_4')
// (16, 14, 'sp4_r_v_b_12')
// (16, 15, 'sp4_r_v_b_1')
// (17, 9, 'sp4_h_l_38')
// (17, 9, 'sp4_h_r_9')
// (17, 9, 'sp4_v_t_44')
// (17, 10, 'sp4_v_b_44')
// (17, 11, 'sp4_h_r_1')
// (17, 11, 'sp4_v_b_33')
// (17, 11, 'sp4_v_t_36')
// (17, 12, 'neigh_op_tnl_4')
// (17, 12, 'sp4_v_b_20')
// (17, 12, 'sp4_v_b_36')
// (17, 13, 'neigh_op_lft_4')
// (17, 13, 'sp4_v_b_25')
// (17, 13, 'sp4_v_b_9')
// (17, 14, 'neigh_op_bnl_4')
// (17, 14, 'sp4_v_b_12')
// (17, 15, 'sp4_v_b_1')
// (18, 9, 'sp4_h_r_20')
// (18, 11, 'sp4_h_r_12')
// (19, 9, 'sp4_h_r_33')
// (19, 11, 'sp4_h_r_25')
// (20, 9, 'local_g3_4')
// (20, 9, 'lutff_1/in_0')
// (20, 9, 'sp4_h_r_44')
// (20, 11, 'sp4_h_r_36')
// (21, 9, 'sp4_h_l_44')
// (21, 11, 'local_g1_4')
// (21, 11, 'lutff_5/in_2')
// (21, 11, 'sp4_h_l_36')
// (21, 11, 'sp4_h_r_4')
// (22, 11, 'sp4_h_r_17')
// (23, 11, 'sp4_h_r_28')
// (24, 11, 'sp4_h_r_41')
// (25, 11, 'sp4_h_l_41')

wire n1939;
// (13, 10, 'neigh_op_tnr_2')
// (13, 11, 'neigh_op_rgt_2')
// (13, 12, 'local_g1_2')
// (13, 12, 'lutff_3/in_0')
// (13, 12, 'neigh_op_bnr_2')
// (14, 10, 'neigh_op_top_2')
// (14, 11, 'lutff_2/out')
// (14, 12, 'neigh_op_bot_2')
// (15, 10, 'neigh_op_tnl_2')
// (15, 11, 'neigh_op_lft_2')
// (15, 12, 'neigh_op_bnl_2')

wire n1940;
// (13, 10, 'neigh_op_tnr_5')
// (13, 11, 'neigh_op_rgt_5')
// (13, 12, 'neigh_op_bnr_5')
// (14, 10, 'neigh_op_top_5')
// (14, 11, 'local_g3_5')
// (14, 11, 'lutff_2/in_2')
// (14, 11, 'lutff_5/out')
// (14, 12, 'neigh_op_bot_5')
// (15, 10, 'neigh_op_tnl_5')
// (15, 11, 'neigh_op_lft_5')
// (15, 12, 'neigh_op_bnl_5')

wire n1941;
// (13, 11, 'neigh_op_tnr_0')
// (13, 12, 'neigh_op_rgt_0')
// (13, 13, 'neigh_op_bnr_0')
// (14, 11, 'neigh_op_top_0')
// (14, 12, 'lutff_0/out')
// (14, 13, 'neigh_op_bot_0')
// (15, 11, 'neigh_op_tnl_0')
// (15, 12, 'local_g0_0')
// (15, 12, 'lutff_4/in_0')
// (15, 12, 'neigh_op_lft_0')
// (15, 13, 'neigh_op_bnl_0')

wire n1942;
// (13, 11, 'neigh_op_tnr_1')
// (13, 12, 'neigh_op_rgt_1')
// (13, 13, 'neigh_op_bnr_1')
// (14, 11, 'neigh_op_top_1')
// (14, 12, 'local_g2_1')
// (14, 12, 'lutff_1/out')
// (14, 12, 'lutff_7/in_2')
// (14, 13, 'neigh_op_bot_1')
// (15, 11, 'neigh_op_tnl_1')
// (15, 12, 'neigh_op_lft_1')
// (15, 13, 'neigh_op_bnl_1')

wire n1943;
// (13, 11, 'neigh_op_tnr_2')
// (13, 12, 'neigh_op_rgt_2')
// (13, 13, 'neigh_op_bnr_2')
// (14, 11, 'neigh_op_top_2')
// (14, 12, 'lutff_2/out')
// (14, 13, 'neigh_op_bot_2')
// (15, 11, 'neigh_op_tnl_2')
// (15, 12, 'neigh_op_lft_2')
// (15, 13, 'local_g3_2')
// (15, 13, 'lutff_6/in_1')
// (15, 13, 'neigh_op_bnl_2')

wire n1944;
// (13, 11, 'neigh_op_tnr_3')
// (13, 12, 'neigh_op_rgt_3')
// (13, 13, 'neigh_op_bnr_3')
// (14, 11, 'neigh_op_top_3')
// (14, 12, 'lutff_3/out')
// (14, 13, 'local_g1_3')
// (14, 13, 'lutff_5/in_3')
// (14, 13, 'neigh_op_bot_3')
// (15, 11, 'neigh_op_tnl_3')
// (15, 12, 'neigh_op_lft_3')
// (15, 13, 'neigh_op_bnl_3')

wire n1945;
// (13, 11, 'neigh_op_tnr_4')
// (13, 12, 'neigh_op_rgt_4')
// (13, 13, 'neigh_op_bnr_4')
// (14, 11, 'neigh_op_top_4')
// (14, 12, 'lutff_4/out')
// (14, 13, 'neigh_op_bot_4')
// (15, 11, 'neigh_op_tnl_4')
// (15, 12, 'local_g1_4')
// (15, 12, 'lutff_4/in_1')
// (15, 12, 'neigh_op_lft_4')
// (15, 13, 'neigh_op_bnl_4')

wire n1946;
// (13, 11, 'neigh_op_tnr_5')
// (13, 12, 'neigh_op_rgt_5')
// (13, 13, 'neigh_op_bnr_5')
// (14, 11, 'neigh_op_top_5')
// (14, 12, 'lutff_5/out')
// (14, 13, 'local_g0_5')
// (14, 13, 'lutff_7/in_0')
// (14, 13, 'neigh_op_bot_5')
// (15, 11, 'neigh_op_tnl_5')
// (15, 12, 'neigh_op_lft_5')
// (15, 13, 'neigh_op_bnl_5')

wire n1947;
// (13, 11, 'neigh_op_tnr_6')
// (13, 12, 'neigh_op_rgt_6')
// (13, 13, 'neigh_op_bnr_6')
// (14, 11, 'neigh_op_top_6')
// (14, 11, 'sp4_r_v_b_40')
// (14, 12, 'lutff_6/out')
// (14, 12, 'sp4_r_v_b_29')
// (14, 13, 'neigh_op_bot_6')
// (14, 13, 'sp4_r_v_b_16')
// (14, 14, 'local_g1_5')
// (14, 14, 'lutff_2/in_2')
// (14, 14, 'sp4_r_v_b_5')
// (15, 10, 'sp4_v_t_40')
// (15, 11, 'neigh_op_tnl_6')
// (15, 11, 'sp4_v_b_40')
// (15, 12, 'neigh_op_lft_6')
// (15, 12, 'sp4_v_b_29')
// (15, 13, 'neigh_op_bnl_6')
// (15, 13, 'sp4_v_b_16')
// (15, 14, 'sp4_v_b_5')

wire n1948;
// (13, 11, 'neigh_op_tnr_7')
// (13, 12, 'neigh_op_rgt_7')
// (13, 13, 'neigh_op_bnr_7')
// (14, 11, 'neigh_op_top_7')
// (14, 12, 'lutff_7/out')
// (14, 13, 'local_g1_7')
// (14, 13, 'lutff_6/in_0')
// (14, 13, 'neigh_op_bot_7')
// (15, 11, 'neigh_op_tnl_7')
// (15, 12, 'neigh_op_lft_7')
// (15, 13, 'neigh_op_bnl_7')

wire n1949;
// (13, 12, 'neigh_op_tnr_1')
// (13, 13, 'local_g3_1')
// (13, 13, 'lutff_7/in_1')
// (13, 13, 'neigh_op_rgt_1')
// (13, 14, 'neigh_op_bnr_1')
// (14, 12, 'neigh_op_top_1')
// (14, 12, 'sp4_r_v_b_46')
// (14, 13, 'lutff_1/out')
// (14, 13, 'sp4_r_v_b_35')
// (14, 14, 'neigh_op_bot_1')
// (14, 14, 'sp4_r_v_b_22')
// (14, 15, 'sp4_r_v_b_11')
// (15, 11, 'sp4_v_t_46')
// (15, 12, 'neigh_op_tnl_1')
// (15, 12, 'sp4_v_b_46')
// (15, 13, 'neigh_op_lft_1')
// (15, 13, 'sp4_v_b_35')
// (15, 14, 'neigh_op_bnl_1')
// (15, 14, 'sp4_v_b_22')
// (15, 15, 'sp4_h_r_5')
// (15, 15, 'sp4_v_b_11')
// (16, 15, 'sp4_h_r_16')
// (17, 15, 'sp4_h_r_29')
// (18, 15, 'sp4_h_r_40')
// (19, 15, 'local_g1_5')
// (19, 15, 'ram/WDATA_8')
// (19, 15, 'sp4_h_l_40')
// (19, 15, 'sp4_h_r_5')
// (20, 15, 'sp4_h_r_16')
// (21, 15, 'sp4_h_r_29')
// (22, 15, 'sp4_h_r_40')
// (23, 15, 'sp4_h_l_40')

wire n1950;
// (13, 12, 'neigh_op_tnr_2')
// (13, 13, 'neigh_op_rgt_2')
// (13, 14, 'neigh_op_bnr_2')
// (14, 12, 'neigh_op_top_2')
// (14, 13, 'lutff_2/out')
// (14, 14, 'local_g0_2')
// (14, 14, 'lutff_0/in_2')
// (14, 14, 'neigh_op_bot_2')
// (15, 12, 'neigh_op_tnl_2')
// (15, 13, 'neigh_op_lft_2')
// (15, 14, 'neigh_op_bnl_2')

wire n1951;
// (13, 12, 'neigh_op_tnr_3')
// (13, 13, 'neigh_op_rgt_3')
// (13, 14, 'neigh_op_bnr_3')
// (14, 12, 'neigh_op_top_3')
// (14, 13, 'local_g3_3')
// (14, 13, 'lutff_3/out')
// (14, 13, 'lutff_7/in_3')
// (14, 14, 'neigh_op_bot_3')
// (15, 12, 'neigh_op_tnl_3')
// (15, 13, 'neigh_op_lft_3')
// (15, 14, 'neigh_op_bnl_3')

wire n1952;
// (13, 12, 'neigh_op_tnr_4')
// (13, 13, 'neigh_op_rgt_4')
// (13, 14, 'neigh_op_bnr_4')
// (14, 12, 'neigh_op_top_4')
// (14, 13, 'local_g1_4')
// (14, 13, 'lutff_4/out')
// (14, 13, 'lutff_7/in_2')
// (14, 14, 'neigh_op_bot_4')
// (15, 12, 'neigh_op_tnl_4')
// (15, 13, 'neigh_op_lft_4')
// (15, 14, 'neigh_op_bnl_4')

wire n1953;
// (13, 12, 'neigh_op_tnr_5')
// (13, 13, 'local_g3_5')
// (13, 13, 'lutff_4/in_0')
// (13, 13, 'neigh_op_rgt_5')
// (13, 14, 'neigh_op_bnr_5')
// (14, 12, 'neigh_op_top_5')
// (14, 13, 'lutff_5/out')
// (14, 13, 'sp4_r_v_b_43')
// (14, 14, 'neigh_op_bot_5')
// (14, 14, 'sp4_r_v_b_30')
// (14, 15, 'sp4_r_v_b_19')
// (14, 16, 'sp4_r_v_b_6')
// (15, 12, 'neigh_op_tnl_5')
// (15, 12, 'sp4_v_t_43')
// (15, 13, 'neigh_op_lft_5')
// (15, 13, 'sp4_v_b_43')
// (15, 14, 'neigh_op_bnl_5')
// (15, 14, 'sp4_v_b_30')
// (15, 15, 'sp4_v_b_19')
// (15, 16, 'sp4_h_r_0')
// (15, 16, 'sp4_v_b_6')
// (16, 16, 'sp4_h_r_13')
// (17, 16, 'sp4_h_r_24')
// (18, 16, 'sp4_h_r_37')
// (19, 16, 'local_g1_3')
// (19, 16, 'ram/WDATA_2')
// (19, 16, 'sp4_h_l_37')
// (19, 16, 'sp4_h_r_3')
// (20, 16, 'sp4_h_r_14')
// (21, 16, 'sp4_h_r_27')
// (22, 16, 'sp4_h_r_38')
// (23, 16, 'sp4_h_l_38')

wire n1954;
// (13, 12, 'neigh_op_tnr_6')
// (13, 13, 'local_g2_6')
// (13, 13, 'lutff_5/in_3')
// (13, 13, 'neigh_op_rgt_6')
// (13, 14, 'neigh_op_bnr_6')
// (14, 12, 'neigh_op_top_6')
// (14, 12, 'sp4_r_v_b_40')
// (14, 13, 'lutff_6/out')
// (14, 13, 'sp4_r_v_b_29')
// (14, 14, 'neigh_op_bot_6')
// (14, 14, 'sp4_r_v_b_16')
// (14, 15, 'sp4_r_v_b_5')
// (15, 11, 'sp4_v_t_40')
// (15, 12, 'neigh_op_tnl_6')
// (15, 12, 'sp4_v_b_40')
// (15, 13, 'neigh_op_lft_6')
// (15, 13, 'sp4_v_b_29')
// (15, 14, 'neigh_op_bnl_6')
// (15, 14, 'sp4_v_b_16')
// (15, 15, 'sp4_h_r_11')
// (15, 15, 'sp4_v_b_5')
// (16, 15, 'sp4_h_r_22')
// (17, 15, 'sp4_h_r_35')
// (18, 15, 'sp4_h_r_46')
// (19, 15, 'local_g0_2')
// (19, 15, 'ram/WDATA_12')
// (19, 15, 'sp4_h_l_46')
// (19, 15, 'sp4_h_r_2')
// (20, 15, 'sp4_h_r_15')
// (21, 15, 'sp4_h_r_26')
// (22, 15, 'sp4_h_r_39')
// (23, 15, 'sp4_h_l_39')

wire n1955;
// (13, 12, 'neigh_op_tnr_7')
// (13, 13, 'local_g3_7')
// (13, 13, 'lutff_6/in_2')
// (13, 13, 'neigh_op_rgt_7')
// (13, 14, 'neigh_op_bnr_7')
// (14, 12, 'neigh_op_top_7')
// (14, 13, 'lutff_7/out')
// (14, 13, 'sp4_r_v_b_47')
// (14, 14, 'neigh_op_bot_7')
// (14, 14, 'sp4_r_v_b_34')
// (14, 15, 'sp4_r_v_b_23')
// (14, 16, 'sp4_r_v_b_10')
// (15, 12, 'neigh_op_tnl_7')
// (15, 12, 'sp4_v_t_47')
// (15, 13, 'neigh_op_lft_7')
// (15, 13, 'sp4_v_b_47')
// (15, 14, 'neigh_op_bnl_7')
// (15, 14, 'sp4_v_b_34')
// (15, 15, 'sp4_v_b_23')
// (15, 16, 'sp4_h_r_4')
// (15, 16, 'sp4_v_b_10')
// (16, 16, 'sp4_h_r_17')
// (17, 16, 'sp4_h_r_28')
// (18, 13, 'sp4_r_v_b_41')
// (18, 14, 'sp4_r_v_b_28')
// (18, 15, 'sp4_r_v_b_17')
// (18, 16, 'sp4_h_r_41')
// (18, 16, 'sp4_r_v_b_4')
// (19, 12, 'sp4_v_t_41')
// (19, 13, 'sp4_v_b_41')
// (19, 14, 'sp4_v_b_28')
// (19, 15, 'local_g1_1')
// (19, 15, 'ram/WDATA_14')
// (19, 15, 'sp4_v_b_17')
// (19, 16, 'sp4_h_l_41')
// (19, 16, 'sp4_v_b_4')

reg n1956 = 0;
// (13, 12, 'sp4_r_v_b_47')
// (13, 13, 'sp4_r_v_b_34')
// (13, 14, 'local_g3_7')
// (13, 14, 'lutff_5/in_1')
// (13, 14, 'lutff_7/in_3')
// (13, 14, 'sp4_r_v_b_23')
// (13, 15, 'sp4_r_v_b_10')
// (13, 16, 'sp4_r_v_b_39')
// (13, 17, 'sp4_r_v_b_26')
// (13, 18, 'neigh_op_tnr_1')
// (13, 18, 'sp4_r_v_b_15')
// (13, 19, 'neigh_op_rgt_1')
// (13, 19, 'sp4_r_v_b_2')
// (13, 20, 'neigh_op_bnr_1')
// (14, 11, 'sp4_v_t_47')
// (14, 12, 'sp4_v_b_47')
// (14, 13, 'sp4_v_b_34')
// (14, 14, 'sp4_v_b_23')
// (14, 15, 'sp4_v_b_10')
// (14, 15, 'sp4_v_t_39')
// (14, 16, 'local_g3_7')
// (14, 16, 'lutff_1/in_3')
// (14, 16, 'sp4_v_b_39')
// (14, 17, 'sp4_v_b_26')
// (14, 18, 'neigh_op_top_1')
// (14, 18, 'sp4_v_b_15')
// (14, 19, 'local_g3_1')
// (14, 19, 'lutff_1/in_1')
// (14, 19, 'lutff_1/out')
// (14, 19, 'sp4_v_b_2')
// (14, 20, 'neigh_op_bot_1')
// (15, 18, 'neigh_op_tnl_1')
// (15, 19, 'neigh_op_lft_1')
// (15, 20, 'neigh_op_bnl_1')

wire n1957;
// (13, 13, 'local_g2_3')
// (13, 13, 'lutff_0/in_3')
// (13, 13, 'lutff_2/in_1')
// (13, 13, 'neigh_op_tnr_3')
// (13, 14, 'local_g3_3')
// (13, 14, 'lutff_2/in_2')
// (13, 14, 'neigh_op_rgt_3')
// (13, 15, 'neigh_op_bnr_3')
// (14, 13, 'neigh_op_top_3')
// (14, 14, 'lutff_3/out')
// (14, 15, 'neigh_op_bot_3')
// (15, 13, 'neigh_op_tnl_3')
// (15, 14, 'neigh_op_lft_3')
// (15, 15, 'neigh_op_bnl_3')

wire n1958;
// (13, 13, 'local_g3_2')
// (13, 13, 'lutff_3/in_2')
// (13, 13, 'neigh_op_tnr_2')
// (13, 14, 'neigh_op_rgt_2')
// (13, 15, 'neigh_op_bnr_2')
// (14, 13, 'neigh_op_top_2')
// (14, 14, 'lutff_2/out')
// (14, 14, 'sp4_r_v_b_37')
// (14, 15, 'neigh_op_bot_2')
// (14, 15, 'sp4_r_v_b_24')
// (14, 16, 'sp4_r_v_b_13')
// (14, 17, 'sp4_r_v_b_0')
// (15, 13, 'neigh_op_tnl_2')
// (15, 13, 'sp4_v_t_37')
// (15, 14, 'neigh_op_lft_2')
// (15, 14, 'sp4_v_b_37')
// (15, 15, 'neigh_op_bnl_2')
// (15, 15, 'sp4_v_b_24')
// (15, 16, 'sp4_v_b_13')
// (15, 17, 'sp4_h_r_0')
// (15, 17, 'sp4_v_b_0')
// (16, 17, 'sp4_h_r_13')
// (17, 17, 'sp4_h_r_24')
// (18, 14, 'sp4_r_v_b_37')
// (18, 15, 'sp4_r_v_b_24')
// (18, 16, 'sp4_r_v_b_13')
// (18, 17, 'sp4_h_r_37')
// (18, 17, 'sp4_r_v_b_0')
// (19, 13, 'sp4_v_t_37')
// (19, 14, 'sp4_v_b_37')
// (19, 15, 'sp4_v_b_24')
// (19, 16, 'local_g1_5')
// (19, 16, 'ram/WDATA_4')
// (19, 16, 'sp4_v_b_13')
// (19, 17, 'sp4_h_l_37')
// (19, 17, 'sp4_v_b_0')

wire n1959;
// (13, 13, 'neigh_op_tnr_0')
// (13, 14, 'neigh_op_rgt_0')
// (13, 15, 'neigh_op_bnr_0')
// (14, 13, 'neigh_op_top_0')
// (14, 14, 'local_g0_0')
// (14, 14, 'lutff_0/out')
// (14, 14, 'lutff_7/in_1')
// (14, 15, 'neigh_op_bot_0')
// (15, 13, 'neigh_op_tnl_0')
// (15, 14, 'neigh_op_lft_0')
// (15, 15, 'neigh_op_bnl_0')

wire n1960;
// (13, 13, 'neigh_op_tnr_1')
// (13, 14, 'local_g3_1')
// (13, 14, 'lutff_4/in_0')
// (13, 14, 'neigh_op_rgt_1')
// (13, 15, 'neigh_op_bnr_1')
// (14, 13, 'neigh_op_top_1')
// (14, 14, 'lutff_1/out')
// (14, 15, 'neigh_op_bot_1')
// (15, 13, 'neigh_op_tnl_1')
// (15, 14, 'neigh_op_lft_1')
// (15, 15, 'neigh_op_bnl_1')

wire n1961;
// (13, 13, 'neigh_op_tnr_4')
// (13, 14, 'neigh_op_rgt_4')
// (13, 15, 'neigh_op_bnr_4')
// (14, 13, 'neigh_op_top_4')
// (14, 14, 'local_g3_4')
// (14, 14, 'lutff_2/in_1')
// (14, 14, 'lutff_4/out')
// (14, 15, 'neigh_op_bot_4')
// (15, 13, 'neigh_op_tnl_4')
// (15, 14, 'neigh_op_lft_4')
// (15, 15, 'neigh_op_bnl_4')

wire n1962;
// (13, 13, 'neigh_op_tnr_5')
// (13, 14, 'neigh_op_rgt_5')
// (13, 15, 'neigh_op_bnr_5')
// (14, 13, 'neigh_op_top_5')
// (14, 14, 'local_g3_5')
// (14, 14, 'lutff_4/in_2')
// (14, 14, 'lutff_5/out')
// (14, 15, 'neigh_op_bot_5')
// (15, 13, 'neigh_op_tnl_5')
// (15, 14, 'neigh_op_lft_5')
// (15, 15, 'neigh_op_bnl_5')

wire n1963;
// (13, 13, 'neigh_op_tnr_6')
// (13, 14, 'neigh_op_rgt_6')
// (13, 15, 'neigh_op_bnr_6')
// (14, 13, 'neigh_op_top_6')
// (14, 14, 'local_g2_6')
// (14, 14, 'lutff_1/in_3')
// (14, 14, 'lutff_6/out')
// (14, 15, 'neigh_op_bot_6')
// (15, 13, 'neigh_op_tnl_6')
// (15, 14, 'neigh_op_lft_6')
// (15, 15, 'neigh_op_bnl_6')

wire n1964;
// (13, 13, 'neigh_op_tnr_7')
// (13, 14, 'neigh_op_rgt_7')
// (13, 15, 'local_g0_7')
// (13, 15, 'lutff_7/in_0')
// (13, 15, 'neigh_op_bnr_7')
// (14, 13, 'neigh_op_top_7')
// (14, 13, 'sp4_r_v_b_42')
// (14, 14, 'lutff_7/out')
// (14, 14, 'sp4_r_v_b_31')
// (14, 15, 'neigh_op_bot_7')
// (14, 15, 'sp4_r_v_b_18')
// (14, 16, 'sp4_r_v_b_7')
// (15, 12, 'sp4_v_t_42')
// (15, 13, 'neigh_op_tnl_7')
// (15, 13, 'sp4_v_b_42')
// (15, 14, 'neigh_op_lft_7')
// (15, 14, 'sp4_v_b_31')
// (15, 15, 'neigh_op_bnl_7')
// (15, 15, 'sp4_v_b_18')
// (15, 16, 'sp4_h_r_7')
// (15, 16, 'sp4_v_b_7')
// (16, 16, 'sp4_h_r_18')
// (17, 16, 'sp4_h_r_31')
// (18, 16, 'sp4_h_r_42')
// (19, 16, 'local_g0_2')
// (19, 16, 'ram/WDATA_6')
// (19, 16, 'sp4_h_l_42')
// (19, 16, 'sp4_h_r_10')
// (20, 16, 'sp4_h_r_23')
// (21, 16, 'sp4_h_r_34')
// (22, 16, 'sp4_h_r_47')
// (23, 16, 'sp4_h_l_47')

reg n1965 = 0;
// (13, 13, 'sp4_h_r_6')
// (14, 7, 'sp4_r_v_b_43')
// (14, 8, 'sp4_r_v_b_30')
// (14, 9, 'local_g3_3')
// (14, 9, 'lutff_7/in_3')
// (14, 9, 'sp4_r_v_b_19')
// (14, 10, 'sp4_r_v_b_6')
// (14, 11, 'sp4_r_v_b_38')
// (14, 12, 'neigh_op_tnr_7')
// (14, 12, 'sp4_r_v_b_27')
// (14, 13, 'neigh_op_rgt_7')
// (14, 13, 'sp4_h_r_19')
// (14, 13, 'sp4_h_r_3')
// (14, 13, 'sp4_r_v_b_14')
// (14, 14, 'neigh_op_bnr_7')
// (14, 14, 'sp4_r_v_b_3')
// (15, 6, 'sp4_v_t_43')
// (15, 7, 'sp4_v_b_43')
// (15, 8, 'local_g3_6')
// (15, 8, 'lutff_1/in_2')
// (15, 8, 'sp4_v_b_30')
// (15, 9, 'sp4_v_b_19')
// (15, 10, 'sp4_h_r_8')
// (15, 10, 'sp4_v_b_6')
// (15, 10, 'sp4_v_t_38')
// (15, 11, 'sp4_v_b_38')
// (15, 12, 'neigh_op_top_7')
// (15, 12, 'sp4_v_b_27')
// (15, 13, 'lutff_7/out')
// (15, 13, 'sp4_h_r_14')
// (15, 13, 'sp4_h_r_30')
// (15, 13, 'sp4_v_b_14')
// (15, 14, 'neigh_op_bot_7')
// (15, 14, 'sp4_v_b_3')
// (16, 6, 'sp4_r_v_b_45')
// (16, 7, 'sp4_r_v_b_32')
// (16, 8, 'sp4_r_v_b_21')
// (16, 9, 'sp4_r_v_b_8')
// (16, 10, 'sp4_h_r_21')
// (16, 10, 'sp4_r_v_b_37')
// (16, 11, 'sp4_r_v_b_24')
// (16, 12, 'neigh_op_tnl_7')
// (16, 12, 'sp4_r_v_b_13')
// (16, 13, 'local_g1_7')
// (16, 13, 'lutff_4/in_0')
// (16, 13, 'neigh_op_lft_7')
// (16, 13, 'sp4_h_r_27')
// (16, 13, 'sp4_h_r_43')
// (16, 13, 'sp4_r_v_b_0')
// (16, 14, 'neigh_op_bnl_7')
// (17, 5, 'sp4_v_t_45')
// (17, 6, 'sp4_r_v_b_44')
// (17, 6, 'sp4_v_b_45')
// (17, 7, 'sp4_r_v_b_33')
// (17, 7, 'sp4_v_b_32')
// (17, 8, 'local_g0_5')
// (17, 8, 'lutff_1/in_0')
// (17, 8, 'sp4_r_v_b_20')
// (17, 8, 'sp4_v_b_21')
// (17, 9, 'sp4_h_r_0')
// (17, 9, 'sp4_r_v_b_9')
// (17, 9, 'sp4_v_b_8')
// (17, 9, 'sp4_v_t_37')
// (17, 10, 'sp4_h_r_32')
// (17, 10, 'sp4_r_v_b_44')
// (17, 10, 'sp4_v_b_37')
// (17, 11, 'sp4_r_v_b_33')
// (17, 11, 'sp4_v_b_24')
// (17, 12, 'sp4_r_v_b_20')
// (17, 12, 'sp4_v_b_13')
// (17, 13, 'sp4_h_l_43')
// (17, 13, 'sp4_h_r_2')
// (17, 13, 'sp4_h_r_38')
// (17, 13, 'sp4_r_v_b_9')
// (17, 13, 'sp4_v_b_0')
// (18, 5, 'sp4_v_t_44')
// (18, 6, 'sp4_v_b_44')
// (18, 7, 'sp4_v_b_33')
// (18, 8, 'local_g0_4')
// (18, 8, 'lutff_5/in_3')
// (18, 8, 'sp4_v_b_20')
// (18, 9, 'local_g0_1')
// (18, 9, 'lutff_5/in_0')
// (18, 9, 'sp4_h_r_13')
// (18, 9, 'sp4_h_r_9')
// (18, 9, 'sp4_v_b_9')
// (18, 9, 'sp4_v_t_44')
// (18, 10, 'sp4_h_r_45')
// (18, 10, 'sp4_v_b_44')
// (18, 11, 'sp4_v_b_33')
// (18, 12, 'sp4_v_b_20')
// (18, 13, 'sp4_h_l_38')
// (18, 13, 'sp4_h_r_15')
// (18, 13, 'sp4_v_b_9')
// (19, 9, 'sp4_h_r_20')
// (19, 9, 'sp4_h_r_24')
// (19, 10, 'sp4_h_l_45')
// (19, 10, 'sp4_h_r_8')
// (19, 13, 'sp4_h_r_26')
// (20, 9, 'local_g3_5')
// (20, 9, 'lutff_6/in_2')
// (20, 9, 'sp4_h_r_33')
// (20, 9, 'sp4_h_r_37')
// (20, 10, 'local_g0_5')
// (20, 10, 'lutff_3/in_2')
// (20, 10, 'sp4_h_r_21')
// (20, 10, 'sp4_r_v_b_39')
// (20, 11, 'sp4_r_v_b_26')
// (20, 12, 'sp4_r_v_b_15')
// (20, 13, 'sp4_h_r_39')
// (20, 13, 'sp4_r_v_b_2')
// (21, 9, 'sp4_h_l_37')
// (21, 9, 'sp4_h_r_44')
// (21, 9, 'sp4_v_t_39')
// (21, 10, 'sp4_h_r_32')
// (21, 10, 'sp4_v_b_39')
// (21, 11, 'local_g2_2')
// (21, 11, 'lutff_4/in_2')
// (21, 11, 'sp4_v_b_26')
// (21, 12, 'sp4_v_b_15')
// (21, 13, 'sp4_h_l_39')
// (21, 13, 'sp4_v_b_2')
// (22, 9, 'sp4_h_l_44')
// (22, 10, 'sp4_h_r_45')
// (23, 10, 'sp4_h_l_45')

reg n1966 = 0;
// (13, 13, 'sp4_r_v_b_43')
// (13, 14, 'sp4_r_v_b_30')
// (13, 15, 'sp4_r_v_b_19')
// (13, 16, 'sp4_r_v_b_6')
// (13, 17, 'sp4_r_v_b_38')
// (13, 18, 'neigh_op_tnr_7')
// (13, 18, 'sp4_r_v_b_27')
// (13, 19, 'neigh_op_rgt_7')
// (13, 19, 'sp4_r_v_b_14')
// (13, 20, 'neigh_op_bnr_7')
// (13, 20, 'sp4_r_v_b_3')
// (14, 12, 'sp4_v_t_43')
// (14, 13, 'sp4_v_b_43')
// (14, 14, 'sp4_v_b_30')
// (14, 15, 'local_g0_3')
// (14, 15, 'lutff_0/in_3')
// (14, 15, 'lutff_1/in_0')
// (14, 15, 'sp4_v_b_19')
// (14, 16, 'local_g1_3')
// (14, 16, 'lutff_7/in_3')
// (14, 16, 'sp4_h_r_3')
// (14, 16, 'sp4_v_b_6')
// (14, 16, 'sp4_v_t_38')
// (14, 17, 'sp4_v_b_38')
// (14, 18, 'neigh_op_top_7')
// (14, 18, 'sp4_v_b_27')
// (14, 19, 'local_g2_7')
// (14, 19, 'lutff_0/in_1')
// (14, 19, 'lutff_7/in_0')
// (14, 19, 'lutff_7/out')
// (14, 19, 'sp4_v_b_14')
// (14, 20, 'neigh_op_bot_7')
// (14, 20, 'sp4_v_b_3')
// (15, 16, 'sp4_h_r_14')
// (15, 18, 'neigh_op_tnl_7')
// (15, 19, 'neigh_op_lft_7')
// (15, 20, 'neigh_op_bnl_7')
// (16, 16, 'sp4_h_r_27')
// (17, 16, 'sp4_h_r_38')
// (18, 16, 'sp4_h_l_38')

wire n1967;
// (13, 13, 'sp4_r_v_b_47')
// (13, 14, 'sp4_r_v_b_34')
// (13, 14, 'sp4_r_v_b_47')
// (13, 15, 'sp4_r_v_b_23')
// (13, 15, 'sp4_r_v_b_34')
// (13, 16, 'neigh_op_tnr_5')
// (13, 16, 'sp4_r_v_b_10')
// (13, 16, 'sp4_r_v_b_23')
// (13, 17, 'neigh_op_rgt_5')
// (13, 17, 'sp4_r_v_b_10')
// (13, 17, 'sp4_r_v_b_42')
// (13, 18, 'local_g3_3')
// (13, 18, 'lutff_global/cen')
// (13, 18, 'neigh_op_bnr_5')
// (13, 18, 'sp4_r_v_b_31')
// (13, 18, 'sp4_r_v_b_41')
// (13, 18, 'sp4_r_v_b_43')
// (13, 19, 'sp4_r_v_b_18')
// (13, 19, 'sp4_r_v_b_28')
// (13, 19, 'sp4_r_v_b_30')
// (13, 20, 'sp4_r_v_b_17')
// (13, 20, 'sp4_r_v_b_19')
// (13, 20, 'sp4_r_v_b_7')
// (13, 21, 'local_g1_4')
// (13, 21, 'lutff_0/in_1')
// (13, 21, 'sp4_r_v_b_4')
// (13, 21, 'sp4_r_v_b_6')
// (14, 12, 'sp4_v_t_47')
// (14, 13, 'sp4_v_b_47')
// (14, 13, 'sp4_v_t_47')
// (14, 14, 'sp4_v_b_34')
// (14, 14, 'sp4_v_b_47')
// (14, 15, 'sp4_v_b_23')
// (14, 15, 'sp4_v_b_34')
// (14, 16, 'local_g0_2')
// (14, 16, 'lutff_global/cen')
// (14, 16, 'neigh_op_top_5')
// (14, 16, 'sp4_v_b_10')
// (14, 16, 'sp4_v_b_23')
// (14, 16, 'sp4_v_t_42')
// (14, 17, 'lutff_5/out')
// (14, 17, 'sp4_h_r_10')
// (14, 17, 'sp4_v_b_10')
// (14, 17, 'sp4_v_b_42')
// (14, 17, 'sp4_v_t_41')
// (14, 17, 'sp4_v_t_43')
// (14, 18, 'neigh_op_bot_5')
// (14, 18, 'sp4_v_b_31')
// (14, 18, 'sp4_v_b_41')
// (14, 18, 'sp4_v_b_43')
// (14, 19, 'sp4_v_b_18')
// (14, 19, 'sp4_v_b_28')
// (14, 19, 'sp4_v_b_30')
// (14, 20, 'sp4_v_b_17')
// (14, 20, 'sp4_v_b_19')
// (14, 20, 'sp4_v_b_7')
// (14, 21, 'sp4_v_b_4')
// (14, 21, 'sp4_v_b_6')
// (15, 16, 'neigh_op_tnl_5')
// (15, 17, 'neigh_op_lft_5')
// (15, 17, 'sp4_h_r_23')
// (15, 18, 'neigh_op_bnl_5')
// (16, 17, 'sp4_h_r_34')
// (17, 17, 'sp4_h_r_47')
// (18, 17, 'sp4_h_l_47')

wire n1968;
// (13, 14, 'neigh_op_tnr_0')
// (13, 15, 'neigh_op_rgt_0')
// (13, 16, 'neigh_op_bnr_0')
// (14, 14, 'neigh_op_top_0')
// (14, 15, 'local_g0_0')
// (14, 15, 'lutff_0/out')
// (14, 15, 'lutff_5/in_1')
// (14, 15, 'sp4_h_r_0')
// (14, 16, 'local_g0_0')
// (14, 16, 'lutff_6/in_0')
// (14, 16, 'neigh_op_bot_0')
// (15, 14, 'neigh_op_tnl_0')
// (15, 15, 'neigh_op_lft_0')
// (15, 15, 'sp4_h_r_13')
// (15, 16, 'neigh_op_bnl_0')
// (16, 15, 'sp4_h_r_24')
// (17, 15, 'sp4_h_r_37')
// (18, 15, 'sp4_h_l_37')
// (18, 15, 'sp4_h_r_3')
// (19, 15, 'local_g1_6')
// (19, 15, 'ram/RADDR_0')
// (19, 15, 'sp4_h_r_14')
// (20, 15, 'sp4_h_r_27')
// (21, 15, 'sp4_h_r_38')
// (22, 15, 'sp4_h_l_38')

wire n1969;
// (13, 14, 'neigh_op_tnr_1')
// (13, 15, 'local_g2_1')
// (13, 15, 'lutff_1/in_2')
// (13, 15, 'neigh_op_rgt_1')
// (13, 16, 'neigh_op_bnr_1')
// (14, 14, 'neigh_op_top_1')
// (14, 15, 'lutff_1/out')
// (14, 16, 'neigh_op_bot_1')
// (15, 14, 'neigh_op_tnl_1')
// (15, 15, 'neigh_op_lft_1')
// (15, 16, 'neigh_op_bnl_1')

wire n1970;
// (13, 14, 'neigh_op_tnr_4')
// (13, 15, 'neigh_op_rgt_4')
// (13, 16, 'neigh_op_bnr_4')
// (14, 14, 'neigh_op_top_4')
// (14, 15, 'lutff_4/out')
// (14, 16, 'neigh_op_bot_4')
// (15, 14, 'local_g2_4')
// (15, 14, 'local_g3_4')
// (15, 14, 'lutff_1/in_2')
// (15, 14, 'lutff_global/s_r')
// (15, 14, 'neigh_op_tnl_4')
// (15, 15, 'neigh_op_lft_4')
// (15, 16, 'neigh_op_bnl_4')

wire n1971;
// (13, 14, 'neigh_op_tnr_5')
// (13, 15, 'local_g2_5')
// (13, 15, 'local_g3_5')
// (13, 15, 'lutff_0/in_1')
// (13, 15, 'lutff_1/in_3')
// (13, 15, 'neigh_op_rgt_5')
// (13, 16, 'neigh_op_bnr_5')
// (14, 14, 'neigh_op_top_5')
// (14, 15, 'lutff_5/out')
// (14, 16, 'neigh_op_bot_5')
// (15, 14, 'neigh_op_tnl_5')
// (15, 15, 'neigh_op_lft_5')
// (15, 16, 'neigh_op_bnl_5')

wire n1972;
// (13, 14, 'neigh_op_tnr_7')
// (13, 15, 'neigh_op_rgt_7')
// (13, 16, 'neigh_op_bnr_7')
// (14, 14, 'neigh_op_top_7')
// (14, 15, 'local_g3_7')
// (14, 15, 'lutff_2/in_0')
// (14, 15, 'lutff_7/out')
// (14, 16, 'neigh_op_bot_7')
// (15, 14, 'neigh_op_tnl_7')
// (15, 15, 'neigh_op_lft_7')
// (15, 16, 'neigh_op_bnl_7')

wire n1973;
// (13, 14, 'sp4_r_v_b_36')
// (13, 15, 'neigh_op_tnr_6')
// (13, 15, 'sp4_r_v_b_25')
// (13, 16, 'local_g2_4')
// (13, 16, 'lutff_global/s_r')
// (13, 16, 'neigh_op_rgt_6')
// (13, 16, 'sp4_r_v_b_12')
// (13, 17, 'neigh_op_bnr_6')
// (13, 17, 'sp4_r_v_b_1')
// (14, 13, 'sp4_v_t_36')
// (14, 14, 'sp4_v_b_36')
// (14, 15, 'neigh_op_top_6')
// (14, 15, 'sp4_v_b_25')
// (14, 16, 'lutff_6/out')
// (14, 16, 'sp4_v_b_12')
// (14, 17, 'neigh_op_bot_6')
// (14, 17, 'sp4_v_b_1')
// (15, 15, 'neigh_op_tnl_6')
// (15, 16, 'neigh_op_lft_6')
// (15, 17, 'neigh_op_bnl_6')

wire n1974;
// (13, 15, 'lutff_1/cout')
// (13, 15, 'lutff_2/in_3')

wire n1975;
// (13, 15, 'lutff_2/cout')
// (13, 15, 'lutff_3/in_3')

wire n1976;
// (13, 15, 'lutff_3/cout')
// (13, 15, 'lutff_4/in_3')

wire n1977;
// (13, 15, 'lutff_4/cout')
// (13, 15, 'lutff_5/in_3')

reg n1978 = 0;
// (13, 15, 'neigh_op_tnr_1')
// (13, 16, 'neigh_op_rgt_1')
// (13, 16, 'sp4_h_r_7')
// (13, 17, 'local_g0_1')
// (13, 17, 'lutff_1/in_2')
// (13, 17, 'neigh_op_bnr_1')
// (14, 15, 'local_g0_1')
// (14, 15, 'lutff_2/in_1')
// (14, 15, 'neigh_op_top_1')
// (14, 16, 'local_g2_1')
// (14, 16, 'lutff_1/in_2')
// (14, 16, 'lutff_1/out')
// (14, 16, 'sp4_h_r_18')
// (14, 17, 'neigh_op_bot_1')
// (15, 15, 'neigh_op_tnl_1')
// (15, 16, 'neigh_op_lft_1')
// (15, 16, 'sp4_h_r_31')
// (15, 17, 'neigh_op_bnl_1')
// (16, 16, 'sp4_h_r_42')
// (17, 16, 'sp4_h_l_42')
// (17, 16, 'sp4_h_r_7')
// (18, 16, 'sp4_h_r_18')
// (19, 16, 'local_g3_7')
// (19, 16, 'ram/WADDR_1')
// (19, 16, 'sp4_h_r_31')
// (20, 16, 'sp4_h_r_42')
// (21, 16, 'sp4_h_l_42')

wire n1979;
// (13, 15, 'neigh_op_tnr_3')
// (13, 16, 'neigh_op_rgt_3')
// (13, 17, 'neigh_op_bnr_3')
// (14, 15, 'neigh_op_top_3')
// (14, 16, 'lutff_3/out')
// (14, 17, 'neigh_op_bot_3')
// (15, 15, 'local_g2_3')
// (15, 15, 'lutff_2/in_1')
// (15, 15, 'neigh_op_tnl_3')
// (15, 16, 'neigh_op_lft_3')
// (15, 17, 'neigh_op_bnl_3')

reg n1980 = 0;
// (13, 15, 'neigh_op_tnr_7')
// (13, 16, 'neigh_op_rgt_7')
// (13, 16, 'sp4_h_r_3')
// (13, 17, 'local_g0_7')
// (13, 17, 'lutff_0/in_1')
// (13, 17, 'neigh_op_bnr_7')
// (14, 15, 'neigh_op_top_7')
// (14, 16, 'local_g1_7')
// (14, 16, 'local_g2_7')
// (14, 16, 'lutff_1/in_1')
// (14, 16, 'lutff_6/in_1')
// (14, 16, 'lutff_7/in_0')
// (14, 16, 'lutff_7/out')
// (14, 16, 'sp4_h_r_14')
// (14, 17, 'neigh_op_bot_7')
// (15, 15, 'neigh_op_tnl_7')
// (15, 16, 'neigh_op_lft_7')
// (15, 16, 'sp4_h_r_27')
// (15, 17, 'neigh_op_bnl_7')
// (16, 16, 'sp4_h_r_38')
// (17, 16, 'sp4_h_l_38')
// (17, 16, 'sp4_h_r_3')
// (18, 16, 'sp4_h_r_14')
// (19, 16, 'local_g2_3')
// (19, 16, 'ram/WADDR_0')
// (19, 16, 'sp4_h_r_27')
// (20, 16, 'sp4_h_r_38')
// (21, 16, 'sp4_h_l_38')

wire n1981;
// (13, 15, 'sp4_r_v_b_38')
// (13, 16, 'local_g0_3')
// (13, 16, 'lutff_4/in_1')
// (13, 16, 'sp4_r_v_b_27')
// (13, 17, 'sp4_r_v_b_14')
// (13, 18, 'sp4_r_v_b_3')
// (13, 19, 'sp4_r_v_b_38')
// (13, 20, 'neigh_op_tnr_7')
// (13, 20, 'sp4_r_v_b_27')
// (13, 21, 'local_g1_3')
// (13, 21, 'lutff_7/in_3')
// (13, 21, 'neigh_op_rgt_7')
// (13, 21, 'sp4_h_r_3')
// (13, 21, 'sp4_r_v_b_14')
// (13, 22, 'neigh_op_bnr_7')
// (13, 22, 'sp4_r_v_b_3')
// (14, 14, 'sp4_v_t_38')
// (14, 15, 'sp4_v_b_38')
// (14, 16, 'sp4_v_b_27')
// (14, 17, 'local_g0_6')
// (14, 17, 'lutff_5/in_1')
// (14, 17, 'sp4_v_b_14')
// (14, 18, 'sp4_v_b_3')
// (14, 18, 'sp4_v_t_38')
// (14, 19, 'sp4_r_v_b_39')
// (14, 19, 'sp4_v_b_38')
// (14, 20, 'neigh_op_top_7')
// (14, 20, 'sp4_r_v_b_26')
// (14, 20, 'sp4_v_b_27')
// (14, 21, 'lutff_7/out')
// (14, 21, 'sp4_h_r_14')
// (14, 21, 'sp4_r_v_b_15')
// (14, 21, 'sp4_v_b_14')
// (14, 22, 'neigh_op_bot_7')
// (14, 22, 'sp4_r_v_b_2')
// (14, 22, 'sp4_v_b_3')
// (15, 18, 'sp4_h_r_2')
// (15, 18, 'sp4_v_t_39')
// (15, 19, 'sp4_v_b_39')
// (15, 20, 'neigh_op_tnl_7')
// (15, 20, 'sp4_v_b_26')
// (15, 21, 'neigh_op_lft_7')
// (15, 21, 'sp4_h_r_27')
// (15, 21, 'sp4_v_b_15')
// (15, 22, 'neigh_op_bnl_7')
// (15, 22, 'sp4_v_b_2')
// (16, 18, 'sp4_h_r_15')
// (16, 21, 'sp4_h_r_38')
// (17, 18, 'sp4_h_r_26')
// (17, 21, 'sp4_h_l_38')
// (18, 15, 'sp4_r_v_b_39')
// (18, 16, 'sp4_r_v_b_26')
// (18, 17, 'sp4_r_v_b_15')
// (18, 18, 'sp4_h_r_39')
// (18, 18, 'sp4_r_v_b_2')
// (19, 14, 'sp4_v_t_39')
// (19, 15, 'sp4_v_b_39')
// (19, 16, 'local_g2_2')
// (19, 16, 'ram/WCLKE')
// (19, 16, 'sp4_v_b_26')
// (19, 17, 'sp4_v_b_15')
// (19, 18, 'sp4_h_l_39')
// (19, 18, 'sp4_v_b_2')

reg n1982 = 0;
// (13, 16, 'local_g3_1')
// (13, 16, 'lutff_6/in_2')
// (13, 16, 'lutff_7/in_3')
// (13, 16, 'sp4_r_v_b_41')
// (13, 17, 'sp4_r_v_b_28')
// (13, 18, 'local_g2_2')
// (13, 18, 'lutff_2/in_2')
// (13, 18, 'neigh_op_tnr_2')
// (13, 18, 'sp4_r_v_b_17')
// (13, 19, 'neigh_op_rgt_2')
// (13, 19, 'sp4_r_v_b_4')
// (13, 20, 'neigh_op_bnr_2')
// (14, 15, 'sp4_v_t_41')
// (14, 16, 'sp4_v_b_41')
// (14, 17, 'sp4_v_b_28')
// (14, 18, 'neigh_op_top_2')
// (14, 18, 'sp4_v_b_17')
// (14, 19, 'local_g1_2')
// (14, 19, 'lutff_2/in_1')
// (14, 19, 'lutff_2/out')
// (14, 19, 'sp4_v_b_4')
// (14, 20, 'neigh_op_bot_2')
// (15, 18, 'neigh_op_tnl_2')
// (15, 19, 'neigh_op_lft_2')
// (15, 20, 'neigh_op_bnl_2')

reg n1983 = 0;
// (13, 16, 'local_g3_3')
// (13, 16, 'lutff_0/in_0')
// (13, 16, 'lutff_1/in_1')
// (13, 16, 'sp4_r_v_b_43')
// (13, 17, 'sp4_r_v_b_30')
// (13, 18, 'local_g2_3')
// (13, 18, 'lutff_6/in_3')
// (13, 18, 'neigh_op_tnr_3')
// (13, 18, 'sp4_r_v_b_19')
// (13, 19, 'neigh_op_rgt_3')
// (13, 19, 'sp4_r_v_b_6')
// (13, 20, 'neigh_op_bnr_3')
// (14, 15, 'sp4_v_t_43')
// (14, 16, 'sp4_v_b_43')
// (14, 17, 'sp4_v_b_30')
// (14, 18, 'neigh_op_top_3')
// (14, 18, 'sp4_v_b_19')
// (14, 19, 'local_g1_3')
// (14, 19, 'lutff_3/in_1')
// (14, 19, 'lutff_3/out')
// (14, 19, 'sp4_v_b_6')
// (14, 20, 'neigh_op_bot_3')
// (15, 18, 'neigh_op_tnl_3')
// (15, 19, 'neigh_op_lft_3')
// (15, 20, 'neigh_op_bnl_3')

reg n1984 = 0;
// (13, 16, 'local_g3_5')
// (13, 16, 'lutff_3/in_3')
// (13, 16, 'lutff_5/in_3')
// (13, 16, 'sp4_r_v_b_45')
// (13, 17, 'sp4_r_v_b_32')
// (13, 18, 'local_g3_4')
// (13, 18, 'lutff_7/in_0')
// (13, 18, 'neigh_op_tnr_4')
// (13, 18, 'sp4_r_v_b_21')
// (13, 19, 'neigh_op_rgt_4')
// (13, 19, 'sp4_r_v_b_8')
// (13, 20, 'neigh_op_bnr_4')
// (14, 15, 'sp4_v_t_45')
// (14, 16, 'sp4_v_b_45')
// (14, 17, 'sp4_v_b_32')
// (14, 18, 'neigh_op_top_4')
// (14, 18, 'sp4_v_b_21')
// (14, 19, 'local_g2_4')
// (14, 19, 'lutff_4/in_2')
// (14, 19, 'lutff_4/out')
// (14, 19, 'sp4_v_b_8')
// (14, 20, 'neigh_op_bot_4')
// (15, 18, 'neigh_op_tnl_4')
// (15, 19, 'neigh_op_lft_4')
// (15, 20, 'neigh_op_bnl_4')

wire n1985;
// (13, 16, 'neigh_op_tnr_3')
// (13, 17, 'neigh_op_rgt_3')
// (13, 17, 'sp4_h_r_11')
// (13, 18, 'neigh_op_bnr_3')
// (14, 16, 'neigh_op_top_3')
// (14, 17, 'lutff_3/out')
// (14, 17, 'sp4_h_r_22')
// (14, 18, 'neigh_op_bot_3')
// (15, 16, 'neigh_op_tnl_3')
// (15, 17, 'neigh_op_lft_3')
// (15, 17, 'sp4_h_r_35')
// (15, 18, 'neigh_op_bnl_3')
// (16, 14, 'sp4_r_v_b_40')
// (16, 15, 'sp4_r_v_b_29')
// (16, 16, 'local_g3_0')
// (16, 16, 'lutff_0/in_1')
// (16, 16, 'sp4_r_v_b_16')
// (16, 17, 'sp4_h_r_46')
// (16, 17, 'sp4_r_v_b_5')
// (17, 13, 'sp4_v_t_40')
// (17, 14, 'sp4_v_b_40')
// (17, 15, 'sp4_v_b_29')
// (17, 16, 'sp4_v_b_16')
// (17, 17, 'sp4_h_l_46')
// (17, 17, 'sp4_v_b_5')

reg n1986 = 0;
// (13, 16, 'neigh_op_tnr_6')
// (13, 17, 'neigh_op_rgt_6')
// (13, 18, 'neigh_op_bnr_6')
// (14, 16, 'neigh_op_top_6')
// (14, 17, 'local_g2_6')
// (14, 17, 'lutff_3/in_1')
// (14, 17, 'lutff_6/out')
// (14, 18, 'neigh_op_bot_6')
// (15, 16, 'neigh_op_tnl_6')
// (15, 17, 'neigh_op_lft_6')
// (15, 18, 'neigh_op_bnl_6')

reg n1987 = 0;
// (13, 16, 'sp4_r_v_b_46')
// (13, 17, 'sp4_r_v_b_35')
// (13, 18, 'sp4_r_v_b_22')
// (13, 19, 'sp4_r_v_b_11')
// (14, 15, 'sp4_v_t_46')
// (14, 16, 'sp4_v_b_46')
// (14, 17, 'sp4_v_b_35')
// (14, 18, 'local_g0_6')
// (14, 18, 'lutff_5/in_1')
// (14, 18, 'sp4_v_b_22')
// (14, 19, 'sp4_h_r_6')
// (14, 19, 'sp4_v_b_11')
// (15, 18, 'neigh_op_tnr_7')
// (15, 19, 'local_g2_7')
// (15, 19, 'lutff_1/in_2')
// (15, 19, 'neigh_op_rgt_7')
// (15, 19, 'sp4_h_r_19')
// (15, 20, 'neigh_op_bnr_7')
// (16, 18, 'neigh_op_top_7')
// (16, 19, 'local_g0_7')
// (16, 19, 'local_g3_7')
// (16, 19, 'lutff_1/in_2')
// (16, 19, 'lutff_7/in_3')
// (16, 19, 'lutff_7/out')
// (16, 19, 'sp4_h_r_30')
// (16, 20, 'neigh_op_bot_7')
// (17, 18, 'neigh_op_tnl_7')
// (17, 19, 'neigh_op_lft_7')
// (17, 19, 'sp4_h_r_43')
// (17, 20, 'neigh_op_bnl_7')
// (18, 19, 'sp4_h_l_43')

wire n1988;
// (13, 17, 'lutff_1/cout')
// (13, 17, 'lutff_2/in_3')

wire n1989;
// (13, 17, 'lutff_3/cout')
// (13, 17, 'lutff_4/in_3')

wire n1990;
// (13, 17, 'lutff_5/cout')
// (13, 17, 'lutff_6/in_3')

wire n1991;
// (13, 17, 'lutff_7/cout')
// (13, 18, 'carry_in')
// (13, 18, 'carry_in_mux')
// (13, 18, 'lutff_0/in_3')

reg n1992 = 0;
// (13, 17, 'neigh_op_tnr_0')
// (13, 18, 'neigh_op_rgt_0')
// (13, 19, 'neigh_op_bnr_0')
// (14, 17, 'neigh_op_top_0')
// (14, 18, 'local_g2_0')
// (14, 18, 'local_g3_0')
// (14, 18, 'lutff_0/in_3')
// (14, 18, 'lutff_0/out')
// (14, 18, 'lutff_5/in_3')
// (14, 18, 'sp4_h_r_0')
// (14, 19, 'neigh_op_bot_0')
// (15, 17, 'neigh_op_tnl_0')
// (15, 18, 'local_g0_0')
// (15, 18, 'lutff_3/in_1')
// (15, 18, 'neigh_op_lft_0')
// (15, 18, 'sp4_h_r_13')
// (15, 19, 'neigh_op_bnl_0')
// (16, 18, 'local_g3_0')
// (16, 18, 'lutff_3/in_2')
// (16, 18, 'sp4_h_r_24')
// (17, 18, 'sp4_h_r_37')
// (18, 18, 'sp4_h_l_37')

reg n1993 = 0;
// (13, 17, 'neigh_op_tnr_1')
// (13, 18, 'neigh_op_rgt_1')
// (13, 19, 'neigh_op_bnr_1')
// (14, 17, 'neigh_op_top_1')
// (14, 18, 'local_g0_1')
// (14, 18, 'local_g3_1')
// (14, 18, 'lutff_1/in_3')
// (14, 18, 'lutff_1/out')
// (14, 18, 'lutff_5/in_2')
// (14, 18, 'sp4_h_r_2')
// (14, 19, 'neigh_op_bot_1')
// (15, 17, 'neigh_op_tnl_1')
// (15, 18, 'local_g1_1')
// (15, 18, 'lutff_5/in_1')
// (15, 18, 'neigh_op_lft_1')
// (15, 18, 'sp4_h_r_15')
// (15, 19, 'neigh_op_bnl_1')
// (16, 18, 'local_g2_2')
// (16, 18, 'lutff_5/in_1')
// (16, 18, 'sp4_h_r_26')
// (17, 18, 'sp4_h_r_39')
// (18, 18, 'sp4_h_l_39')

wire n1994;
// (13, 17, 'neigh_op_tnr_2')
// (13, 18, 'neigh_op_rgt_2')
// (13, 18, 'sp4_h_r_9')
// (13, 19, 'neigh_op_bnr_2')
// (14, 17, 'neigh_op_top_2')
// (14, 18, 'lutff_2/out')
// (14, 18, 'sp4_h_r_20')
// (14, 19, 'neigh_op_bot_2')
// (15, 17, 'neigh_op_tnl_2')
// (15, 18, 'neigh_op_lft_2')
// (15, 18, 'sp4_h_r_33')
// (15, 19, 'neigh_op_bnl_2')
// (16, 15, 'sp4_r_v_b_38')
// (16, 16, 'sp4_r_v_b_27')
// (16, 17, 'local_g2_6')
// (16, 17, 'lutff_0/in_0')
// (16, 17, 'lutff_3/in_1')
// (16, 17, 'sp4_r_v_b_14')
// (16, 18, 'sp4_h_r_44')
// (16, 18, 'sp4_r_v_b_3')
// (17, 14, 'sp4_v_t_38')
// (17, 15, 'sp4_v_b_38')
// (17, 16, 'sp4_v_b_27')
// (17, 17, 'sp4_v_b_14')
// (17, 18, 'sp4_h_l_44')
// (17, 18, 'sp4_v_b_3')

reg n1995 = 0;
// (13, 17, 'neigh_op_tnr_3')
// (13, 18, 'neigh_op_rgt_3')
// (13, 19, 'neigh_op_bnr_3')
// (14, 17, 'neigh_op_top_3')
// (14, 18, 'local_g2_3')
// (14, 18, 'lutff_3/in_0')
// (14, 18, 'lutff_3/out')
// (14, 18, 'lutff_5/in_0')
// (14, 18, 'sp4_h_r_6')
// (14, 19, 'neigh_op_bot_3')
// (15, 17, 'neigh_op_tnl_3')
// (15, 18, 'local_g1_3')
// (15, 18, 'lutff_7/in_1')
// (15, 18, 'neigh_op_lft_3')
// (15, 18, 'sp4_h_r_19')
// (15, 19, 'neigh_op_bnl_3')
// (16, 18, 'local_g3_6')
// (16, 18, 'lutff_7/in_2')
// (16, 18, 'sp4_h_r_30')
// (17, 18, 'sp4_h_r_43')
// (18, 18, 'sp4_h_l_43')

wire n1996;
// (13, 17, 'neigh_op_tnr_5')
// (13, 18, 'neigh_op_rgt_5')
// (13, 19, 'neigh_op_bnr_5')
// (14, 17, 'neigh_op_top_5')
// (14, 18, 'local_g2_5')
// (14, 18, 'lutff_2/in_1')
// (14, 18, 'lutff_5/out')
// (14, 19, 'neigh_op_bot_5')
// (15, 17, 'neigh_op_tnl_5')
// (15, 18, 'neigh_op_lft_5')
// (15, 19, 'neigh_op_bnl_5')

reg n1997 = 0;
// (13, 17, 'neigh_op_tnr_7')
// (13, 18, 'neigh_op_rgt_7')
// (13, 18, 'sp4_h_r_3')
// (13, 19, 'neigh_op_bnr_7')
// (14, 17, 'neigh_op_top_7')
// (14, 18, 'local_g3_7')
// (14, 18, 'lutff_2/in_2')
// (14, 18, 'lutff_7/in_1')
// (14, 18, 'lutff_7/out')
// (14, 18, 'sp4_h_r_14')
// (14, 19, 'neigh_op_bot_7')
// (15, 17, 'neigh_op_tnl_7')
// (15, 18, 'local_g0_7')
// (15, 18, 'lutff_0/in_1')
// (15, 18, 'neigh_op_lft_7')
// (15, 18, 'sp4_h_r_27')
// (15, 19, 'neigh_op_bnl_7')
// (16, 18, 'local_g2_6')
// (16, 18, 'lutff_0/in_2')
// (16, 18, 'lutff_1/in_3')
// (16, 18, 'sp4_h_r_38')
// (17, 18, 'sp4_h_l_38')

wire n1998;
// (13, 18, 'neigh_op_tnr_6')
// (13, 19, 'neigh_op_rgt_6')
// (13, 20, 'neigh_op_bnr_6')
// (14, 18, 'neigh_op_top_6')
// (14, 19, 'lutff_6/out')
// (14, 20, 'neigh_op_bot_6')
// (15, 18, 'neigh_op_tnl_6')
// (15, 19, 'local_g0_6')
// (15, 19, 'lutff_7/in_1')
// (15, 19, 'neigh_op_lft_6')
// (15, 20, 'local_g3_6')
// (15, 20, 'lutff_5/in_0')
// (15, 20, 'neigh_op_bnl_6')

wire n1999;
// (13, 18, 'sp4_h_r_1')
// (14, 18, 'local_g0_4')
// (14, 18, 'lutff_0/in_2')
// (14, 18, 'sp4_h_r_12')
// (15, 17, 'neigh_op_tnr_2')
// (15, 18, 'neigh_op_rgt_2')
// (15, 18, 'sp4_h_r_25')
// (15, 19, 'neigh_op_bnr_2')
// (16, 17, 'neigh_op_top_2')
// (16, 18, 'lutff_2/out')
// (16, 18, 'sp4_h_r_36')
// (16, 19, 'neigh_op_bot_2')
// (17, 17, 'neigh_op_tnl_2')
// (17, 18, 'neigh_op_lft_2')
// (17, 18, 'sp4_h_l_36')
// (17, 19, 'neigh_op_bnl_2')

wire n2000;
// (13, 18, 'sp4_h_r_5')
// (14, 18, 'local_g1_0')
// (14, 18, 'lutff_1/in_0')
// (14, 18, 'sp4_h_r_16')
// (15, 17, 'neigh_op_tnr_4')
// (15, 18, 'neigh_op_rgt_4')
// (15, 18, 'sp4_h_r_29')
// (15, 19, 'neigh_op_bnr_4')
// (16, 17, 'neigh_op_top_4')
// (16, 18, 'lutff_4/out')
// (16, 18, 'sp4_h_r_40')
// (16, 19, 'neigh_op_bot_4')
// (17, 17, 'neigh_op_tnl_4')
// (17, 18, 'neigh_op_lft_4')
// (17, 18, 'sp4_h_l_40')
// (17, 19, 'neigh_op_bnl_4')

wire n2001;
// (13, 19, 'lutff_1/cout')
// (13, 19, 'lutff_2/in_3')

wire n2002;
// (13, 19, 'lutff_2/cout')
// (13, 19, 'lutff_3/in_3')

wire n2003;
// (13, 19, 'lutff_3/cout')
// (13, 19, 'lutff_4/in_3')

wire n2004;
// (13, 19, 'lutff_4/cout')
// (13, 19, 'lutff_5/in_3')

wire n2005;
// (13, 19, 'lutff_5/cout')
// (13, 19, 'lutff_6/in_3')

reg n2006 = 0;
// (13, 19, 'neigh_op_tnr_0')
// (13, 20, 'neigh_op_rgt_0')
// (13, 21, 'neigh_op_bnr_0')
// (14, 19, 'local_g0_0')
// (14, 19, 'lutff_2/in_2')
// (14, 19, 'neigh_op_top_0')
// (14, 19, 'sp4_r_v_b_44')
// (14, 20, 'lutff_0/out')
// (14, 20, 'sp4_r_v_b_33')
// (14, 21, 'neigh_op_bot_0')
// (14, 21, 'sp4_r_v_b_20')
// (14, 22, 'local_g2_1')
// (14, 22, 'lutff_3/in_2')
// (14, 22, 'sp4_r_v_b_9')
// (15, 18, 'sp4_v_t_44')
// (15, 19, 'neigh_op_tnl_0')
// (15, 19, 'sp4_v_b_44')
// (15, 20, 'neigh_op_lft_0')
// (15, 20, 'sp4_v_b_33')
// (15, 21, 'neigh_op_bnl_0')
// (15, 21, 'sp4_v_b_20')
// (15, 22, 'sp4_v_b_9')

reg n2007 = 0;
// (13, 19, 'neigh_op_tnr_2')
// (13, 20, 'neigh_op_rgt_2')
// (13, 21, 'neigh_op_bnr_2')
// (14, 19, 'local_g0_2')
// (14, 19, 'lutff_0/in_2')
// (14, 19, 'lutff_7/in_3')
// (14, 19, 'neigh_op_top_2')
// (14, 20, 'lutff_2/out')
// (14, 21, 'local_g1_2')
// (14, 21, 'lutff_0/in_1')
// (14, 21, 'neigh_op_bot_2')
// (15, 19, 'neigh_op_tnl_2')
// (15, 20, 'neigh_op_lft_2')
// (15, 21, 'neigh_op_bnl_2')

reg n2008 = 0;
// (13, 19, 'neigh_op_tnr_3')
// (13, 20, 'neigh_op_rgt_3')
// (13, 20, 'sp4_r_v_b_38')
// (13, 21, 'neigh_op_bnr_3')
// (13, 21, 'sp4_r_v_b_27')
// (13, 22, 'sp4_r_v_b_14')
// (13, 23, 'sp4_r_v_b_3')
// (14, 19, 'local_g0_3')
// (14, 19, 'lutff_3/in_2')
// (14, 19, 'neigh_op_top_3')
// (14, 19, 'sp4_v_t_38')
// (14, 20, 'lutff_3/out')
// (14, 20, 'sp4_v_b_38')
// (14, 21, 'neigh_op_bot_3')
// (14, 21, 'sp4_v_b_27')
// (14, 22, 'local_g1_6')
// (14, 22, 'lutff_0/in_3')
// (14, 22, 'sp4_v_b_14')
// (14, 23, 'sp4_v_b_3')
// (15, 19, 'neigh_op_tnl_3')
// (15, 20, 'neigh_op_lft_3')
// (15, 21, 'neigh_op_bnl_3')

reg n2009 = 0;
// (13, 19, 'neigh_op_tnr_4')
// (13, 20, 'neigh_op_rgt_4')
// (13, 20, 'sp4_r_v_b_40')
// (13, 21, 'neigh_op_bnr_4')
// (13, 21, 'sp4_r_v_b_29')
// (13, 22, 'sp4_r_v_b_16')
// (13, 23, 'sp4_r_v_b_5')
// (14, 19, 'local_g1_4')
// (14, 19, 'lutff_1/in_2')
// (14, 19, 'neigh_op_top_4')
// (14, 19, 'sp4_v_t_40')
// (14, 20, 'lutff_4/out')
// (14, 20, 'sp4_v_b_40')
// (14, 21, 'neigh_op_bot_4')
// (14, 21, 'sp4_v_b_29')
// (14, 22, 'local_g1_0')
// (14, 22, 'lutff_4/in_3')
// (14, 22, 'sp4_v_b_16')
// (14, 23, 'sp4_v_b_5')
// (15, 19, 'neigh_op_tnl_4')
// (15, 20, 'neigh_op_lft_4')
// (15, 21, 'neigh_op_bnl_4')

reg n2010 = 0;
// (13, 19, 'sp4_h_r_2')
// (14, 18, 'neigh_op_tnr_5')
// (14, 19, 'neigh_op_rgt_5')
// (14, 19, 'sp4_h_r_15')
// (14, 20, 'neigh_op_bnr_5')
// (15, 18, 'neigh_op_top_5')
// (15, 19, 'lutff_5/out')
// (15, 19, 'sp4_h_r_26')
// (15, 20, 'neigh_op_bot_5')
// (16, 16, 'sp4_r_v_b_45')
// (16, 17, 'sp4_r_v_b_32')
// (16, 18, 'neigh_op_tnl_5')
// (16, 18, 'sp4_r_v_b_21')
// (16, 19, 'neigh_op_lft_5')
// (16, 19, 'sp4_h_r_39')
// (16, 19, 'sp4_r_v_b_8')
// (16, 20, 'neigh_op_bnl_5')
// (17, 15, 'sp4_v_t_45')
// (17, 16, 'sp4_v_b_45')
// (17, 17, 'sp4_v_b_32')
// (17, 18, 'local_g1_5')
// (17, 18, 'lutff_6/in_0')
// (17, 18, 'sp4_v_b_21')
// (17, 19, 'sp4_h_l_39')
// (17, 19, 'sp4_v_b_8')

wire n2011;
// (13, 19, 'sp4_h_r_6')
// (14, 18, 'neigh_op_tnr_7')
// (14, 19, 'neigh_op_rgt_7')
// (14, 19, 'sp4_h_r_19')
// (14, 20, 'neigh_op_bnr_7')
// (15, 17, 'sp4_r_v_b_39')
// (15, 18, 'neigh_op_top_7')
// (15, 18, 'sp4_r_v_b_26')
// (15, 18, 'sp4_r_v_b_42')
// (15, 19, 'lutff_7/out')
// (15, 19, 'sp4_h_r_30')
// (15, 19, 'sp4_r_v_b_15')
// (15, 19, 'sp4_r_v_b_31')
// (15, 20, 'neigh_op_bot_7')
// (15, 20, 'sp4_r_v_b_18')
// (15, 20, 'sp4_r_v_b_2')
// (15, 21, 'sp4_r_v_b_7')
// (16, 16, 'sp4_h_r_2')
// (16, 16, 'sp4_r_v_b_43')
// (16, 16, 'sp4_v_t_39')
// (16, 17, 'sp4_h_r_7')
// (16, 17, 'sp4_r_v_b_30')
// (16, 17, 'sp4_v_b_39')
// (16, 17, 'sp4_v_t_42')
// (16, 18, 'neigh_op_tnl_7')
// (16, 18, 'sp4_r_v_b_19')
// (16, 18, 'sp4_v_b_26')
// (16, 18, 'sp4_v_b_42')
// (16, 19, 'neigh_op_lft_7')
// (16, 19, 'sp4_h_r_43')
// (16, 19, 'sp4_r_v_b_6')
// (16, 19, 'sp4_v_b_15')
// (16, 19, 'sp4_v_b_31')
// (16, 20, 'neigh_op_bnl_7')
// (16, 20, 'sp4_v_b_18')
// (16, 20, 'sp4_v_b_2')
// (16, 21, 'sp4_v_b_7')
// (17, 15, 'sp4_v_t_43')
// (17, 16, 'sp4_h_r_15')
// (17, 16, 'sp4_v_b_43')
// (17, 17, 'local_g0_2')
// (17, 17, 'lutff_1/in_3')
// (17, 17, 'lutff_2/in_2')
// (17, 17, 'lutff_3/in_3')
// (17, 17, 'lutff_4/in_0')
// (17, 17, 'lutff_5/in_3')
// (17, 17, 'lutff_7/in_3')
// (17, 17, 'sp4_h_r_18')
// (17, 17, 'sp4_v_b_30')
// (17, 18, 'local_g1_3')
// (17, 18, 'lutff_global/cen')
// (17, 18, 'sp4_v_b_19')
// (17, 19, 'sp4_h_l_43')
// (17, 19, 'sp4_v_b_6')
// (18, 16, 'local_g2_2')
// (18, 16, 'lutff_global/cen')
// (18, 16, 'sp4_h_r_26')
// (18, 17, 'sp4_h_r_31')
// (19, 16, 'sp4_h_r_39')
// (19, 17, 'sp4_h_r_42')
// (20, 16, 'sp4_h_l_39')
// (20, 17, 'sp4_h_l_42')

wire n2012;
// (13, 20, 'local_g2_6')
// (13, 20, 'lutff_7/in_3')
// (13, 20, 'neigh_op_tnr_6')
// (13, 21, 'neigh_op_rgt_6')
// (13, 21, 'sp4_h_r_1')
// (13, 22, 'neigh_op_bnr_6')
// (14, 16, 'sp4_r_v_b_45')
// (14, 17, 'sp4_r_v_b_32')
// (14, 18, 'sp4_r_v_b_21')
// (14, 19, 'sp4_r_v_b_37')
// (14, 19, 'sp4_r_v_b_8')
// (14, 20, 'neigh_op_top_6')
// (14, 20, 'sp4_r_v_b_24')
// (14, 20, 'sp4_r_v_b_40')
// (14, 21, 'lutff_6/out')
// (14, 21, 'sp4_h_r_12')
// (14, 21, 'sp4_r_v_b_13')
// (14, 21, 'sp4_r_v_b_29')
// (14, 21, 'sp4_r_v_b_45')
// (14, 22, 'neigh_op_bot_6')
// (14, 22, 'sp4_r_v_b_0')
// (14, 22, 'sp4_r_v_b_16')
// (14, 22, 'sp4_r_v_b_32')
// (14, 23, 'sp4_r_v_b_21')
// (14, 23, 'sp4_r_v_b_5')
// (14, 24, 'sp4_r_v_b_8')
// (15, 15, 'sp4_h_r_8')
// (15, 15, 'sp4_v_t_45')
// (15, 16, 'sp4_v_b_45')
// (15, 17, 'sp4_v_b_32')
// (15, 18, 'sp4_h_r_0')
// (15, 18, 'sp4_v_b_21')
// (15, 18, 'sp4_v_t_37')
// (15, 19, 'local_g2_5')
// (15, 19, 'lutff_5/in_2')
// (15, 19, 'sp4_h_r_5')
// (15, 19, 'sp4_v_b_37')
// (15, 19, 'sp4_v_b_8')
// (15, 19, 'sp4_v_t_40')
// (15, 20, 'neigh_op_tnl_6')
// (15, 20, 'sp4_h_r_8')
// (15, 20, 'sp4_v_b_24')
// (15, 20, 'sp4_v_b_40')
// (15, 20, 'sp4_v_t_45')
// (15, 21, 'neigh_op_lft_6')
// (15, 21, 'sp4_h_r_25')
// (15, 21, 'sp4_v_b_13')
// (15, 21, 'sp4_v_b_29')
// (15, 21, 'sp4_v_b_45')
// (15, 22, 'local_g2_6')
// (15, 22, 'lutff_4/in_2')
// (15, 22, 'neigh_op_bnl_6')
// (15, 22, 'sp4_h_r_0')
// (15, 22, 'sp4_h_r_6')
// (15, 22, 'sp4_v_b_0')
// (15, 22, 'sp4_v_b_16')
// (15, 22, 'sp4_v_b_32')
// (15, 23, 'local_g1_5')
// (15, 23, 'lutff_1/in_3')
// (15, 23, 'sp4_h_r_11')
// (15, 23, 'sp4_v_b_21')
// (15, 23, 'sp4_v_b_5')
// (15, 24, 'sp4_h_r_2')
// (15, 24, 'sp4_v_b_8')
// (16, 15, 'sp4_h_r_21')
// (16, 18, 'sp4_h_r_13')
// (16, 18, 'sp4_r_v_b_42')
// (16, 19, 'sp4_h_r_16')
// (16, 19, 'sp4_r_v_b_31')
// (16, 20, 'local_g3_2')
// (16, 20, 'lutff_4/in_3')
// (16, 20, 'sp4_h_r_21')
// (16, 20, 'sp4_r_v_b_18')
// (16, 21, 'local_g3_4')
// (16, 21, 'lutff_6/in_3')
// (16, 21, 'sp4_h_r_36')
// (16, 21, 'sp4_r_v_b_7')
// (16, 22, 'local_g1_5')
// (16, 22, 'lutff_6/in_0')
// (16, 22, 'sp4_h_r_13')
// (16, 22, 'sp4_h_r_19')
// (16, 23, 'local_g1_6')
// (16, 23, 'lutff_3/in_2')
// (16, 23, 'sp4_h_r_22')
// (16, 24, 'local_g0_7')
// (16, 24, 'lutff_7/in_0')
// (16, 24, 'sp4_h_r_15')
// (17, 15, 'sp4_h_r_32')
// (17, 17, 'sp4_h_r_0')
// (17, 17, 'sp4_v_t_42')
// (17, 18, 'sp4_h_r_24')
// (17, 18, 'sp4_v_b_42')
// (17, 19, 'sp4_h_r_29')
// (17, 19, 'sp4_v_b_31')
// (17, 20, 'sp4_h_r_32')
// (17, 20, 'sp4_v_b_18')
// (17, 21, 'local_g0_7')
// (17, 21, 'lutff_3/in_0')
// (17, 21, 'sp4_h_l_36')
// (17, 21, 'sp4_h_r_1')
// (17, 21, 'sp4_v_b_7')
// (17, 22, 'local_g3_6')
// (17, 22, 'lutff_1/in_2')
// (17, 22, 'sp4_h_r_24')
// (17, 22, 'sp4_h_r_30')
// (17, 23, 'local_g3_3')
// (17, 23, 'lutff_1/in_1')
// (17, 23, 'sp4_h_r_35')
// (17, 24, 'local_g3_2')
// (17, 24, 'lutff_2/in_1')
// (17, 24, 'sp4_h_r_26')
// (18, 15, 'local_g2_5')
// (18, 15, 'lutff_2/in_1')
// (18, 15, 'sp4_h_r_45')
// (18, 15, 'sp4_r_v_b_37')
// (18, 16, 'sp4_r_v_b_24')
// (18, 16, 'sp4_r_v_b_40')
// (18, 17, 'local_g2_5')
// (18, 17, 'lutff_0/in_3')
// (18, 17, 'sp4_h_r_13')
// (18, 17, 'sp4_r_v_b_13')
// (18, 17, 'sp4_r_v_b_29')
// (18, 18, 'local_g3_5')
// (18, 18, 'lutff_0/in_0')
// (18, 18, 'sp4_h_r_37')
// (18, 18, 'sp4_r_v_b_0')
// (18, 18, 'sp4_r_v_b_16')
// (18, 19, 'local_g3_0')
// (18, 19, 'lutff_0/in_3')
// (18, 19, 'sp4_h_r_40')
// (18, 19, 'sp4_r_v_b_5')
// (18, 20, 'local_g2_5')
// (18, 20, 'lutff_3/in_0')
// (18, 20, 'sp4_h_r_45')
// (18, 21, 'local_g1_4')
// (18, 21, 'lutff_7/in_0')
// (18, 21, 'sp4_h_r_12')
// (18, 22, 'local_g2_3')
// (18, 22, 'lutff_3/in_2')
// (18, 22, 'sp4_h_r_37')
// (18, 22, 'sp4_h_r_43')
// (18, 23, 'local_g2_6')
// (18, 23, 'lutff_1/in_3')
// (18, 23, 'sp4_h_r_46')
// (18, 24, 'local_g3_7')
// (18, 24, 'lutff_3/in_1')
// (18, 24, 'sp4_h_r_39')
// (19, 14, 'sp4_v_t_37')
// (19, 15, 'sp4_h_l_45')
// (19, 15, 'sp4_h_r_10')
// (19, 15, 'sp4_v_b_37')
// (19, 15, 'sp4_v_t_40')
// (19, 16, 'sp4_v_b_24')
// (19, 16, 'sp4_v_b_40')
// (19, 17, 'sp4_h_r_24')
// (19, 17, 'sp4_v_b_13')
// (19, 17, 'sp4_v_b_29')
// (19, 18, 'sp4_h_l_37')
// (19, 18, 'sp4_h_r_0')
// (19, 18, 'sp4_v_b_0')
// (19, 18, 'sp4_v_b_16')
// (19, 19, 'sp4_h_l_40')
// (19, 19, 'sp4_h_r_5')
// (19, 19, 'sp4_v_b_5')
// (19, 20, 'sp4_h_l_45')
// (19, 20, 'sp4_h_r_4')
// (19, 20, 'sp4_h_r_8')
// (19, 21, 'sp4_h_r_25')
// (19, 22, 'sp4_h_l_37')
// (19, 22, 'sp4_h_l_43')
// (19, 22, 'sp4_h_r_8')
// (19, 23, 'sp4_h_l_46')
// (19, 23, 'sp4_h_r_11')
// (19, 23, 'sp4_h_r_2')
// (19, 24, 'sp4_h_l_39')
// (19, 24, 'sp4_h_r_5')
// (20, 14, 'sp4_r_v_b_42')
// (20, 14, 'sp4_r_v_b_43')
// (20, 15, 'local_g1_7')
// (20, 15, 'lutff_1/in_3')
// (20, 15, 'sp4_h_r_23')
// (20, 15, 'sp4_r_v_b_30')
// (20, 15, 'sp4_r_v_b_31')
// (20, 16, 'local_g3_3')
// (20, 16, 'lutff_3/in_1')
// (20, 16, 'sp4_r_v_b_18')
// (20, 16, 'sp4_r_v_b_19')
// (20, 17, 'local_g3_5')
// (20, 17, 'lutff_4/in_0')
// (20, 17, 'sp4_h_r_37')
// (20, 17, 'sp4_r_v_b_6')
// (20, 17, 'sp4_r_v_b_7')
// (20, 18, 'local_g0_5')
// (20, 18, 'lutff_2/in_1')
// (20, 18, 'sp4_h_r_13')
// (20, 18, 'sp4_r_v_b_42')
// (20, 19, 'local_g1_0')
// (20, 19, 'lutff_6/in_3')
// (20, 19, 'sp4_h_r_16')
// (20, 19, 'sp4_r_v_b_31')
// (20, 20, 'local_g1_1')
// (20, 20, 'lutff_2/in_2')
// (20, 20, 'sp4_h_r_17')
// (20, 20, 'sp4_h_r_21')
// (20, 20, 'sp4_r_v_b_18')
// (20, 21, 'local_g3_4')
// (20, 21, 'lutff_2/in_1')
// (20, 21, 'sp4_h_r_36')
// (20, 21, 'sp4_r_v_b_7')
// (20, 22, 'local_g1_5')
// (20, 22, 'lutff_0/in_0')
// (20, 22, 'sp4_h_r_21')
// (20, 23, 'local_g1_6')
// (20, 23, 'lutff_4/in_3')
// (20, 23, 'sp4_h_r_15')
// (20, 23, 'sp4_h_r_22')
// (20, 24, 'sp4_h_r_16')
// (21, 13, 'sp4_v_t_42')
// (21, 13, 'sp4_v_t_43')
// (21, 14, 'sp4_v_b_42')
// (21, 14, 'sp4_v_b_43')
// (21, 15, 'local_g2_6')
// (21, 15, 'lutff_3/in_1')
// (21, 15, 'sp4_h_r_34')
// (21, 15, 'sp4_v_b_30')
// (21, 15, 'sp4_v_b_31')
// (21, 16, 'local_g1_2')
// (21, 16, 'lutff_7/in_0')
// (21, 16, 'sp4_v_b_18')
// (21, 16, 'sp4_v_b_19')
// (21, 17, 'local_g0_7')
// (21, 17, 'lutff_7/in_0')
// (21, 17, 'sp4_h_l_37')
// (21, 17, 'sp4_h_r_3')
// (21, 17, 'sp4_v_b_6')
// (21, 17, 'sp4_v_b_7')
// (21, 17, 'sp4_v_t_42')
// (21, 18, 'local_g3_0')
// (21, 18, 'lutff_0/in_3')
// (21, 18, 'sp4_h_r_24')
// (21, 18, 'sp4_v_b_42')
// (21, 19, 'local_g2_7')
// (21, 19, 'lutff_4/in_1')
// (21, 19, 'sp4_h_r_29')
// (21, 19, 'sp4_v_b_31')
// (21, 20, 'local_g1_2')
// (21, 20, 'lutff_6/in_3')
// (21, 20, 'sp4_h_r_28')
// (21, 20, 'sp4_h_r_32')
// (21, 20, 'sp4_v_b_18')
// (21, 21, 'local_g0_4')
// (21, 21, 'lutff_0/in_2')
// (21, 21, 'sp4_h_l_36')
// (21, 21, 'sp4_h_r_4')
// (21, 21, 'sp4_v_b_7')
// (21, 22, 'local_g2_0')
// (21, 22, 'lutff_3/in_3')
// (21, 22, 'sp4_h_r_32')
// (21, 23, 'local_g3_2')
// (21, 23, 'lutff_1/in_0')
// (21, 23, 'sp4_h_r_26')
// (21, 23, 'sp4_h_r_35')
// (21, 24, 'local_g3_5')
// (21, 24, 'lutff_6/in_0')
// (21, 24, 'sp4_h_r_29')
// (22, 15, 'sp4_h_r_47')
// (22, 15, 'sp4_r_v_b_43')
// (22, 16, 'local_g1_6')
// (22, 16, 'lutff_3/in_2')
// (22, 16, 'sp4_r_v_b_30')
// (22, 16, 'sp4_r_v_b_40')
// (22, 17, 'local_g3_3')
// (22, 17, 'lutff_2/in_0')
// (22, 17, 'sp4_h_r_14')
// (22, 17, 'sp4_r_v_b_19')
// (22, 17, 'sp4_r_v_b_29')
// (22, 18, 'local_g3_5')
// (22, 18, 'lutff_6/in_0')
// (22, 18, 'sp4_h_r_37')
// (22, 18, 'sp4_r_v_b_16')
// (22, 18, 'sp4_r_v_b_6')
// (22, 19, 'local_g2_0')
// (22, 19, 'lutff_1/in_1')
// (22, 19, 'sp4_h_r_40')
// (22, 19, 'sp4_r_v_b_5')
// (22, 20, 'local_g2_5')
// (22, 20, 'lutff_1/in_2')
// (22, 20, 'sp4_h_r_41')
// (22, 20, 'sp4_h_r_45')
// (22, 21, 'local_g1_1')
// (22, 21, 'lutff_3/in_1')
// (22, 21, 'sp4_h_r_17')
// (22, 22, 'local_g2_5')
// (22, 22, 'lutff_4/in_3')
// (22, 22, 'sp4_h_r_45')
// (22, 23, 'local_g2_6')
// (22, 23, 'lutff_6/in_2')
// (22, 23, 'sp4_h_r_39')
// (22, 23, 'sp4_h_r_46')
// (22, 24, 'sp4_h_r_40')
// (23, 14, 'sp4_v_t_43')
// (23, 15, 'local_g3_3')
// (23, 15, 'lutff_6/in_2')
// (23, 15, 'sp4_h_l_47')
// (23, 15, 'sp4_h_r_10')
// (23, 15, 'sp4_v_b_43')
// (23, 15, 'sp4_v_t_40')
// (23, 16, 'local_g3_6')
// (23, 16, 'lutff_6/in_1')
// (23, 16, 'sp4_v_b_30')
// (23, 16, 'sp4_v_b_40')
// (23, 17, 'local_g3_3')
// (23, 17, 'lutff_0/in_0')
// (23, 17, 'sp4_h_r_27')
// (23, 17, 'sp4_v_b_19')
// (23, 17, 'sp4_v_b_29')
// (23, 18, 'local_g0_0')
// (23, 18, 'lutff_1/in_1')
// (23, 18, 'sp4_h_l_37')
// (23, 18, 'sp4_h_r_8')
// (23, 18, 'sp4_v_b_16')
// (23, 18, 'sp4_v_b_6')
// (23, 19, 'local_g0_5')
// (23, 19, 'lutff_3/in_2')
// (23, 19, 'sp4_h_l_40')
// (23, 19, 'sp4_h_r_5')
// (23, 19, 'sp4_v_b_5')
// (23, 20, 'local_g0_7')
// (23, 20, 'lutff_7/in_2')
// (23, 20, 'sp4_h_l_41')
// (23, 20, 'sp4_h_l_45')
// (23, 20, 'sp4_h_r_7')
// (23, 21, 'local_g3_4')
// (23, 21, 'lutff_4/in_3')
// (23, 21, 'sp4_h_r_28')
// (23, 22, 'local_g0_0')
// (23, 22, 'lutff_0/in_2')
// (23, 22, 'sp4_h_l_45')
// (23, 22, 'sp4_h_r_8')
// (23, 23, 'sp4_h_l_39')
// (23, 23, 'sp4_h_l_46')
// (23, 24, 'sp4_h_l_40')
// (24, 14, 'sp4_r_v_b_44')
// (24, 15, 'local_g0_7')
// (24, 15, 'lutff_1/in_2')
// (24, 15, 'sp4_h_r_23')
// (24, 15, 'sp4_r_v_b_33')
// (24, 16, 'local_g3_4')
// (24, 16, 'lutff_5/in_2')
// (24, 16, 'sp4_r_v_b_20')
// (24, 17, 'local_g3_6')
// (24, 17, 'lutff_3/in_0')
// (24, 17, 'sp4_h_r_38')
// (24, 17, 'sp4_r_v_b_9')
// (24, 18, 'local_g0_5')
// (24, 18, 'lutff_3/in_0')
// (24, 18, 'sp4_h_r_21')
// (24, 18, 'sp4_r_v_b_47')
// (24, 19, 'local_g1_0')
// (24, 19, 'lutff_0/in_1')
// (24, 19, 'sp4_h_r_16')
// (24, 19, 'sp4_r_v_b_34')
// (24, 20, 'local_g3_7')
// (24, 20, 'lutff_2/in_2')
// (24, 20, 'sp4_h_r_18')
// (24, 20, 'sp4_r_v_b_23')
// (24, 21, 'local_g3_1')
// (24, 21, 'lutff_1/in_3')
// (24, 21, 'sp4_h_r_41')
// (24, 21, 'sp4_r_v_b_10')
// (24, 22, 'sp4_h_r_21')
// (25, 13, 'sp4_v_t_44')
// (25, 14, 'sp4_v_b_44')
// (25, 15, 'sp4_h_r_34')
// (25, 15, 'sp4_v_b_33')
// (25, 16, 'sp4_v_b_20')
// (25, 17, 'sp4_h_l_38')
// (25, 17, 'sp4_v_b_9')
// (25, 17, 'sp4_v_t_47')
// (25, 18, 'sp4_h_r_32')
// (25, 18, 'sp4_v_b_47')
// (25, 19, 'sp4_h_r_29')
// (25, 19, 'sp4_v_b_34')
// (25, 20, 'sp4_h_r_31')
// (25, 20, 'sp4_v_b_23')
// (25, 21, 'sp4_h_l_41')
// (25, 21, 'sp4_v_b_10')
// (25, 22, 'sp4_h_r_32')

wire n2013;
// (13, 20, 'lutff_1/cout')
// (13, 20, 'lutff_2/in_3')

wire n2014;
// (13, 20, 'lutff_2/cout')
// (13, 20, 'lutff_3/in_3')

wire n2015;
// (13, 20, 'lutff_3/cout')
// (13, 20, 'lutff_4/in_3')

wire n2016;
// (13, 20, 'lutff_4/cout')
// (13, 20, 'lutff_5/in_3')

wire n2017;
// (13, 20, 'lutff_5/cout')
// (13, 20, 'lutff_6/in_3')

wire n2018;
// (13, 20, 'neigh_op_tnr_0')
// (13, 20, 'sp4_r_v_b_45')
// (13, 21, 'neigh_op_rgt_0')
// (13, 21, 'sp4_r_v_b_32')
// (13, 22, 'neigh_op_bnr_0')
// (13, 22, 'sp4_r_v_b_21')
// (13, 23, 'sp4_r_v_b_8')
// (14, 19, 'sp4_v_t_45')
// (14, 20, 'neigh_op_top_0')
// (14, 20, 'sp4_v_b_45')
// (14, 21, 'lutff_0/out')
// (14, 21, 'sp4_v_b_32')
// (14, 22, 'local_g0_0')
// (14, 22, 'lutff_6/in_0')
// (14, 22, 'neigh_op_bot_0')
// (14, 22, 'sp4_v_b_21')
// (14, 23, 'local_g0_0')
// (14, 23, 'lutff_0/in_2')
// (14, 23, 'sp4_v_b_8')
// (15, 20, 'neigh_op_tnl_0')
// (15, 21, 'neigh_op_lft_0')
// (15, 22, 'neigh_op_bnl_0')

reg n2019 = 0;
// (13, 20, 'neigh_op_tnr_1')
// (13, 21, 'neigh_op_rgt_1')
// (13, 22, 'neigh_op_bnr_1')
// (14, 20, 'neigh_op_top_1')
// (14, 21, 'local_g3_1')
// (14, 21, 'lutff_1/out')
// (14, 21, 'lutff_3/in_3')
// (14, 22, 'neigh_op_bot_1')
// (15, 20, 'neigh_op_tnl_1')
// (15, 21, 'neigh_op_lft_1')
// (15, 22, 'neigh_op_bnl_1')

wire n2020;
// (13, 20, 'neigh_op_tnr_3')
// (13, 21, 'neigh_op_rgt_3')
// (13, 22, 'neigh_op_bnr_3')
// (14, 20, 'neigh_op_top_3')
// (14, 21, 'local_g2_3')
// (14, 21, 'lutff_1/in_2')
// (14, 21, 'lutff_3/out')
// (14, 21, 'lutff_6/in_3')
// (14, 22, 'neigh_op_bot_3')
// (15, 20, 'neigh_op_tnl_3')
// (15, 21, 'neigh_op_lft_3')
// (15, 22, 'neigh_op_bnl_3')

reg n2021 = 0;
// (13, 20, 'neigh_op_tnr_5')
// (13, 21, 'local_g3_5')
// (13, 21, 'lutff_0/in_2')
// (13, 21, 'lutff_1/in_3')
// (13, 21, 'lutff_2/in_2')
// (13, 21, 'lutff_3/in_1')
// (13, 21, 'lutff_6/in_2')
// (13, 21, 'neigh_op_rgt_5')
// (13, 22, 'neigh_op_bnr_5')
// (14, 20, 'neigh_op_top_5')
// (14, 21, 'local_g1_5')
// (14, 21, 'lutff_1/in_3')
// (14, 21, 'lutff_5/out')
// (14, 22, 'neigh_op_bot_5')
// (15, 20, 'local_g3_5')
// (15, 20, 'lutff_0/in_2')
// (15, 20, 'lutff_5/in_1')
// (15, 20, 'neigh_op_tnl_5')
// (15, 21, 'neigh_op_lft_5')
// (15, 22, 'neigh_op_bnl_5')

wire n2022;
// (13, 20, 'sp4_h_r_3')
// (14, 20, 'sp4_h_r_14')
// (15, 19, 'neigh_op_tnr_3')
// (15, 20, 'neigh_op_rgt_3')
// (15, 20, 'sp4_h_r_11')
// (15, 20, 'sp4_h_r_27')
// (15, 21, 'neigh_op_bnr_3')
// (16, 18, 'sp4_r_v_b_47')
// (16, 19, 'neigh_op_top_3')
// (16, 19, 'sp4_r_v_b_34')
// (16, 20, 'lutff_3/out')
// (16, 20, 'sp4_h_r_22')
// (16, 20, 'sp4_h_r_38')
// (16, 20, 'sp4_r_v_b_23')
// (16, 21, 'local_g1_3')
// (16, 21, 'lutff_1/in_1')
// (16, 21, 'neigh_op_bot_3')
// (16, 21, 'sp4_r_v_b_10')
// (17, 17, 'sp4_v_t_47')
// (17, 18, 'sp4_v_b_47')
// (17, 19, 'neigh_op_tnl_3')
// (17, 19, 'sp4_v_b_34')
// (17, 20, 'local_g0_3')
// (17, 20, 'lutff_0/in_1')
// (17, 20, 'lutff_1/in_2')
// (17, 20, 'lutff_2/in_1')
// (17, 20, 'lutff_3/in_0')
// (17, 20, 'lutff_4/in_1')
// (17, 20, 'lutff_5/in_0')
// (17, 20, 'lutff_6/in_3')
// (17, 20, 'lutff_7/in_0')
// (17, 20, 'neigh_op_lft_3')
// (17, 20, 'sp4_h_l_38')
// (17, 20, 'sp4_h_r_3')
// (17, 20, 'sp4_h_r_35')
// (17, 20, 'sp4_v_b_23')
// (17, 21, 'local_g2_3')
// (17, 21, 'lutff_0/in_3')
// (17, 21, 'lutff_5/in_0')
// (17, 21, 'lutff_7/in_2')
// (17, 21, 'neigh_op_bnl_3')
// (17, 21, 'sp4_h_r_4')
// (17, 21, 'sp4_v_b_10')
// (18, 20, 'sp4_h_r_14')
// (18, 20, 'sp4_h_r_46')
// (18, 21, 'sp4_h_r_17')
// (19, 20, 'sp4_h_l_46')
// (19, 20, 'sp4_h_r_27')
// (19, 20, 'sp4_h_r_7')
// (19, 21, 'sp4_h_r_28')
// (20, 17, 'sp4_r_v_b_38')
// (20, 18, 'sp4_r_v_b_27')
// (20, 19, 'sp4_r_v_b_14')
// (20, 20, 'sp4_h_r_18')
// (20, 20, 'sp4_h_r_38')
// (20, 20, 'sp4_r_v_b_3')
// (20, 21, 'sp4_h_r_41')
// (21, 16, 'sp4_v_t_38')
// (21, 17, 'sp4_v_b_38')
// (21, 18, 'sp4_v_b_27')
// (21, 19, 'local_g0_6')
// (21, 19, 'lutff_3/in_1')
// (21, 19, 'sp4_v_b_14')
// (21, 20, 'sp4_h_l_38')
// (21, 20, 'sp4_h_r_31')
// (21, 20, 'sp4_v_b_3')
// (21, 21, 'local_g0_7')
// (21, 21, 'lutff_6/in_1')
// (21, 21, 'sp4_h_l_41')
// (21, 21, 'sp4_h_r_7')
// (22, 17, 'sp4_r_v_b_36')
// (22, 18, 'sp4_r_v_b_25')
// (22, 19, 'local_g2_4')
// (22, 19, 'lutff_5/in_1')
// (22, 19, 'lutff_7/in_3')
// (22, 19, 'sp4_r_v_b_12')
// (22, 20, 'sp4_h_r_42')
// (22, 20, 'sp4_r_v_b_1')
// (22, 21, 'sp4_h_r_18')
// (23, 16, 'sp4_v_t_36')
// (23, 17, 'sp4_v_b_36')
// (23, 18, 'sp4_v_b_25')
// (23, 19, 'sp4_v_b_12')
// (23, 20, 'sp4_h_l_42')
// (23, 20, 'sp4_v_b_1')
// (23, 21, 'sp4_h_r_31')
// (24, 21, 'sp4_h_r_42')
// (25, 21, 'sp4_h_l_42')

wire n2023;
// (13, 20, 'sp4_h_r_8')
// (14, 20, 'sp4_h_r_21')
// (15, 20, 'sp4_h_r_32')
// (16, 17, 'sp4_r_v_b_39')
// (16, 18, 'sp4_r_v_b_26')
// (16, 19, 'neigh_op_tnr_4')
// (16, 19, 'sp4_r_v_b_15')
// (16, 20, 'neigh_op_rgt_4')
// (16, 20, 'sp4_h_r_45')
// (16, 20, 'sp4_r_v_b_2')
// (16, 21, 'neigh_op_bnr_4')
// (17, 16, 'sp4_v_t_39')
// (17, 17, 'sp4_v_b_39')
// (17, 18, 'sp4_v_b_26')
// (17, 19, 'neigh_op_top_4')
// (17, 19, 'sp4_v_b_15')
// (17, 20, 'local_g0_2')
// (17, 20, 'lutff_4/out')
// (17, 20, 'lutff_global/cen')
// (17, 20, 'sp4_h_l_45')
// (17, 20, 'sp4_h_r_8')
// (17, 20, 'sp4_v_b_2')
// (17, 21, 'neigh_op_bot_4')
// (18, 19, 'neigh_op_tnl_4')
// (18, 20, 'neigh_op_lft_4')
// (18, 20, 'sp4_h_r_21')
// (18, 21, 'neigh_op_bnl_4')
// (19, 20, 'sp4_h_r_32')
// (20, 20, 'sp4_h_r_45')
// (21, 20, 'sp4_h_l_45')

wire n2024;
// (13, 20, 'sp4_h_r_9')
// (14, 20, 'sp4_h_r_20')
// (15, 19, 'neigh_op_tnr_6')
// (15, 20, 'neigh_op_rgt_6')
// (15, 20, 'sp4_h_r_33')
// (15, 21, 'neigh_op_bnr_6')
// (16, 17, 'sp4_r_v_b_38')
// (16, 18, 'sp4_r_v_b_27')
// (16, 19, 'neigh_op_top_6')
// (16, 19, 'sp4_r_v_b_14')
// (16, 20, 'local_g1_3')
// (16, 20, 'lutff_6/out')
// (16, 20, 'lutff_global/cen')
// (16, 20, 'sp4_h_r_44')
// (16, 20, 'sp4_r_v_b_3')
// (16, 21, 'neigh_op_bot_6')
// (17, 16, 'sp4_v_t_38')
// (17, 17, 'sp4_v_b_38')
// (17, 18, 'sp4_v_b_27')
// (17, 19, 'neigh_op_tnl_6')
// (17, 19, 'sp4_v_b_14')
// (17, 20, 'neigh_op_lft_6')
// (17, 20, 'sp4_h_l_44')
// (17, 20, 'sp4_v_b_3')
// (17, 21, 'neigh_op_bnl_6')

wire n2025;
// (13, 21, 'local_g2_5')
// (13, 21, 'lutff_4/in_3')
// (13, 21, 'neigh_op_tnr_5')
// (13, 22, 'local_g2_5')
// (13, 22, 'lutff_3/in_2')
// (13, 22, 'neigh_op_rgt_5')
// (13, 23, 'neigh_op_bnr_5')
// (14, 21, 'local_g0_5')
// (14, 21, 'lutff_3/in_2')
// (14, 21, 'lutff_7/in_2')
// (14, 21, 'neigh_op_top_5')
// (14, 22, 'lutff_5/out')
// (14, 23, 'neigh_op_bot_5')
// (15, 21, 'neigh_op_tnl_5')
// (15, 22, 'neigh_op_lft_5')
// (15, 23, 'neigh_op_bnl_5')

wire n2026;
// (13, 21, 'neigh_op_tnr_0')
// (13, 22, 'neigh_op_rgt_0')
// (13, 23, 'neigh_op_bnr_0')
// (14, 21, 'neigh_op_top_0')
// (14, 22, 'lutff_0/out')
// (14, 23, 'local_g1_0')
// (14, 23, 'lutff_3/in_2')
// (14, 23, 'neigh_op_bot_0')
// (15, 21, 'neigh_op_tnl_0')
// (15, 22, 'neigh_op_lft_0')
// (15, 23, 'neigh_op_bnl_0')

wire n2027;
// (13, 21, 'neigh_op_tnr_1')
// (13, 22, 'neigh_op_rgt_1')
// (13, 23, 'neigh_op_bnr_1')
// (14, 21, 'neigh_op_top_1')
// (14, 22, 'local_g3_1')
// (14, 22, 'lutff_1/out')
// (14, 22, 'lutff_5/in_1')
// (14, 23, 'neigh_op_bot_1')
// (15, 21, 'neigh_op_tnl_1')
// (15, 22, 'neigh_op_lft_1')
// (15, 23, 'neigh_op_bnl_1')

wire n2028;
// (13, 21, 'neigh_op_tnr_3')
// (13, 22, 'neigh_op_rgt_3')
// (13, 23, 'neigh_op_bnr_3')
// (14, 21, 'neigh_op_top_3')
// (14, 22, 'lutff_3/out')
// (14, 23, 'local_g1_3')
// (14, 23, 'lutff_2/in_2')
// (14, 23, 'neigh_op_bot_3')
// (15, 21, 'neigh_op_tnl_3')
// (15, 22, 'neigh_op_lft_3')
// (15, 23, 'neigh_op_bnl_3')

wire n2029;
// (13, 21, 'neigh_op_tnr_4')
// (13, 22, 'neigh_op_rgt_4')
// (13, 23, 'neigh_op_bnr_4')
// (14, 21, 'neigh_op_top_4')
// (14, 22, 'lutff_4/out')
// (14, 23, 'local_g1_4')
// (14, 23, 'lutff_1/in_2')
// (14, 23, 'neigh_op_bot_4')
// (15, 21, 'neigh_op_tnl_4')
// (15, 22, 'neigh_op_lft_4')
// (15, 23, 'neigh_op_bnl_4')

wire n2030;
// (13, 21, 'neigh_op_tnr_6')
// (13, 22, 'local_g3_6')
// (13, 22, 'lutff_0/in_1')
// (13, 22, 'neigh_op_rgt_6')
// (13, 23, 'local_g0_6')
// (13, 23, 'local_g1_6')
// (13, 23, 'lutff_0/in_1')
// (13, 23, 'lutff_1/in_3')
// (13, 23, 'neigh_op_bnr_6')
// (14, 21, 'neigh_op_top_6')
// (14, 22, 'lutff_6/out')
// (14, 23, 'neigh_op_bot_6')
// (15, 21, 'neigh_op_tnl_6')
// (15, 22, 'neigh_op_lft_6')
// (15, 23, 'neigh_op_bnl_6')

wire n2031;
// (13, 22, 'neigh_op_tnr_1')
// (13, 23, 'local_g2_1')
// (13, 23, 'lutff_1/in_2')
// (13, 23, 'neigh_op_rgt_1')
// (13, 24, 'neigh_op_bnr_1')
// (14, 22, 'neigh_op_top_1')
// (14, 23, 'lutff_1/out')
// (14, 24, 'neigh_op_bot_1')
// (15, 22, 'neigh_op_tnl_1')
// (15, 23, 'neigh_op_lft_1')
// (15, 24, 'neigh_op_bnl_1')

wire n2032;
// (13, 22, 'neigh_op_tnr_2')
// (13, 23, 'local_g3_2')
// (13, 23, 'lutff_2/in_1')
// (13, 23, 'neigh_op_rgt_2')
// (13, 24, 'neigh_op_bnr_2')
// (14, 22, 'neigh_op_top_2')
// (14, 23, 'lutff_2/out')
// (14, 24, 'neigh_op_bot_2')
// (15, 22, 'neigh_op_tnl_2')
// (15, 23, 'neigh_op_lft_2')
// (15, 24, 'neigh_op_bnl_2')

wire n2033;
// (13, 22, 'neigh_op_tnr_3')
// (13, 23, 'local_g3_3')
// (13, 23, 'lutff_3/in_1')
// (13, 23, 'neigh_op_rgt_3')
// (13, 24, 'neigh_op_bnr_3')
// (14, 22, 'neigh_op_top_3')
// (14, 23, 'lutff_3/out')
// (14, 24, 'neigh_op_bot_3')
// (15, 22, 'neigh_op_tnl_3')
// (15, 23, 'neigh_op_lft_3')
// (15, 24, 'neigh_op_bnl_3')

wire n2034;
// (13, 22, 'neigh_op_tnr_4')
// (13, 23, 'local_g3_4')
// (13, 23, 'lutff_4/in_1')
// (13, 23, 'neigh_op_rgt_4')
// (13, 24, 'neigh_op_bnr_4')
// (14, 22, 'neigh_op_top_4')
// (14, 23, 'lutff_4/out')
// (14, 24, 'neigh_op_bot_4')
// (15, 22, 'neigh_op_tnl_4')
// (15, 23, 'neigh_op_lft_4')
// (15, 24, 'neigh_op_bnl_4')

wire n2035;
// (13, 22, 'neigh_op_tnr_5')
// (13, 23, 'local_g3_5')
// (13, 23, 'lutff_5/in_1')
// (13, 23, 'neigh_op_rgt_5')
// (13, 24, 'neigh_op_bnr_5')
// (14, 22, 'neigh_op_top_5')
// (14, 23, 'lutff_5/out')
// (14, 24, 'neigh_op_bot_5')
// (15, 22, 'neigh_op_tnl_5')
// (15, 23, 'neigh_op_lft_5')
// (15, 24, 'neigh_op_bnl_5')

wire n2036;
// (13, 22, 'neigh_op_tnr_6')
// (13, 23, 'local_g3_6')
// (13, 23, 'lutff_6/in_1')
// (13, 23, 'neigh_op_rgt_6')
// (13, 24, 'neigh_op_bnr_6')
// (14, 22, 'neigh_op_top_6')
// (14, 23, 'lutff_6/out')
// (14, 24, 'neigh_op_bot_6')
// (15, 22, 'neigh_op_tnl_6')
// (15, 23, 'neigh_op_lft_6')
// (15, 24, 'neigh_op_bnl_6')

wire n2037;
// (13, 22, 'sp4_h_r_11')
// (14, 22, 'sp4_h_r_22')
// (15, 20, 'neigh_op_tnr_1')
// (15, 21, 'neigh_op_rgt_1')
// (15, 22, 'local_g3_3')
// (15, 22, 'lutff_global/cen')
// (15, 22, 'neigh_op_bnr_1')
// (15, 22, 'sp4_h_r_35')
// (16, 19, 'sp4_r_v_b_43')
// (16, 20, 'neigh_op_top_1')
// (16, 20, 'sp4_r_v_b_30')
// (16, 21, 'lutff_1/out')
// (16, 21, 'sp4_r_v_b_19')
// (16, 22, 'neigh_op_bot_1')
// (16, 22, 'sp4_h_r_46')
// (16, 22, 'sp4_r_v_b_6')
// (17, 18, 'sp4_v_t_43')
// (17, 19, 'sp4_v_b_43')
// (17, 20, 'neigh_op_tnl_1')
// (17, 20, 'sp4_v_b_30')
// (17, 21, 'neigh_op_lft_1')
// (17, 21, 'sp4_v_b_19')
// (17, 22, 'neigh_op_bnl_1')
// (17, 22, 'sp4_h_l_46')
// (17, 22, 'sp4_v_b_6')

wire n2038;
// (13, 22, 'sp4_r_v_b_43')
// (13, 23, 'sp4_r_v_b_30')
// (13, 24, 'sp4_r_v_b_19')
// (13, 25, 'sp4_r_v_b_6')
// (14, 21, 'sp4_h_r_11')
// (14, 21, 'sp4_h_r_6')
// (14, 21, 'sp4_v_t_43')
// (14, 22, 'sp4_v_b_43')
// (14, 23, 'sp4_v_b_30')
// (14, 24, 'sp4_v_b_19')
// (14, 25, 'sp4_v_b_6')
// (15, 20, 'neigh_op_tnr_7')
// (15, 21, 'neigh_op_rgt_7')
// (15, 21, 'sp4_h_r_19')
// (15, 21, 'sp4_h_r_22')
// (15, 22, 'neigh_op_bnr_7')
// (16, 20, 'neigh_op_top_7')
// (16, 21, 'local_g3_3')
// (16, 21, 'lutff_7/out')
// (16, 21, 'lutff_global/cen')
// (16, 21, 'sp4_h_r_30')
// (16, 21, 'sp4_h_r_35')
// (16, 22, 'neigh_op_bot_7')
// (17, 20, 'neigh_op_tnl_7')
// (17, 21, 'neigh_op_lft_7')
// (17, 21, 'sp4_h_r_43')
// (17, 21, 'sp4_h_r_46')
// (17, 22, 'neigh_op_bnl_7')
// (18, 21, 'sp4_h_l_43')
// (18, 21, 'sp4_h_l_46')

wire n2039;
// (13, 23, 'lutff_1/cout')
// (13, 23, 'lutff_2/in_3')

wire n2040;
// (13, 23, 'lutff_2/cout')
// (13, 23, 'lutff_3/in_3')

wire n2041;
// (13, 23, 'lutff_3/cout')
// (13, 23, 'lutff_4/in_3')

wire n2042;
// (13, 23, 'lutff_4/cout')
// (13, 23, 'lutff_5/in_3')

wire n2043;
// (13, 23, 'lutff_5/cout')
// (13, 23, 'lutff_6/in_3')

wire n2044;
// (14, 1, 'neigh_op_tnr_1')
// (14, 2, 'neigh_op_rgt_1')
// (14, 3, 'neigh_op_bnr_1')
// (15, 1, 'neigh_op_top_1')
// (15, 2, 'local_g3_1')
// (15, 2, 'lutff_1/out')
// (15, 2, 'lutff_5/in_1')
// (15, 3, 'neigh_op_bot_1')
// (16, 1, 'neigh_op_tnl_1')
// (16, 2, 'neigh_op_lft_1')
// (16, 3, 'neigh_op_bnl_1')

wire n2045;
// (14, 1, 'neigh_op_tnr_3')
// (14, 2, 'local_g2_3')
// (14, 2, 'lutff_4/in_3')
// (14, 2, 'neigh_op_rgt_3')
// (14, 3, 'neigh_op_bnr_3')
// (15, 1, 'neigh_op_top_3')
// (15, 2, 'lutff_3/out')
// (15, 3, 'neigh_op_bot_3')
// (16, 1, 'neigh_op_tnl_3')
// (16, 2, 'neigh_op_lft_3')
// (16, 3, 'neigh_op_bnl_3')

wire n2046;
// (14, 1, 'neigh_op_tnr_5')
// (14, 2, 'neigh_op_rgt_5')
// (14, 3, 'local_g0_5')
// (14, 3, 'lutff_5/in_0')
// (14, 3, 'neigh_op_bnr_5')
// (15, 1, 'neigh_op_top_5')
// (15, 2, 'lutff_5/out')
// (15, 3, 'neigh_op_bot_5')
// (16, 1, 'neigh_op_tnl_5')
// (16, 2, 'neigh_op_lft_5')
// (16, 3, 'neigh_op_bnl_5')

wire n2047;
// (14, 1, 'neigh_op_tnr_6')
// (14, 2, 'neigh_op_rgt_6')
// (14, 3, 'neigh_op_bnr_6')
// (15, 1, 'neigh_op_top_6')
// (15, 2, 'local_g1_6')
// (15, 2, 'lutff_5/in_0')
// (15, 2, 'lutff_6/out')
// (15, 3, 'neigh_op_bot_6')
// (16, 1, 'neigh_op_tnl_6')
// (16, 2, 'neigh_op_lft_6')
// (16, 3, 'neigh_op_bnl_6')

wire n2048;
// (14, 1, 'neigh_op_tnr_7')
// (14, 2, 'neigh_op_rgt_7')
// (14, 3, 'neigh_op_bnr_7')
// (15, 1, 'neigh_op_top_7')
// (15, 1, 'sp4_r_v_b_42')
// (15, 2, 'lutff_7/out')
// (15, 2, 'sp4_r_v_b_31')
// (15, 3, 'neigh_op_bot_7')
// (15, 3, 'sp4_r_v_b_18')
// (15, 4, 'local_g1_7')
// (15, 4, 'lutff_4/in_0')
// (15, 4, 'sp4_r_v_b_7')
// (16, 0, 'span4_vert_42')
// (16, 1, 'neigh_op_tnl_7')
// (16, 1, 'sp4_v_b_42')
// (16, 2, 'neigh_op_lft_7')
// (16, 2, 'sp4_v_b_31')
// (16, 3, 'neigh_op_bnl_7')
// (16, 3, 'sp4_v_b_18')
// (16, 4, 'sp4_v_b_7')

reg n2049 = 0;
// (14, 2, 'neigh_op_tnr_0')
// (14, 2, 'sp4_r_v_b_45')
// (14, 3, 'local_g3_0')
// (14, 3, 'lutff_0/in_3')
// (14, 3, 'neigh_op_rgt_0')
// (14, 3, 'sp4_r_v_b_32')
// (14, 4, 'neigh_op_bnr_0')
// (14, 4, 'sp4_r_v_b_21')
// (14, 4, 'sp4_r_v_b_37')
// (14, 5, 'sp4_r_v_b_24')
// (14, 5, 'sp4_r_v_b_8')
// (14, 6, 'sp4_r_v_b_13')
// (14, 6, 'sp4_r_v_b_46')
// (14, 7, 'sp4_r_v_b_0')
// (14, 7, 'sp4_r_v_b_35')
// (14, 8, 'local_g3_6')
// (14, 8, 'lutff_2/in_1')
// (14, 8, 'sp4_r_v_b_22')
// (14, 8, 'sp4_r_v_b_37')
// (14, 9, 'sp4_r_v_b_11')
// (14, 9, 'sp4_r_v_b_24')
// (14, 10, 'local_g2_5')
// (14, 10, 'lutff_5/in_2')
// (14, 10, 'sp4_r_v_b_13')
// (14, 11, 'sp4_r_v_b_0')
// (15, 0, 'span12_vert_20')
// (15, 1, 'sp12_v_b_20')
// (15, 1, 'sp4_v_t_45')
// (15, 2, 'neigh_op_top_0')
// (15, 2, 'sp12_v_b_19')
// (15, 2, 'sp4_v_b_45')
// (15, 3, 'lutff_0/out')
// (15, 3, 'sp12_v_b_16')
// (15, 3, 'sp4_h_r_0')
// (15, 3, 'sp4_v_b_32')
// (15, 3, 'sp4_v_t_37')
// (15, 4, 'neigh_op_bot_0')
// (15, 4, 'sp12_v_b_15')
// (15, 4, 'sp4_v_b_21')
// (15, 4, 'sp4_v_b_37')
// (15, 5, 'sp12_v_b_12')
// (15, 5, 'sp4_v_b_24')
// (15, 5, 'sp4_v_b_8')
// (15, 5, 'sp4_v_t_46')
// (15, 6, 'local_g3_6')
// (15, 6, 'lutff_2/in_3')
// (15, 6, 'sp12_v_b_11')
// (15, 6, 'sp4_v_b_13')
// (15, 6, 'sp4_v_b_46')
// (15, 7, 'sp12_v_b_8')
// (15, 7, 'sp4_v_b_0')
// (15, 7, 'sp4_v_b_35')
// (15, 7, 'sp4_v_t_37')
// (15, 8, 'sp12_v_b_7')
// (15, 8, 'sp4_v_b_22')
// (15, 8, 'sp4_v_b_37')
// (15, 9, 'sp12_v_b_4')
// (15, 9, 'sp4_v_b_11')
// (15, 9, 'sp4_v_b_24')
// (15, 10, 'local_g2_3')
// (15, 10, 'lutff_1/in_0')
// (15, 10, 'sp12_v_b_3')
// (15, 10, 'sp4_v_b_13')
// (15, 11, 'sp12_v_b_0')
// (15, 11, 'sp4_v_b_0')
// (16, 2, 'neigh_op_tnl_0')
// (16, 3, 'neigh_op_lft_0')
// (16, 3, 'sp4_h_r_13')
// (16, 4, 'neigh_op_bnl_0')
// (17, 3, 'sp4_h_r_24')
// (18, 3, 'sp4_h_r_37')
// (19, 3, 'sp4_h_l_37')

wire n2050;
// (14, 3, 'neigh_op_tnr_4')
// (14, 4, 'neigh_op_rgt_4')
// (14, 5, 'neigh_op_bnr_4')
// (15, 3, 'neigh_op_top_4')
// (15, 4, 'local_g0_4')
// (15, 4, 'lutff_4/out')
// (15, 4, 'lutff_7/in_1')
// (15, 5, 'neigh_op_bot_4')
// (16, 3, 'neigh_op_tnl_4')
// (16, 4, 'neigh_op_lft_4')
// (16, 5, 'neigh_op_bnl_4')

wire n2051;
// (14, 3, 'neigh_op_tnr_5')
// (14, 4, 'neigh_op_rgt_5')
// (14, 5, 'neigh_op_bnr_5')
// (15, 3, 'neigh_op_top_5')
// (15, 4, 'local_g0_5')
// (15, 4, 'lutff_4/in_1')
// (15, 4, 'lutff_5/out')
// (15, 5, 'neigh_op_bot_5')
// (16, 3, 'neigh_op_tnl_5')
// (16, 4, 'neigh_op_lft_5')
// (16, 5, 'neigh_op_bnl_5')

wire n2052;
// (14, 3, 'neigh_op_tnr_7')
// (14, 4, 'neigh_op_rgt_7')
// (14, 5, 'neigh_op_bnr_7')
// (15, 3, 'neigh_op_top_7')
// (15, 4, 'local_g0_7')
// (15, 4, 'lutff_6/in_1')
// (15, 4, 'lutff_7/out')
// (15, 5, 'neigh_op_bot_7')
// (16, 3, 'neigh_op_tnl_7')
// (16, 4, 'neigh_op_lft_7')
// (16, 5, 'neigh_op_bnl_7')

reg n2053 = 0;
// (14, 3, 'sp4_r_v_b_40')
// (14, 4, 'sp4_r_v_b_29')
// (14, 5, 'sp4_r_v_b_16')
// (14, 6, 'sp4_r_v_b_5')
// (14, 7, 'sp4_r_v_b_45')
// (14, 8, 'local_g0_3')
// (14, 8, 'lutff_1/in_0')
// (14, 8, 'sp4_r_v_b_32')
// (14, 9, 'sp4_r_v_b_21')
// (14, 10, 'sp4_r_v_b_8')
// (15, 1, 'neigh_op_tnr_3')
// (15, 2, 'local_g3_3')
// (15, 2, 'lutff_3/in_3')
// (15, 2, 'neigh_op_rgt_3')
// (15, 2, 'sp4_h_r_11')
// (15, 2, 'sp4_r_v_b_38')
// (15, 2, 'sp4_v_t_40')
// (15, 3, 'neigh_op_bnr_3')
// (15, 3, 'sp4_r_v_b_27')
// (15, 3, 'sp4_v_b_40')
// (15, 4, 'sp4_r_v_b_14')
// (15, 4, 'sp4_v_b_29')
// (15, 5, 'sp4_r_v_b_3')
// (15, 5, 'sp4_v_b_16')
// (15, 6, 'sp4_r_v_b_43')
// (15, 6, 'sp4_v_b_5')
// (15, 6, 'sp4_v_t_45')
// (15, 7, 'sp4_r_v_b_30')
// (15, 7, 'sp4_v_b_45')
// (15, 8, 'sp4_r_v_b_19')
// (15, 8, 'sp4_v_b_32')
// (15, 9, 'sp4_r_v_b_6')
// (15, 9, 'sp4_v_b_21')
// (15, 10, 'sp4_v_b_8')
// (16, 1, 'neigh_op_top_3')
// (16, 1, 'sp4_v_t_38')
// (16, 2, 'lutff_3/out')
// (16, 2, 'sp4_h_r_22')
// (16, 2, 'sp4_v_b_38')
// (16, 3, 'neigh_op_bot_3')
// (16, 3, 'sp4_v_b_27')
// (16, 4, 'sp4_v_b_14')
// (16, 5, 'sp4_v_b_3')
// (16, 5, 'sp4_v_t_43')
// (16, 6, 'sp4_v_b_43')
// (16, 7, 'sp4_v_b_30')
// (16, 8, 'local_g0_3')
// (16, 8, 'lutff_0/in_3')
// (16, 8, 'lutff_4/in_3')
// (16, 8, 'sp4_v_b_19')
// (16, 9, 'sp4_v_b_6')
// (17, 1, 'neigh_op_tnl_3')
// (17, 2, 'neigh_op_lft_3')
// (17, 2, 'sp4_h_r_35')
// (17, 3, 'neigh_op_bnl_3')
// (18, 2, 'sp4_h_r_46')
// (19, 2, 'sp4_h_l_46')

wire n2054;
// (14, 4, 'neigh_op_tnr_2')
// (14, 5, 'neigh_op_rgt_2')
// (14, 6, 'neigh_op_bnr_2')
// (15, 4, 'neigh_op_top_2')
// (15, 5, 'lutff_2/out')
// (15, 6, 'local_g1_2')
// (15, 6, 'lutff_1/in_0')
// (15, 6, 'neigh_op_bot_2')
// (16, 4, 'neigh_op_tnl_2')
// (16, 5, 'neigh_op_lft_2')
// (16, 6, 'neigh_op_bnl_2')

wire n2055;
// (14, 5, 'neigh_op_tnr_1')
// (14, 6, 'neigh_op_rgt_1')
// (14, 7, 'neigh_op_bnr_1')
// (15, 5, 'neigh_op_top_1')
// (15, 6, 'lutff_1/out')
// (15, 7, 'local_g1_1')
// (15, 7, 'lutff_0/in_0')
// (15, 7, 'neigh_op_bot_1')
// (16, 5, 'neigh_op_tnl_1')
// (16, 6, 'neigh_op_lft_1')
// (16, 7, 'neigh_op_bnl_1')

wire n2056;
// (14, 5, 'neigh_op_tnr_2')
// (14, 6, 'neigh_op_rgt_2')
// (14, 7, 'neigh_op_bnr_2')
// (15, 5, 'neigh_op_top_2')
// (15, 6, 'lutff_2/out')
// (15, 7, 'local_g0_2')
// (15, 7, 'lutff_7/in_3')
// (15, 7, 'neigh_op_bot_2')
// (16, 5, 'neigh_op_tnl_2')
// (16, 6, 'neigh_op_lft_2')
// (16, 7, 'neigh_op_bnl_2')

wire n2057;
// (14, 5, 'neigh_op_tnr_6')
// (14, 6, 'neigh_op_rgt_6')
// (14, 7, 'neigh_op_bnr_6')
// (15, 5, 'neigh_op_top_6')
// (15, 6, 'lutff_6/out')
// (15, 7, 'local_g1_6')
// (15, 7, 'lutff_7/in_2')
// (15, 7, 'neigh_op_bot_6')
// (16, 5, 'neigh_op_tnl_6')
// (16, 6, 'neigh_op_lft_6')
// (16, 7, 'neigh_op_bnl_6')

wire n2058;
// (14, 5, 'neigh_op_tnr_7')
// (14, 6, 'neigh_op_rgt_7')
// (14, 7, 'neigh_op_bnr_7')
// (15, 5, 'neigh_op_top_7')
// (15, 6, 'lutff_7/out')
// (15, 7, 'local_g1_7')
// (15, 7, 'lutff_2/in_0')
// (15, 7, 'neigh_op_bot_7')
// (16, 5, 'neigh_op_tnl_7')
// (16, 6, 'neigh_op_lft_7')
// (16, 7, 'neigh_op_bnl_7')

wire n2059;
// (14, 6, 'neigh_op_tnr_1')
// (14, 7, 'neigh_op_rgt_1')
// (14, 8, 'neigh_op_bnr_1')
// (15, 6, 'neigh_op_top_1')
// (15, 7, 'local_g2_1')
// (15, 7, 'lutff_1/out')
// (15, 7, 'lutff_7/in_0')
// (15, 8, 'neigh_op_bot_1')
// (16, 6, 'neigh_op_tnl_1')
// (16, 7, 'neigh_op_lft_1')
// (16, 8, 'neigh_op_bnl_1')

wire n2060;
// (14, 6, 'neigh_op_tnr_2')
// (14, 7, 'neigh_op_rgt_2')
// (14, 7, 'sp4_r_v_b_36')
// (14, 8, 'neigh_op_bnr_2')
// (14, 8, 'sp4_r_v_b_25')
// (14, 9, 'sp4_r_v_b_12')
// (14, 10, 'sp4_r_v_b_1')
// (15, 6, 'neigh_op_top_2')
// (15, 6, 'sp4_v_t_36')
// (15, 7, 'lutff_2/out')
// (15, 7, 'sp4_v_b_36')
// (15, 8, 'neigh_op_bot_2')
// (15, 8, 'sp4_v_b_25')
// (15, 9, 'sp4_v_b_12')
// (15, 10, 'local_g0_1')
// (15, 10, 'lutff_5/in_0')
// (15, 10, 'sp4_v_b_1')
// (16, 6, 'neigh_op_tnl_2')
// (16, 7, 'neigh_op_lft_2')
// (16, 8, 'neigh_op_bnl_2')

wire n2061;
// (14, 6, 'neigh_op_tnr_3')
// (14, 7, 'neigh_op_rgt_3')
// (14, 8, 'neigh_op_bnr_3')
// (15, 6, 'neigh_op_top_3')
// (15, 7, 'local_g3_3')
// (15, 7, 'lutff_3/out')
// (15, 7, 'lutff_7/in_1')
// (15, 8, 'neigh_op_bot_3')
// (16, 6, 'neigh_op_tnl_3')
// (16, 7, 'neigh_op_lft_3')
// (16, 8, 'neigh_op_bnl_3')

wire n2062;
// (14, 6, 'neigh_op_tnr_4')
// (14, 7, 'neigh_op_rgt_4')
// (14, 7, 'sp4_r_v_b_40')
// (14, 8, 'neigh_op_bnr_4')
// (14, 8, 'sp4_r_v_b_29')
// (14, 9, 'sp4_r_v_b_16')
// (14, 10, 'sp4_r_v_b_5')
// (15, 6, 'neigh_op_top_4')
// (15, 6, 'sp4_v_t_40')
// (15, 7, 'lutff_4/out')
// (15, 7, 'sp4_v_b_40')
// (15, 8, 'neigh_op_bot_4')
// (15, 8, 'sp4_v_b_29')
// (15, 9, 'sp4_v_b_16')
// (15, 10, 'local_g0_5')
// (15, 10, 'lutff_7/in_0')
// (15, 10, 'sp4_v_b_5')
// (16, 6, 'neigh_op_tnl_4')
// (16, 7, 'neigh_op_lft_4')
// (16, 8, 'neigh_op_bnl_4')

wire n2063;
// (14, 6, 'neigh_op_tnr_6')
// (14, 7, 'neigh_op_rgt_6')
// (14, 8, 'neigh_op_bnr_6')
// (15, 6, 'neigh_op_top_6')
// (15, 7, 'local_g2_6')
// (15, 7, 'lutff_0/in_2')
// (15, 7, 'lutff_6/out')
// (15, 8, 'neigh_op_bot_6')
// (16, 6, 'neigh_op_tnl_6')
// (16, 7, 'neigh_op_lft_6')
// (16, 8, 'neigh_op_bnl_6')

wire n2064;
// (14, 6, 'neigh_op_tnr_7')
// (14, 7, 'neigh_op_rgt_7')
// (14, 8, 'neigh_op_bnr_7')
// (15, 6, 'neigh_op_top_7')
// (15, 7, 'local_g2_7')
// (15, 7, 'lutff_0/in_3')
// (15, 7, 'lutff_7/out')
// (15, 8, 'neigh_op_bot_7')
// (16, 6, 'neigh_op_tnl_7')
// (16, 7, 'neigh_op_lft_7')
// (16, 8, 'neigh_op_bnl_7')

wire n2065;
// (14, 6, 'sp4_h_r_3')
// (15, 6, 'local_g1_6')
// (15, 6, 'lutff_4/in_3')
// (15, 6, 'sp4_h_r_14')
// (16, 5, 'neigh_op_tnr_3')
// (16, 6, 'neigh_op_rgt_3')
// (16, 6, 'sp4_h_r_27')
// (16, 7, 'neigh_op_bnr_3')
// (17, 5, 'neigh_op_top_3')
// (17, 6, 'lutff_3/out')
// (17, 6, 'sp4_h_r_38')
// (17, 7, 'neigh_op_bot_3')
// (18, 5, 'neigh_op_tnl_3')
// (18, 6, 'neigh_op_lft_3')
// (18, 6, 'sp4_h_l_38')
// (18, 7, 'neigh_op_bnl_3')

wire n2066;
// (14, 6, 'sp4_h_r_5')
// (15, 5, 'sp4_r_v_b_44')
// (15, 6, 'local_g0_0')
// (15, 6, 'local_g2_1')
// (15, 6, 'lutff_0/in_0')
// (15, 6, 'lutff_3/in_2')
// (15, 6, 'lutff_4/in_2')
// (15, 6, 'lutff_5/in_1')
// (15, 6, 'sp4_h_r_16')
// (15, 6, 'sp4_r_v_b_33')
// (15, 7, 'sp4_r_v_b_20')
// (15, 8, 'sp4_r_v_b_9')
// (16, 4, 'sp4_v_t_44')
// (16, 5, 'sp4_r_v_b_45')
// (16, 5, 'sp4_v_b_44')
// (16, 6, 'sp4_h_r_29')
// (16, 6, 'sp4_r_v_b_32')
// (16, 6, 'sp4_v_b_33')
// (16, 7, 'sp4_r_v_b_21')
// (16, 7, 'sp4_v_b_20')
// (16, 8, 'sp4_h_r_4')
// (16, 8, 'sp4_r_v_b_8')
// (16, 8, 'sp4_v_b_9')
// (16, 12, 'sp4_h_r_8')
// (17, 1, 'sp4_r_v_b_46')
// (17, 2, 'sp4_r_v_b_35')
// (17, 3, 'sp4_r_v_b_22')
// (17, 4, 'sp4_r_v_b_11')
// (17, 4, 'sp4_v_t_45')
// (17, 5, 'sp4_v_b_45')
// (17, 6, 'sp4_h_r_40')
// (17, 6, 'sp4_v_b_32')
// (17, 7, 'local_g0_5')
// (17, 7, 'lutff_5/in_2')
// (17, 7, 'sp4_v_b_21')
// (17, 8, 'sp4_h_r_17')
// (17, 8, 'sp4_h_r_8')
// (17, 8, 'sp4_v_b_8')
// (17, 12, 'local_g0_5')
// (17, 12, 'lutff_1/in_2')
// (17, 12, 'sp4_h_r_21')
// (18, 0, 'span4_vert_46')
// (18, 1, 'sp4_v_b_46')
// (18, 2, 'sp4_v_b_35')
// (18, 3, 'local_g0_6')
// (18, 3, 'lutff_1/in_3')
// (18, 3, 'lutff_2/in_0')
// (18, 3, 'lutff_7/in_3')
// (18, 3, 'sp4_v_b_22')
// (18, 4, 'sp4_h_r_6')
// (18, 4, 'sp4_v_b_11')
// (18, 6, 'sp4_h_l_40')
// (18, 6, 'sp4_h_r_2')
// (18, 8, 'sp4_h_r_21')
// (18, 8, 'sp4_h_r_28')
// (18, 12, 'sp4_h_r_32')
// (19, 4, 'sp4_h_r_19')
// (19, 6, 'sp4_h_r_15')
// (19, 8, 'sp4_h_r_32')
// (19, 8, 'sp4_h_r_41')
// (19, 9, 'sp4_r_v_b_45')
// (19, 10, 'sp4_r_v_b_32')
// (19, 11, 'sp4_r_v_b_21')
// (19, 12, 'sp4_h_r_45')
// (19, 12, 'sp4_r_v_b_8')
// (20, 4, 'sp4_h_r_30')
// (20, 6, 'sp4_h_r_26')
// (20, 8, 'sp4_h_l_41')
// (20, 8, 'sp4_h_r_45')
// (20, 8, 'sp4_h_r_8')
// (20, 8, 'sp4_v_t_45')
// (20, 9, 'sp4_v_b_45')
// (20, 10, 'sp4_v_b_32')
// (20, 11, 'sp4_v_b_21')
// (20, 12, 'sp4_h_l_45')
// (20, 12, 'sp4_v_b_8')
// (21, 4, 'sp4_h_r_43')
// (21, 5, 'sp4_r_v_b_37')
// (21, 6, 'sp4_h_r_39')
// (21, 6, 'sp4_r_v_b_24')
// (21, 7, 'neigh_op_tnr_0')
// (21, 7, 'sp4_r_v_b_13')
// (21, 7, 'sp4_r_v_b_45')
// (21, 8, 'neigh_op_rgt_0')
// (21, 8, 'sp4_h_l_45')
// (21, 8, 'sp4_h_r_21')
// (21, 8, 'sp4_h_r_5')
// (21, 8, 'sp4_r_v_b_0')
// (21, 8, 'sp4_r_v_b_32')
// (21, 9, 'neigh_op_bnr_0')
// (21, 9, 'sp4_r_v_b_21')
// (21, 10, 'sp4_r_v_b_8')
// (22, 4, 'sp4_h_l_43')
// (22, 4, 'sp4_v_t_37')
// (22, 5, 'sp4_v_b_37')
// (22, 6, 'sp4_h_l_39')
// (22, 6, 'sp4_v_b_24')
// (22, 6, 'sp4_v_t_45')
// (22, 7, 'neigh_op_top_0')
// (22, 7, 'sp4_v_b_13')
// (22, 7, 'sp4_v_b_45')
// (22, 8, 'lutff_0/out')
// (22, 8, 'sp4_h_r_16')
// (22, 8, 'sp4_h_r_32')
// (22, 8, 'sp4_v_b_0')
// (22, 8, 'sp4_v_b_32')
// (22, 9, 'neigh_op_bot_0')
// (22, 9, 'sp4_v_b_21')
// (22, 10, 'local_g0_0')
// (22, 10, 'lutff_3/in_1')
// (22, 10, 'lutff_4/in_0')
// (22, 10, 'sp4_v_b_8')
// (23, 7, 'neigh_op_tnl_0')
// (23, 8, 'neigh_op_lft_0')
// (23, 8, 'sp4_h_r_29')
// (23, 8, 'sp4_h_r_45')
// (23, 9, 'neigh_op_bnl_0')
// (24, 8, 'sp4_h_l_45')
// (24, 8, 'sp4_h_r_40')
// (25, 8, 'sp4_h_l_40')

reg n2067 = 0;
// (14, 6, 'sp4_r_v_b_43')
// (14, 6, 'sp4_r_v_b_44')
// (14, 7, 'sp4_r_v_b_30')
// (14, 7, 'sp4_r_v_b_33')
// (14, 8, 'local_g3_3')
// (14, 8, 'lutff_5/in_1')
// (14, 8, 'sp4_r_v_b_19')
// (14, 8, 'sp4_r_v_b_20')
// (14, 9, 'local_g2_1')
// (14, 9, 'lutff_4/in_3')
// (14, 9, 'sp4_r_v_b_6')
// (14, 9, 'sp4_r_v_b_9')
// (14, 10, 'sp4_r_v_b_43')
// (14, 11, 'sp4_r_v_b_30')
// (14, 12, 'sp4_r_v_b_19')
// (14, 13, 'sp4_r_v_b_6')
// (15, 5, 'sp4_v_t_43')
// (15, 5, 'sp4_v_t_44')
// (15, 6, 'sp4_v_b_43')
// (15, 6, 'sp4_v_b_44')
// (15, 7, 'sp4_r_v_b_44')
// (15, 7, 'sp4_v_b_30')
// (15, 7, 'sp4_v_b_33')
// (15, 8, 'sp4_r_v_b_33')
// (15, 8, 'sp4_v_b_19')
// (15, 8, 'sp4_v_b_20')
// (15, 9, 'local_g3_4')
// (15, 9, 'lutff_3/in_0')
// (15, 9, 'sp4_r_v_b_20')
// (15, 9, 'sp4_v_b_6')
// (15, 9, 'sp4_v_b_9')
// (15, 9, 'sp4_v_t_43')
// (15, 10, 'sp4_r_v_b_9')
// (15, 10, 'sp4_v_b_43')
// (15, 11, 'sp4_r_v_b_36')
// (15, 11, 'sp4_v_b_30')
// (15, 12, 'neigh_op_tnr_6')
// (15, 12, 'sp4_r_v_b_25')
// (15, 12, 'sp4_v_b_19')
// (15, 13, 'neigh_op_rgt_6')
// (15, 13, 'sp4_h_r_1')
// (15, 13, 'sp4_r_v_b_12')
// (15, 13, 'sp4_v_b_6')
// (15, 14, 'neigh_op_bnr_6')
// (15, 14, 'sp4_r_v_b_1')
// (16, 6, 'sp4_v_t_44')
// (16, 7, 'sp4_r_v_b_37')
// (16, 7, 'sp4_v_b_44')
// (16, 8, 'sp4_r_v_b_24')
// (16, 8, 'sp4_r_v_b_45')
// (16, 8, 'sp4_v_b_33')
// (16, 9, 'sp4_r_v_b_13')
// (16, 9, 'sp4_r_v_b_32')
// (16, 9, 'sp4_v_b_20')
// (16, 10, 'local_g1_1')
// (16, 10, 'lutff_5/in_3')
// (16, 10, 'sp4_h_r_1')
// (16, 10, 'sp4_r_v_b_0')
// (16, 10, 'sp4_r_v_b_21')
// (16, 10, 'sp4_v_b_9')
// (16, 10, 'sp4_v_t_36')
// (16, 11, 'sp4_r_v_b_37')
// (16, 11, 'sp4_r_v_b_8')
// (16, 11, 'sp4_v_b_36')
// (16, 12, 'neigh_op_top_6')
// (16, 12, 'sp4_r_v_b_24')
// (16, 12, 'sp4_r_v_b_40')
// (16, 12, 'sp4_v_b_25')
// (16, 13, 'local_g2_6')
// (16, 13, 'lutff_2/in_2')
// (16, 13, 'lutff_6/out')
// (16, 13, 'sp4_h_r_12')
// (16, 13, 'sp4_r_v_b_13')
// (16, 13, 'sp4_r_v_b_29')
// (16, 13, 'sp4_v_b_12')
// (16, 14, 'neigh_op_bot_6')
// (16, 14, 'sp4_r_v_b_0')
// (16, 14, 'sp4_r_v_b_16')
// (16, 14, 'sp4_v_b_1')
// (16, 15, 'sp4_r_v_b_5')
// (17, 6, 'sp4_v_t_37')
// (17, 7, 'sp4_v_b_37')
// (17, 7, 'sp4_v_t_45')
// (17, 8, 'local_g2_0')
// (17, 8, 'lutff_5/in_3')
// (17, 8, 'sp4_v_b_24')
// (17, 8, 'sp4_v_b_45')
// (17, 9, 'local_g3_0')
// (17, 9, 'lutff_0/in_3')
// (17, 9, 'sp4_v_b_13')
// (17, 9, 'sp4_v_b_32')
// (17, 10, 'sp4_h_r_12')
// (17, 10, 'sp4_v_b_0')
// (17, 10, 'sp4_v_b_21')
// (17, 10, 'sp4_v_t_37')
// (17, 11, 'sp4_v_b_37')
// (17, 11, 'sp4_v_b_8')
// (17, 11, 'sp4_v_t_40')
// (17, 12, 'neigh_op_tnl_6')
// (17, 12, 'sp4_v_b_24')
// (17, 12, 'sp4_v_b_40')
// (17, 13, 'neigh_op_lft_6')
// (17, 13, 'sp4_h_r_25')
// (17, 13, 'sp4_v_b_13')
// (17, 13, 'sp4_v_b_29')
// (17, 14, 'neigh_op_bnl_6')
// (17, 14, 'sp4_v_b_0')
// (17, 14, 'sp4_v_b_16')
// (17, 15, 'sp4_v_b_5')
// (18, 10, 'local_g3_1')
// (18, 10, 'lutff_4/in_2')
// (18, 10, 'sp4_h_r_25')
// (18, 10, 'sp4_r_v_b_36')
// (18, 11, 'sp4_r_v_b_25')
// (18, 12, 'sp4_r_v_b_12')
// (18, 13, 'sp4_h_r_36')
// (18, 13, 'sp4_r_v_b_1')
// (19, 9, 'sp4_h_r_1')
// (19, 9, 'sp4_v_t_36')
// (19, 10, 'sp4_h_r_36')
// (19, 10, 'sp4_v_b_36')
// (19, 11, 'sp4_v_b_25')
// (19, 12, 'sp4_v_b_12')
// (19, 13, 'sp4_h_l_36')
// (19, 13, 'sp4_v_b_1')
// (20, 9, 'local_g0_4')
// (20, 9, 'lutff_7/in_1')
// (20, 9, 'sp4_h_r_12')
// (20, 10, 'sp4_h_l_36')
// (21, 9, 'sp4_h_r_25')
// (22, 9, 'sp4_h_r_36')
// (23, 9, 'sp4_h_l_36')

wire n2068;
// (14, 7, 'neigh_op_tnr_0')
// (14, 8, 'neigh_op_rgt_0')
// (14, 9, 'neigh_op_bnr_0')
// (15, 7, 'neigh_op_top_0')
// (15, 8, 'local_g1_0')
// (15, 8, 'lutff_0/out')
// (15, 8, 'lutff_7/in_2')
// (15, 9, 'neigh_op_bot_0')
// (16, 7, 'neigh_op_tnl_0')
// (16, 8, 'neigh_op_lft_0')
// (16, 9, 'neigh_op_bnl_0')

reg n2069 = 0;
// (14, 7, 'neigh_op_tnr_1')
// (14, 8, 'neigh_op_rgt_1')
// (14, 8, 'sp4_h_r_7')
// (14, 9, 'neigh_op_bnr_1')
// (15, 7, 'neigh_op_top_1')
// (15, 8, 'lutff_1/out')
// (15, 8, 'sp4_h_r_18')
// (15, 9, 'neigh_op_bot_1')
// (16, 7, 'local_g3_1')
// (16, 7, 'lutff_0/in_0')
// (16, 7, 'neigh_op_tnl_1')
// (16, 8, 'neigh_op_lft_1')
// (16, 8, 'sp4_h_r_31')
// (16, 9, 'neigh_op_bnl_1')
// (17, 8, 'sp4_h_r_42')
// (17, 9, 'sp4_r_v_b_42')
// (17, 10, 'sp4_r_v_b_31')
// (17, 11, 'sp4_r_v_b_18')
// (17, 12, 'sp4_r_v_b_7')
// (18, 8, 'sp4_h_l_42')
// (18, 8, 'sp4_v_t_42')
// (18, 9, 'local_g2_2')
// (18, 9, 'lutff_6/in_0')
// (18, 9, 'sp4_v_b_42')
// (18, 10, 'sp4_v_b_31')
// (18, 11, 'sp4_v_b_18')
// (18, 12, 'sp4_v_b_7')

wire n2070;
// (14, 7, 'neigh_op_tnr_2')
// (14, 8, 'local_g3_2')
// (14, 8, 'lutff_3/in_2')
// (14, 8, 'neigh_op_rgt_2')
// (14, 9, 'neigh_op_bnr_2')
// (15, 7, 'neigh_op_top_2')
// (15, 8, 'lutff_2/out')
// (15, 9, 'neigh_op_bot_2')
// (16, 7, 'neigh_op_tnl_2')
// (16, 8, 'neigh_op_lft_2')
// (16, 9, 'neigh_op_bnl_2')

wire n2071;
// (14, 7, 'neigh_op_tnr_3')
// (14, 8, 'neigh_op_rgt_3')
// (14, 9, 'neigh_op_bnr_3')
// (15, 7, 'neigh_op_top_3')
// (15, 8, 'lutff_3/out')
// (15, 9, 'local_g0_3')
// (15, 9, 'lutff_4/in_1')
// (15, 9, 'neigh_op_bot_3')
// (16, 7, 'neigh_op_tnl_3')
// (16, 8, 'neigh_op_lft_3')
// (16, 9, 'neigh_op_bnl_3')

reg n2072 = 0;
// (14, 7, 'neigh_op_tnr_4')
// (14, 8, 'neigh_op_rgt_4')
// (14, 9, 'neigh_op_bnr_4')
// (15, 7, 'neigh_op_top_4')
// (15, 8, 'lutff_4/out')
// (15, 8, 'sp4_h_r_8')
// (15, 9, 'neigh_op_bot_4')
// (16, 7, 'local_g3_4')
// (16, 7, 'lutff_5/in_0')
// (16, 7, 'neigh_op_tnl_4')
// (16, 8, 'neigh_op_lft_4')
// (16, 8, 'sp4_h_r_21')
// (16, 9, 'neigh_op_bnl_4')
// (17, 8, 'local_g3_0')
// (17, 8, 'lutff_2/in_3')
// (17, 8, 'sp4_h_r_32')
// (18, 8, 'sp4_h_r_45')
// (19, 8, 'sp4_h_l_45')

wire n2073;
// (14, 7, 'neigh_op_tnr_5')
// (14, 8, 'neigh_op_rgt_5')
// (14, 9, 'neigh_op_bnr_5')
// (15, 7, 'neigh_op_top_5')
// (15, 8, 'lutff_5/out')
// (15, 9, 'local_g1_5')
// (15, 9, 'lutff_7/in_1')
// (15, 9, 'neigh_op_bot_5')
// (16, 7, 'neigh_op_tnl_5')
// (16, 8, 'neigh_op_lft_5')
// (16, 9, 'neigh_op_bnl_5')

wire n2074;
// (14, 7, 'neigh_op_tnr_6')
// (14, 8, 'neigh_op_rgt_6')
// (14, 9, 'neigh_op_bnr_6')
// (15, 7, 'neigh_op_top_6')
// (15, 8, 'local_g1_6')
// (15, 8, 'lutff_3/in_2')
// (15, 8, 'lutff_6/out')
// (15, 9, 'neigh_op_bot_6')
// (16, 7, 'neigh_op_tnl_6')
// (16, 8, 'neigh_op_lft_6')
// (16, 9, 'neigh_op_bnl_6')

wire n2075;
// (14, 7, 'neigh_op_tnr_7')
// (14, 8, 'neigh_op_rgt_7')
// (14, 9, 'neigh_op_bnr_7')
// (15, 7, 'neigh_op_top_7')
// (15, 8, 'lutff_7/out')
// (15, 9, 'local_g1_7')
// (15, 9, 'lutff_6/in_2')
// (15, 9, 'neigh_op_bot_7')
// (16, 7, 'neigh_op_tnl_7')
// (16, 8, 'neigh_op_lft_7')
// (16, 9, 'neigh_op_bnl_7')

wire n2076;
// (14, 8, 'local_g1_3')
// (14, 8, 'lutff_global/cen')
// (14, 8, 'sp4_h_r_11')
// (15, 8, 'sp4_h_r_22')
// (15, 9, 'sp4_r_v_b_43')
// (15, 10, 'sp4_r_v_b_30')
// (15, 11, 'sp4_r_v_b_19')
// (15, 12, 'sp4_r_v_b_6')
// (16, 8, 'sp4_h_r_0')
// (16, 8, 'sp4_h_r_35')
// (16, 8, 'sp4_v_t_43')
// (16, 9, 'sp4_v_b_43')
// (16, 10, 'sp4_v_b_30')
// (16, 11, 'local_g1_3')
// (16, 11, 'lutff_global/cen')
// (16, 11, 'sp4_v_b_19')
// (16, 12, 'sp4_v_b_6')
// (17, 7, 'neigh_op_tnr_4')
// (17, 8, 'neigh_op_rgt_4')
// (17, 8, 'sp4_h_r_13')
// (17, 8, 'sp4_h_r_46')
// (17, 9, 'neigh_op_bnr_4')
// (18, 0, 'span12_vert_23')
// (18, 1, 'sp12_v_b_23')
// (18, 2, 'sp12_v_b_20')
// (18, 3, 'sp12_v_b_19')
// (18, 4, 'sp12_v_b_16')
// (18, 5, 'sp12_v_b_15')
// (18, 6, 'sp12_v_b_12')
// (18, 7, 'local_g3_3')
// (18, 7, 'lutff_global/cen')
// (18, 7, 'neigh_op_top_4')
// (18, 7, 'sp12_v_b_11')
// (18, 7, 'sp4_r_v_b_36')
// (18, 7, 'sp4_r_v_b_43')
// (18, 8, 'lutff_4/out')
// (18, 8, 'sp12_v_b_8')
// (18, 8, 'sp4_h_l_46')
// (18, 8, 'sp4_h_r_24')
// (18, 8, 'sp4_h_r_8')
// (18, 8, 'sp4_r_v_b_25')
// (18, 8, 'sp4_r_v_b_30')
// (18, 9, 'local_g3_3')
// (18, 9, 'lutff_global/cen')
// (18, 9, 'neigh_op_bot_4')
// (18, 9, 'sp12_v_b_7')
// (18, 9, 'sp4_r_v_b_12')
// (18, 9, 'sp4_r_v_b_19')
// (18, 10, 'sp12_v_b_4')
// (18, 10, 'sp4_r_v_b_1')
// (18, 10, 'sp4_r_v_b_6')
// (18, 11, 'sp12_v_b_3')
// (18, 12, 'sp12_v_b_0')
// (19, 6, 'sp4_v_t_36')
// (19, 6, 'sp4_v_t_43')
// (19, 7, 'neigh_op_tnl_4')
// (19, 7, 'sp4_v_b_36')
// (19, 7, 'sp4_v_b_43')
// (19, 8, 'neigh_op_lft_4')
// (19, 8, 'sp4_h_r_21')
// (19, 8, 'sp4_h_r_37')
// (19, 8, 'sp4_v_b_25')
// (19, 8, 'sp4_v_b_30')
// (19, 9, 'neigh_op_bnl_4')
// (19, 9, 'sp4_v_b_12')
// (19, 9, 'sp4_v_b_19')
// (19, 10, 'sp4_h_r_1')
// (19, 10, 'sp4_v_b_1')
// (19, 10, 'sp4_v_b_6')
// (20, 8, 'sp4_h_l_37')
// (20, 8, 'sp4_h_r_32')
// (20, 10, 'sp4_h_r_12')
// (21, 8, 'sp4_h_r_45')
// (21, 10, 'sp4_h_r_25')
// (22, 8, 'sp4_h_l_45')
// (22, 10, 'sp4_h_r_36')
// (23, 10, 'sp4_h_l_36')

wire n2077;
// (14, 8, 'neigh_op_tnr_0')
// (14, 9, 'neigh_op_rgt_0')
// (14, 10, 'neigh_op_bnr_0')
// (15, 8, 'neigh_op_top_0')
// (15, 9, 'lutff_0/out')
// (15, 10, 'local_g0_0')
// (15, 10, 'lutff_1/in_1')
// (15, 10, 'neigh_op_bot_0')
// (16, 8, 'neigh_op_tnl_0')
// (16, 9, 'neigh_op_lft_0')
// (16, 10, 'neigh_op_bnl_0')

wire n2078;
// (14, 8, 'neigh_op_tnr_1')
// (14, 9, 'neigh_op_rgt_1')
// (14, 10, 'neigh_op_bnr_1')
// (15, 8, 'neigh_op_top_1')
// (15, 9, 'local_g3_1')
// (15, 9, 'lutff_1/out')
// (15, 9, 'lutff_4/in_2')
// (15, 10, 'neigh_op_bot_1')
// (16, 8, 'neigh_op_tnl_1')
// (16, 9, 'neigh_op_lft_1')
// (16, 10, 'neigh_op_bnl_1')

wire n2079;
// (14, 8, 'neigh_op_tnr_2')
// (14, 9, 'neigh_op_rgt_2')
// (14, 10, 'neigh_op_bnr_2')
// (15, 8, 'neigh_op_top_2')
// (15, 9, 'local_g3_2')
// (15, 9, 'lutff_2/out')
// (15, 9, 'lutff_6/in_3')
// (15, 10, 'neigh_op_bot_2')
// (16, 8, 'neigh_op_tnl_2')
// (16, 9, 'neigh_op_lft_2')
// (16, 10, 'neigh_op_bnl_2')

reg n2080 = 0;
// (14, 8, 'neigh_op_tnr_3')
// (14, 9, 'neigh_op_rgt_3')
// (14, 10, 'neigh_op_bnr_3')
// (15, 8, 'neigh_op_top_3')
// (15, 9, 'lutff_3/out')
// (15, 10, 'neigh_op_bot_3')
// (16, 8, 'neigh_op_tnl_3')
// (16, 9, 'local_g1_3')
// (16, 9, 'lutff_6/in_2')
// (16, 9, 'neigh_op_lft_3')
// (16, 10, 'neigh_op_bnl_3')

wire n2081;
// (14, 8, 'neigh_op_tnr_4')
// (14, 9, 'neigh_op_rgt_4')
// (14, 10, 'neigh_op_bnr_4')
// (15, 8, 'neigh_op_top_4')
// (15, 9, 'lutff_4/out')
// (15, 10, 'local_g0_4')
// (15, 10, 'lutff_5/in_3')
// (15, 10, 'neigh_op_bot_4')
// (16, 8, 'neigh_op_tnl_4')
// (16, 9, 'neigh_op_lft_4')
// (16, 10, 'neigh_op_bnl_4')

wire n2082;
// (14, 8, 'neigh_op_tnr_5')
// (14, 9, 'neigh_op_rgt_5')
// (14, 10, 'neigh_op_bnr_5')
// (15, 8, 'neigh_op_top_5')
// (15, 9, 'local_g3_5')
// (15, 9, 'lutff_5/out')
// (15, 9, 'lutff_6/in_0')
// (15, 10, 'neigh_op_bot_5')
// (16, 8, 'neigh_op_tnl_5')
// (16, 9, 'neigh_op_lft_5')
// (16, 10, 'neigh_op_bnl_5')

wire n2083;
// (14, 8, 'neigh_op_tnr_6')
// (14, 9, 'neigh_op_rgt_6')
// (14, 10, 'neigh_op_bnr_6')
// (15, 8, 'neigh_op_top_6')
// (15, 9, 'local_g2_6')
// (15, 9, 'lutff_0/in_0')
// (15, 9, 'lutff_6/out')
// (15, 10, 'neigh_op_bot_6')
// (16, 8, 'neigh_op_tnl_6')
// (16, 9, 'neigh_op_lft_6')
// (16, 10, 'neigh_op_bnl_6')

wire n2084;
// (14, 8, 'neigh_op_tnr_7')
// (14, 9, 'neigh_op_rgt_7')
// (14, 10, 'neigh_op_bnr_7')
// (15, 8, 'neigh_op_top_7')
// (15, 9, 'local_g2_7')
// (15, 9, 'lutff_4/in_3')
// (15, 9, 'lutff_7/out')
// (15, 10, 'neigh_op_bot_7')
// (16, 8, 'neigh_op_tnl_7')
// (16, 9, 'neigh_op_lft_7')
// (16, 10, 'neigh_op_bnl_7')

reg n2085 = 0;
// (14, 9, 'neigh_op_tnr_0')
// (14, 10, 'neigh_op_rgt_0')
// (14, 11, 'neigh_op_bnr_0')
// (15, 8, 'sp4_r_v_b_41')
// (15, 9, 'neigh_op_top_0')
// (15, 9, 'sp4_r_v_b_28')
// (15, 10, 'lutff_0/out')
// (15, 10, 'sp4_r_v_b_17')
// (15, 11, 'neigh_op_bot_0')
// (15, 11, 'sp4_r_v_b_4')
// (16, 7, 'sp4_v_t_41')
// (16, 8, 'local_g2_1')
// (16, 8, 'lutff_1/in_0')
// (16, 8, 'sp4_v_b_41')
// (16, 9, 'local_g2_0')
// (16, 9, 'lutff_0/in_2')
// (16, 9, 'neigh_op_tnl_0')
// (16, 9, 'sp4_v_b_28')
// (16, 10, 'neigh_op_lft_0')
// (16, 10, 'sp4_v_b_17')
// (16, 11, 'neigh_op_bnl_0')
// (16, 11, 'sp4_v_b_4')

wire n2086;
// (14, 9, 'neigh_op_tnr_1')
// (14, 10, 'neigh_op_rgt_1')
// (14, 11, 'neigh_op_bnr_1')
// (15, 9, 'neigh_op_top_1')
// (15, 10, 'local_g2_1')
// (15, 10, 'lutff_1/out')
// (15, 10, 'lutff_2/in_3')
// (15, 11, 'neigh_op_bot_1')
// (16, 9, 'neigh_op_tnl_1')
// (16, 10, 'neigh_op_lft_1')
// (16, 11, 'neigh_op_bnl_1')

reg n2087 = 0;
// (14, 9, 'neigh_op_tnr_3')
// (14, 10, 'neigh_op_rgt_3')
// (14, 11, 'neigh_op_bnr_3')
// (15, 7, 'local_g3_2')
// (15, 7, 'lutff_4/in_3')
// (15, 7, 'sp4_r_v_b_42')
// (15, 8, 'sp4_r_v_b_31')
// (15, 9, 'neigh_op_top_3')
// (15, 9, 'sp4_r_v_b_18')
// (15, 10, 'lutff_3/out')
// (15, 10, 'sp4_r_v_b_7')
// (15, 11, 'neigh_op_bot_3')
// (16, 6, 'sp4_v_t_42')
// (16, 7, 'sp4_v_b_42')
// (16, 8, 'sp4_v_b_31')
// (16, 9, 'neigh_op_tnl_3')
// (16, 9, 'sp4_v_b_18')
// (16, 10, 'local_g0_3')
// (16, 10, 'lutff_7/in_0')
// (16, 10, 'neigh_op_lft_3')
// (16, 10, 'sp4_v_b_7')
// (16, 11, 'neigh_op_bnl_3')

wire n2088;
// (14, 9, 'neigh_op_tnr_4')
// (14, 10, 'neigh_op_rgt_4')
// (14, 11, 'neigh_op_bnr_4')
// (15, 9, 'neigh_op_top_4')
// (15, 10, 'local_g2_4')
// (15, 10, 'lutff_2/in_0')
// (15, 10, 'lutff_4/out')
// (15, 11, 'neigh_op_bot_4')
// (16, 9, 'neigh_op_tnl_4')
// (16, 10, 'neigh_op_lft_4')
// (16, 11, 'neigh_op_bnl_4')

wire n2089;
// (14, 9, 'neigh_op_tnr_5')
// (14, 10, 'neigh_op_rgt_5')
// (14, 11, 'neigh_op_bnr_5')
// (15, 9, 'neigh_op_top_5')
// (15, 10, 'local_g1_5')
// (15, 10, 'lutff_2/in_2')
// (15, 10, 'lutff_5/out')
// (15, 11, 'neigh_op_bot_5')
// (16, 9, 'neigh_op_tnl_5')
// (16, 10, 'neigh_op_lft_5')
// (16, 11, 'neigh_op_bnl_5')

reg n2090 = 0;
// (14, 9, 'neigh_op_tnr_6')
// (14, 10, 'neigh_op_rgt_6')
// (14, 11, 'neigh_op_bnr_6')
// (15, 9, 'neigh_op_top_6')
// (15, 10, 'local_g0_6')
// (15, 10, 'lutff_6/out')
// (15, 10, 'lutff_7/in_3')
// (15, 11, 'neigh_op_bot_6')
// (16, 9, 'neigh_op_tnl_6')
// (16, 10, 'local_g0_6')
// (16, 10, 'lutff_2/in_0')
// (16, 10, 'neigh_op_lft_6')
// (16, 11, 'neigh_op_bnl_6')

wire n2091;
// (14, 9, 'neigh_op_tnr_7')
// (14, 10, 'neigh_op_rgt_7')
// (14, 11, 'neigh_op_bnr_7')
// (15, 9, 'neigh_op_top_7')
// (15, 10, 'local_g1_7')
// (15, 10, 'lutff_4/in_2')
// (15, 10, 'lutff_7/out')
// (15, 11, 'neigh_op_bot_7')
// (16, 9, 'neigh_op_tnl_7')
// (16, 10, 'neigh_op_lft_7')
// (16, 11, 'neigh_op_bnl_7')

reg n2092 = 0;
// (14, 9, 'sp4_h_r_0')
// (15, 8, 'neigh_op_tnr_4')
// (15, 9, 'neigh_op_rgt_4')
// (15, 9, 'sp4_h_r_13')
// (15, 10, 'neigh_op_bnr_4')
// (16, 8, 'neigh_op_top_4')
// (16, 9, 'lutff_4/out')
// (16, 9, 'sp4_h_r_24')
// (16, 10, 'neigh_op_bot_4')
// (17, 8, 'neigh_op_tnl_4')
// (17, 9, 'neigh_op_lft_4')
// (17, 9, 'sp4_h_r_37')
// (17, 10, 'neigh_op_bnl_4')
// (17, 10, 'sp4_r_v_b_40')
// (17, 11, 'sp4_r_v_b_29')
// (17, 12, 'sp4_r_v_b_16')
// (17, 13, 'sp4_r_v_b_5')
// (18, 9, 'sp4_h_l_37')
// (18, 9, 'sp4_v_t_40')
// (18, 10, 'sp4_v_b_40')
// (18, 11, 'local_g3_5')
// (18, 11, 'lutff_2/in_2')
// (18, 11, 'sp4_v_b_29')
// (18, 12, 'sp4_v_b_16')
// (18, 13, 'sp4_v_b_5')

wire n2093;
// (14, 9, 'sp4_h_r_11')
// (15, 9, 'sp4_h_r_22')
// (16, 7, 'local_g0_2')
// (16, 7, 'lutff_global/cen')
// (16, 7, 'sp4_h_r_2')
// (16, 9, 'local_g3_3')
// (16, 9, 'lutff_global/cen')
// (16, 9, 'sp4_h_r_35')
// (17, 7, 'sp4_h_r_15')
// (17, 9, 'sp4_h_r_46')
// (18, 7, 'sp4_h_r_26')
// (18, 9, 'sp4_h_l_46')
// (18, 9, 'sp4_h_r_8')
// (19, 7, 'sp4_h_r_39')
// (19, 8, 'neigh_op_tnr_0')
// (19, 8, 'sp4_r_v_b_45')
// (19, 9, 'neigh_op_rgt_0')
// (19, 9, 'sp4_h_r_21')
// (19, 9, 'sp4_r_v_b_32')
// (19, 10, 'neigh_op_bnr_0')
// (19, 10, 'sp4_r_v_b_21')
// (19, 11, 'sp4_r_v_b_8')
// (20, 7, 'sp4_h_l_39')
// (20, 7, 'sp4_v_t_45')
// (20, 8, 'neigh_op_top_0')
// (20, 8, 'sp4_r_v_b_44')
// (20, 8, 'sp4_v_b_45')
// (20, 9, 'local_g0_2')
// (20, 9, 'lutff_0/out')
// (20, 9, 'lutff_global/cen')
// (20, 9, 'sp4_h_r_32')
// (20, 9, 'sp4_r_v_b_33')
// (20, 9, 'sp4_v_b_32')
// (20, 10, 'neigh_op_bot_0')
// (20, 10, 'sp4_r_v_b_20')
// (20, 10, 'sp4_v_b_21')
// (20, 11, 'sp4_r_v_b_9')
// (20, 11, 'sp4_v_b_8')
// (21, 7, 'sp4_v_t_44')
// (21, 8, 'neigh_op_tnl_0')
// (21, 8, 'sp4_v_b_44')
// (21, 9, 'neigh_op_lft_0')
// (21, 9, 'sp4_h_r_45')
// (21, 9, 'sp4_v_b_33')
// (21, 10, 'neigh_op_bnl_0')
// (21, 10, 'sp4_v_b_20')
// (21, 11, 'sp4_v_b_9')
// (22, 9, 'sp4_h_l_45')

wire n2094;
// (14, 10, 'neigh_op_tnr_0')
// (14, 11, 'neigh_op_rgt_0')
// (14, 12, 'neigh_op_bnr_0')
// (15, 10, 'neigh_op_top_0')
// (15, 11, 'lutff_0/out')
// (15, 12, 'local_g1_0')
// (15, 12, 'lutff_7/in_0')
// (15, 12, 'neigh_op_bot_0')
// (16, 10, 'neigh_op_tnl_0')
// (16, 11, 'neigh_op_lft_0')
// (16, 12, 'neigh_op_bnl_0')

wire n2095;
// (14, 10, 'neigh_op_tnr_1')
// (14, 11, 'neigh_op_rgt_1')
// (14, 12, 'neigh_op_bnr_1')
// (15, 10, 'neigh_op_top_1')
// (15, 11, 'local_g1_1')
// (15, 11, 'lutff_1/out')
// (15, 11, 'lutff_3/in_1')
// (15, 12, 'neigh_op_bot_1')
// (16, 10, 'neigh_op_tnl_1')
// (16, 11, 'neigh_op_lft_1')
// (16, 12, 'neigh_op_bnl_1')

wire n2096;
// (14, 10, 'neigh_op_tnr_2')
// (14, 11, 'neigh_op_rgt_2')
// (14, 12, 'neigh_op_bnr_2')
// (15, 10, 'neigh_op_top_2')
// (15, 11, 'lutff_2/out')
// (15, 12, 'local_g1_2')
// (15, 12, 'lutff_5/in_2')
// (15, 12, 'neigh_op_bot_2')
// (16, 10, 'neigh_op_tnl_2')
// (16, 11, 'neigh_op_lft_2')
// (16, 12, 'neigh_op_bnl_2')

wire n2097;
// (14, 10, 'neigh_op_tnr_3')
// (14, 11, 'local_g2_3')
// (14, 11, 'lutff_2/in_1')
// (14, 11, 'neigh_op_rgt_3')
// (14, 12, 'neigh_op_bnr_3')
// (15, 10, 'neigh_op_top_3')
// (15, 11, 'lutff_3/out')
// (15, 12, 'neigh_op_bot_3')
// (16, 10, 'neigh_op_tnl_3')
// (16, 11, 'neigh_op_lft_3')
// (16, 12, 'neigh_op_bnl_3')

wire n2098;
// (14, 10, 'neigh_op_tnr_4')
// (14, 11, 'neigh_op_rgt_4')
// (14, 12, 'neigh_op_bnr_4')
// (15, 10, 'local_g1_4')
// (15, 10, 'lutff_4/in_3')
// (15, 10, 'lutff_5/in_2')
// (15, 10, 'neigh_op_top_4')
// (15, 11, 'lutff_4/out')
// (15, 12, 'neigh_op_bot_4')
// (16, 10, 'neigh_op_tnl_4')
// (16, 11, 'neigh_op_lft_4')
// (16, 12, 'neigh_op_bnl_4')

reg n2099 = 0;
// (14, 10, 'neigh_op_tnr_5')
// (14, 11, 'neigh_op_rgt_5')
// (14, 12, 'neigh_op_bnr_5')
// (15, 10, 'neigh_op_top_5')
// (15, 11, 'lutff_5/out')
// (15, 12, 'neigh_op_bot_5')
// (16, 10, 'neigh_op_tnl_5')
// (16, 11, 'local_g1_5')
// (16, 11, 'lutff_6/in_0')
// (16, 11, 'neigh_op_lft_5')
// (16, 12, 'neigh_op_bnl_5')

wire n2100;
// (14, 10, 'neigh_op_tnr_6')
// (14, 11, 'neigh_op_rgt_6')
// (14, 12, 'local_g1_6')
// (14, 12, 'lutff_5/in_0')
// (14, 12, 'neigh_op_bnr_6')
// (15, 10, 'neigh_op_top_6')
// (15, 11, 'lutff_6/out')
// (15, 12, 'neigh_op_bot_6')
// (16, 10, 'neigh_op_tnl_6')
// (16, 11, 'neigh_op_lft_6')
// (16, 12, 'neigh_op_bnl_6')

reg n2101 = 0;
// (14, 10, 'neigh_op_tnr_7')
// (14, 11, 'neigh_op_rgt_7')
// (14, 12, 'neigh_op_bnr_7')
// (15, 10, 'neigh_op_top_7')
// (15, 11, 'lutff_7/out')
// (15, 12, 'neigh_op_bot_7')
// (16, 10, 'neigh_op_tnl_7')
// (16, 11, 'local_g1_7')
// (16, 11, 'lutff_5/in_1')
// (16, 11, 'neigh_op_lft_7')
// (16, 12, 'neigh_op_bnl_7')

wire n2102;
// (14, 10, 'sp4_r_v_b_45')
// (14, 11, 'local_g0_3')
// (14, 11, 'lutff_2/in_3')
// (14, 11, 'lutff_5/in_0')
// (14, 11, 'sp4_r_v_b_32')
// (14, 12, 'local_g2_4')
// (14, 12, 'lutff_0/in_0')
// (14, 12, 'lutff_1/in_1')
// (14, 12, 'lutff_2/in_0')
// (14, 12, 'lutff_5/in_1')
// (14, 12, 'neigh_op_tnr_4')
// (14, 12, 'sp4_r_v_b_21')
// (14, 13, 'local_g2_4')
// (14, 13, 'lutff_3/in_1')
// (14, 13, 'neigh_op_rgt_4')
// (14, 13, 'sp4_r_v_b_8')
// (14, 14, 'local_g1_4')
// (14, 14, 'lutff_5/in_2')
// (14, 14, 'lutff_6/in_1')
// (14, 14, 'neigh_op_bnr_4')
// (15, 9, 'sp4_v_t_45')
// (15, 10, 'sp4_v_b_45')
// (15, 11, 'sp4_v_b_32')
// (15, 12, 'local_g0_4')
// (15, 12, 'lutff_2/in_0')
// (15, 12, 'neigh_op_top_4')
// (15, 12, 'sp4_v_b_21')
// (15, 13, 'local_g2_4')
// (15, 13, 'lutff_0/in_0')
// (15, 13, 'lutff_2/in_2')
// (15, 13, 'lutff_4/out')
// (15, 13, 'sp4_v_b_8')
// (15, 14, 'neigh_op_bot_4')
// (16, 12, 'neigh_op_tnl_4')
// (16, 13, 'neigh_op_lft_4')
// (16, 14, 'neigh_op_bnl_4')

wire n2103;
// (14, 10, 'sp4_r_v_b_46')
// (14, 11, 'neigh_op_tnr_3')
// (14, 11, 'sp4_r_v_b_35')
// (14, 12, 'neigh_op_rgt_3')
// (14, 12, 'sp4_r_v_b_22')
// (14, 13, 'neigh_op_bnr_3')
// (14, 13, 'sp4_r_v_b_11')
// (15, 9, 'sp4_v_t_46')
// (15, 10, 'sp4_v_b_46')
// (15, 11, 'local_g1_3')
// (15, 11, 'local_g2_3')
// (15, 11, 'lutff_3/in_0')
// (15, 11, 'lutff_6/in_2')
// (15, 11, 'neigh_op_top_3')
// (15, 11, 'sp4_v_b_35')
// (15, 12, 'lutff_3/out')
// (15, 12, 'sp4_v_b_22')
// (15, 13, 'neigh_op_bot_3')
// (15, 13, 'sp4_v_b_11')
// (16, 11, 'neigh_op_tnl_3')
// (16, 12, 'local_g1_3')
// (16, 12, 'lutff_5/in_3')
// (16, 12, 'neigh_op_lft_3')
// (16, 13, 'neigh_op_bnl_3')

wire n2104;
// (14, 11, 'local_g3_7')
// (14, 11, 'lutff_5/in_3')
// (14, 11, 'sp4_r_v_b_47')
// (14, 12, 'local_g0_1')
// (14, 12, 'lutff_1/in_2')
// (14, 12, 'lutff_5/in_2')
// (14, 12, 'sp4_r_v_b_34')
// (14, 13, 'neigh_op_tnr_5')
// (14, 13, 'sp4_r_v_b_23')
// (14, 14, 'neigh_op_rgt_5')
// (14, 14, 'sp4_r_v_b_10')
// (14, 15, 'neigh_op_bnr_5')
// (15, 10, 'sp4_v_t_47')
// (15, 11, 'sp4_v_b_47')
// (15, 12, 'local_g3_2')
// (15, 12, 'lutff_2/in_1')
// (15, 12, 'lutff_3/in_0')
// (15, 12, 'sp4_v_b_34')
// (15, 13, 'local_g0_5')
// (15, 13, 'lutff_0/in_3')
// (15, 13, 'lutff_2/in_3')
// (15, 13, 'neigh_op_top_5')
// (15, 13, 'sp4_v_b_23')
// (15, 14, 'lutff_5/out')
// (15, 14, 'sp4_v_b_10')
// (15, 15, 'neigh_op_bot_5')
// (16, 13, 'neigh_op_tnl_5')
// (16, 14, 'neigh_op_lft_5')
// (16, 15, 'neigh_op_bnl_5')

wire n2105;
// (14, 11, 'neigh_op_tnr_0')
// (14, 12, 'local_g2_0')
// (14, 12, 'lutff_7/in_3')
// (14, 12, 'neigh_op_rgt_0')
// (14, 13, 'neigh_op_bnr_0')
// (15, 11, 'neigh_op_top_0')
// (15, 12, 'lutff_0/out')
// (15, 13, 'neigh_op_bot_0')
// (16, 11, 'neigh_op_tnl_0')
// (16, 12, 'neigh_op_lft_0')
// (16, 13, 'neigh_op_bnl_0')

wire n2106;
// (14, 11, 'neigh_op_tnr_1')
// (14, 12, 'neigh_op_rgt_1')
// (14, 13, 'neigh_op_bnr_1')
// (15, 11, 'neigh_op_top_1')
// (15, 12, 'local_g1_1')
// (15, 12, 'lutff_0/in_0')
// (15, 12, 'lutff_1/out')
// (15, 13, 'neigh_op_bot_1')
// (16, 11, 'neigh_op_tnl_1')
// (16, 12, 'neigh_op_lft_1')
// (16, 13, 'neigh_op_bnl_1')

wire n2107;
// (14, 11, 'neigh_op_tnr_4')
// (14, 12, 'neigh_op_rgt_4')
// (14, 13, 'local_g0_4')
// (14, 13, 'lutff_1/in_3')
// (14, 13, 'neigh_op_bnr_4')
// (15, 11, 'neigh_op_top_4')
// (15, 12, 'lutff_4/out')
// (15, 13, 'neigh_op_bot_4')
// (16, 11, 'neigh_op_tnl_4')
// (16, 12, 'neigh_op_lft_4')
// (16, 13, 'neigh_op_bnl_4')

wire n2108;
// (14, 11, 'neigh_op_tnr_5')
// (14, 12, 'neigh_op_rgt_5')
// (14, 13, 'local_g1_5')
// (14, 13, 'lutff_2/in_0')
// (14, 13, 'neigh_op_bnr_5')
// (15, 11, 'neigh_op_top_5')
// (15, 12, 'lutff_5/out')
// (15, 13, 'neigh_op_bot_5')
// (16, 11, 'neigh_op_tnl_5')
// (16, 12, 'neigh_op_lft_5')
// (16, 13, 'neigh_op_bnl_5')

wire n2109;
// (14, 11, 'neigh_op_tnr_7')
// (14, 12, 'neigh_op_rgt_7')
// (14, 13, 'neigh_op_bnr_7')
// (15, 11, 'neigh_op_top_7')
// (15, 12, 'lutff_7/out')
// (15, 13, 'local_g0_7')
// (15, 13, 'lutff_6/in_3')
// (15, 13, 'neigh_op_bot_7')
// (16, 11, 'neigh_op_tnl_7')
// (16, 12, 'neigh_op_lft_7')
// (16, 13, 'neigh_op_bnl_7')

wire n2110;
// (14, 11, 'sp4_h_r_8')
// (15, 10, 'neigh_op_tnr_0')
// (15, 11, 'local_g0_5')
// (15, 11, 'lutff_6/in_1')
// (15, 11, 'neigh_op_rgt_0')
// (15, 11, 'sp4_h_r_21')
// (15, 12, 'neigh_op_bnr_0')
// (16, 10, 'neigh_op_top_0')
// (16, 11, 'lutff_0/out')
// (16, 11, 'sp4_h_r_32')
// (16, 12, 'neigh_op_bot_0')
// (17, 10, 'neigh_op_tnl_0')
// (17, 11, 'neigh_op_lft_0')
// (17, 11, 'sp4_h_r_45')
// (17, 12, 'neigh_op_bnl_0')
// (18, 11, 'sp4_h_l_45')

wire n2111;
// (14, 11, 'sp4_h_r_9')
// (15, 11, 'sp4_h_r_20')
// (16, 10, 'neigh_op_tnr_6')
// (16, 11, 'local_g2_1')
// (16, 11, 'lutff_3/in_2')
// (16, 11, 'neigh_op_rgt_6')
// (16, 11, 'sp4_h_r_33')
// (16, 12, 'neigh_op_bnr_6')
// (17, 10, 'neigh_op_top_6')
// (17, 11, 'lutff_6/out')
// (17, 11, 'sp4_h_r_44')
// (17, 12, 'neigh_op_bot_6')
// (18, 10, 'neigh_op_tnl_6')
// (18, 11, 'neigh_op_lft_6')
// (18, 11, 'sp4_h_l_44')
// (18, 12, 'neigh_op_bnl_6')

wire n2112;
// (14, 11, 'sp4_r_v_b_42')
// (14, 12, 'sp4_r_v_b_31')
// (14, 13, 'sp4_r_v_b_18')
// (14, 14, 'sp4_r_v_b_7')
// (15, 10, 'sp4_h_r_7')
// (15, 10, 'sp4_v_t_42')
// (15, 11, 'local_g2_2')
// (15, 11, 'lutff_global/cen')
// (15, 11, 'sp4_v_b_42')
// (15, 12, 'sp4_v_b_31')
// (15, 13, 'sp4_v_b_18')
// (15, 14, 'sp4_v_b_7')
// (16, 10, 'local_g0_2')
// (16, 10, 'lutff_global/cen')
// (16, 10, 'sp4_h_r_18')
// (17, 10, 'sp4_h_r_31')
// (18, 10, 'sp4_h_r_42')
// (19, 9, 'neigh_op_tnr_1')
// (19, 9, 'sp4_r_v_b_47')
// (19, 10, 'neigh_op_rgt_1')
// (19, 10, 'sp4_h_l_42')
// (19, 10, 'sp4_h_r_7')
// (19, 10, 'sp4_r_v_b_34')
// (19, 11, 'neigh_op_bnr_1')
// (19, 11, 'sp4_r_v_b_23')
// (19, 12, 'sp4_r_v_b_10')
// (20, 8, 'sp4_v_t_47')
// (20, 9, 'neigh_op_top_1')
// (20, 9, 'sp4_v_b_47')
// (20, 10, 'local_g0_2')
// (20, 10, 'lutff_1/out')
// (20, 10, 'lutff_global/cen')
// (20, 10, 'sp4_h_r_18')
// (20, 10, 'sp4_v_b_34')
// (20, 11, 'neigh_op_bot_1')
// (20, 11, 'sp4_v_b_23')
// (20, 12, 'local_g0_2')
// (20, 12, 'lutff_global/cen')
// (20, 12, 'sp4_v_b_10')
// (21, 9, 'neigh_op_tnl_1')
// (21, 10, 'neigh_op_lft_1')
// (21, 10, 'sp4_h_r_31')
// (21, 11, 'neigh_op_bnl_1')
// (22, 10, 'sp4_h_r_42')
// (23, 10, 'sp4_h_l_42')

wire n2113;
// (14, 11, 'sp4_r_v_b_44')
// (14, 12, 'sp4_r_v_b_33')
// (14, 13, 'sp4_r_v_b_20')
// (14, 14, 'sp4_r_v_b_9')
// (15, 10, 'sp4_h_r_3')
// (15, 10, 'sp4_v_t_44')
// (15, 11, 'sp4_v_b_44')
// (15, 12, 'sp4_v_b_33')
// (15, 13, 'sp4_v_b_20')
// (15, 14, 'local_g1_1')
// (15, 14, 'lutff_1/in_1')
// (15, 14, 'lutff_2/in_2')
// (15, 14, 'sp4_v_b_9')
// (16, 10, 'sp4_h_r_14')
// (17, 10, 'sp4_h_r_27')
// (17, 10, 'sp4_r_v_b_45')
// (17, 11, 'sp4_r_v_b_32')
// (17, 12, 'local_g3_5')
// (17, 12, 'lutff_1/in_3')
// (17, 12, 'sp4_r_v_b_21')
// (17, 13, 'sp4_r_v_b_8')
// (18, 9, 'sp4_v_t_45')
// (18, 10, 'sp4_h_r_38')
// (18, 10, 'sp4_v_b_45')
// (18, 11, 'sp4_v_b_32')
// (18, 12, 'sp4_v_b_21')
// (18, 13, 'sp4_h_r_3')
// (18, 13, 'sp4_v_b_8')
// (19, 10, 'sp4_h_l_38')
// (19, 10, 'sp4_h_r_3')
// (19, 13, 'sp4_h_r_14')
// (20, 10, 'sp4_h_r_14')
// (20, 13, 'sp4_h_r_27')
// (21, 9, 'neigh_op_tnr_3')
// (21, 10, 'neigh_op_rgt_3')
// (21, 10, 'sp4_h_r_27')
// (21, 10, 'sp4_r_v_b_38')
// (21, 11, 'neigh_op_bnr_3')
// (21, 11, 'sp4_r_v_b_27')
// (21, 12, 'sp4_r_v_b_14')
// (21, 13, 'sp4_h_r_38')
// (21, 13, 'sp4_r_v_b_3')
// (22, 9, 'neigh_op_top_3')
// (22, 9, 'sp4_v_t_38')
// (22, 10, 'local_g3_3')
// (22, 10, 'lutff_3/out')
// (22, 10, 'lutff_global/cen')
// (22, 10, 'sp4_h_r_38')
// (22, 10, 'sp4_v_b_38')
// (22, 11, 'neigh_op_bot_3')
// (22, 11, 'sp4_v_b_27')
// (22, 12, 'sp4_v_b_14')
// (22, 13, 'sp4_h_l_38')
// (22, 13, 'sp4_v_b_3')
// (23, 9, 'neigh_op_tnl_3')
// (23, 10, 'neigh_op_lft_3')
// (23, 10, 'sp4_h_l_38')
// (23, 11, 'neigh_op_bnl_3')

wire n2114;
// (14, 12, 'neigh_op_tnr_0')
// (14, 13, 'local_g3_0')
// (14, 13, 'lutff_2/in_3')
// (14, 13, 'neigh_op_rgt_0')
// (14, 14, 'neigh_op_bnr_0')
// (15, 12, 'neigh_op_top_0')
// (15, 13, 'lutff_0/out')
// (15, 14, 'neigh_op_bot_0')
// (16, 12, 'neigh_op_tnl_0')
// (16, 13, 'neigh_op_lft_0')
// (16, 14, 'neigh_op_bnl_0')

wire n2115;
// (14, 12, 'neigh_op_tnr_1')
// (14, 13, 'neigh_op_rgt_1')
// (14, 14, 'neigh_op_bnr_1')
// (15, 12, 'neigh_op_top_1')
// (15, 13, 'local_g1_1')
// (15, 13, 'lutff_1/out')
// (15, 13, 'lutff_5/in_1')
// (15, 14, 'neigh_op_bot_1')
// (16, 12, 'neigh_op_tnl_1')
// (16, 13, 'neigh_op_lft_1')
// (16, 14, 'neigh_op_bnl_1')

wire n2116;
// (14, 12, 'neigh_op_tnr_2')
// (14, 13, 'neigh_op_rgt_2')
// (14, 14, 'neigh_op_bnr_2')
// (15, 12, 'local_g0_2')
// (15, 12, 'lutff_0/in_2')
// (15, 12, 'neigh_op_top_2')
// (15, 13, 'local_g2_2')
// (15, 13, 'lutff_1/in_1')
// (15, 13, 'lutff_2/out')
// (15, 14, 'local_g0_2')
// (15, 14, 'local_g1_2')
// (15, 14, 'lutff_3/in_3')
// (15, 14, 'lutff_6/in_1')
// (15, 14, 'neigh_op_bot_2')
// (16, 12, 'neigh_op_tnl_2')
// (16, 13, 'neigh_op_lft_2')
// (16, 14, 'neigh_op_bnl_2')

wire n2117;
// (14, 12, 'neigh_op_tnr_3')
// (14, 13, 'neigh_op_rgt_3')
// (14, 14, 'neigh_op_bnr_3')
// (15, 12, 'local_g0_3')
// (15, 12, 'lutff_0/in_1')
// (15, 12, 'lutff_1/in_2')
// (15, 12, 'lutff_3/in_2')
// (15, 12, 'neigh_op_top_3')
// (15, 13, 'local_g1_3')
// (15, 13, 'lutff_1/in_3')
// (15, 13, 'lutff_3/out')
// (15, 13, 'lutff_5/in_3')
// (15, 14, 'local_g0_3')
// (15, 14, 'lutff_0/in_1')
// (15, 14, 'lutff_6/in_3')
// (15, 14, 'lutff_7/in_0')
// (15, 14, 'neigh_op_bot_3')
// (16, 12, 'neigh_op_tnl_3')
// (16, 13, 'neigh_op_lft_3')
// (16, 14, 'neigh_op_bnl_3')

wire n2118;
// (14, 12, 'neigh_op_tnr_5')
// (14, 13, 'neigh_op_rgt_5')
// (14, 14, 'local_g0_5')
// (14, 14, 'lutff_1/in_0')
// (14, 14, 'neigh_op_bnr_5')
// (15, 12, 'neigh_op_top_5')
// (15, 13, 'lutff_5/out')
// (15, 14, 'neigh_op_bot_5')
// (16, 12, 'neigh_op_tnl_5')
// (16, 13, 'neigh_op_lft_5')
// (16, 14, 'neigh_op_bnl_5')

wire n2119;
// (14, 12, 'neigh_op_tnr_6')
// (14, 13, 'local_g3_6')
// (14, 13, 'lutff_5/in_2')
// (14, 13, 'neigh_op_rgt_6')
// (14, 14, 'neigh_op_bnr_6')
// (15, 12, 'neigh_op_top_6')
// (15, 13, 'lutff_6/out')
// (15, 14, 'neigh_op_bot_6')
// (16, 12, 'neigh_op_tnl_6')
// (16, 13, 'neigh_op_lft_6')
// (16, 14, 'neigh_op_bnl_6')

wire n2120;
// (14, 12, 'sp4_h_r_11')
// (15, 12, 'sp4_h_r_22')
// (16, 12, 'local_g3_3')
// (16, 12, 'lutff_global/cen')
// (16, 12, 'sp4_h_r_35')
// (17, 7, 'neigh_op_tnr_3')
// (17, 8, 'neigh_op_rgt_3')
// (17, 9, 'neigh_op_bnr_3')
// (17, 9, 'sp4_r_v_b_43')
// (17, 10, 'sp4_r_v_b_30')
// (17, 11, 'sp4_r_v_b_19')
// (17, 12, 'sp4_h_r_46')
// (17, 12, 'sp4_r_v_b_6')
// (18, 0, 'span12_vert_21')
// (18, 1, 'sp12_v_b_21')
// (18, 2, 'sp12_v_b_18')
// (18, 3, 'sp12_v_b_17')
// (18, 4, 'sp12_v_b_14')
// (18, 5, 'sp12_v_b_13')
// (18, 6, 'sp12_v_b_10')
// (18, 7, 'neigh_op_top_3')
// (18, 7, 'sp12_v_b_9')
// (18, 8, 'local_g1_3')
// (18, 8, 'lutff_3/out')
// (18, 8, 'lutff_global/cen')
// (18, 8, 'sp12_v_b_6')
// (18, 8, 'sp4_h_r_6')
// (18, 8, 'sp4_v_t_43')
// (18, 9, 'neigh_op_bot_3')
// (18, 9, 'sp12_v_b_5')
// (18, 9, 'sp4_v_b_43')
// (18, 10, 'local_g2_2')
// (18, 10, 'lutff_global/cen')
// (18, 10, 'sp12_v_b_2')
// (18, 10, 'sp4_v_b_30')
// (18, 11, 'sp12_v_b_1')
// (18, 11, 'sp4_v_b_19')
// (18, 12, 'sp4_h_l_46')
// (18, 12, 'sp4_v_b_6')
// (19, 7, 'neigh_op_tnl_3')
// (19, 8, 'neigh_op_lft_3')
// (19, 8, 'sp4_h_r_19')
// (19, 9, 'neigh_op_bnl_3')
// (20, 8, 'sp4_h_r_30')
// (21, 8, 'sp4_h_r_43')
// (22, 8, 'sp4_h_l_43')

wire n2121;
// (14, 12, 'sp4_r_v_b_45')
// (14, 13, 'sp4_r_v_b_32')
// (14, 14, 'neigh_op_tnr_4')
// (14, 14, 'sp4_r_v_b_21')
// (14, 15, 'neigh_op_rgt_4')
// (14, 15, 'sp4_r_v_b_8')
// (14, 16, 'neigh_op_bnr_4')
// (15, 11, 'sp4_v_t_45')
// (15, 12, 'sp4_v_b_45')
// (15, 13, 'local_g2_0')
// (15, 13, 'lutff_4/in_0')
// (15, 13, 'sp4_v_b_32')
// (15, 14, 'neigh_op_top_4')
// (15, 14, 'sp4_v_b_21')
// (15, 15, 'lutff_4/out')
// (15, 15, 'sp4_v_b_8')
// (15, 16, 'neigh_op_bot_4')
// (16, 14, 'neigh_op_tnl_4')
// (16, 15, 'neigh_op_lft_4')
// (16, 16, 'neigh_op_bnl_4')

wire n2122;
// (14, 13, 'local_g1_6')
// (14, 13, 'lutff_2/in_1')
// (14, 13, 'sp4_h_r_6')
// (15, 12, 'local_g2_7')
// (15, 12, 'lutff_7/in_2')
// (15, 12, 'neigh_op_tnr_7')
// (15, 13, 'local_g2_7')
// (15, 13, 'lutff_3/in_0')
// (15, 13, 'lutff_5/in_2')
// (15, 13, 'neigh_op_rgt_7')
// (15, 13, 'sp4_h_r_19')
// (15, 14, 'local_g0_7')
// (15, 14, 'lutff_3/in_0')
// (15, 14, 'neigh_op_bnr_7')
// (16, 12, 'local_g0_7')
// (16, 12, 'lutff_2/in_1')
// (16, 12, 'neigh_op_top_7')
// (16, 13, 'local_g0_7')
// (16, 13, 'lutff_0/in_1')
// (16, 13, 'lutff_7/out')
// (16, 13, 'sp4_h_r_30')
// (16, 14, 'neigh_op_bot_7')
// (17, 12, 'neigh_op_tnl_7')
// (17, 13, 'neigh_op_lft_7')
// (17, 13, 'sp4_h_r_43')
// (17, 14, 'neigh_op_bnl_7')
// (18, 13, 'sp4_h_l_43')

wire n2123;
// (14, 13, 'local_g2_6')
// (14, 13, 'lutff_2/in_2')
// (14, 13, 'neigh_op_tnr_6')
// (14, 14, 'neigh_op_rgt_6')
// (14, 15, 'neigh_op_bnr_6')
// (15, 13, 'neigh_op_top_6')
// (15, 14, 'lutff_6/out')
// (15, 15, 'neigh_op_bot_6')
// (16, 13, 'neigh_op_tnl_6')
// (16, 14, 'neigh_op_lft_6')
// (16, 15, 'neigh_op_bnl_6')

wire n2124;
// (14, 13, 'neigh_op_tnr_0')
// (14, 14, 'local_g2_0')
// (14, 14, 'lutff_4/in_0')
// (14, 14, 'neigh_op_rgt_0')
// (14, 15, 'neigh_op_bnr_0')
// (15, 13, 'neigh_op_top_0')
// (15, 14, 'lutff_0/out')
// (15, 15, 'neigh_op_bot_0')
// (16, 13, 'neigh_op_tnl_0')
// (16, 14, 'neigh_op_lft_0')
// (16, 15, 'neigh_op_bnl_0')

reg n2125 = 0;
// (14, 13, 'neigh_op_tnr_2')
// (14, 14, 'neigh_op_rgt_2')
// (14, 15, 'neigh_op_bnr_2')
// (15, 13, 'neigh_op_top_2')
// (15, 14, 'lutff_2/out')
// (15, 14, 'sp4_r_v_b_37')
// (15, 15, 'neigh_op_bot_2')
// (15, 15, 'sp4_r_v_b_24')
// (15, 16, 'sp4_r_v_b_13')
// (15, 17, 'sp4_r_v_b_0')
// (16, 13, 'neigh_op_tnl_2')
// (16, 13, 'sp4_v_t_37')
// (16, 14, 'neigh_op_lft_2')
// (16, 14, 'sp4_v_b_37')
// (16, 15, 'neigh_op_bnl_2')
// (16, 15, 'sp4_v_b_24')
// (16, 16, 'local_g1_5')
// (16, 16, 'lutff_7/in_1')
// (16, 16, 'sp4_v_b_13')
// (16, 17, 'sp4_v_b_0')

wire n2126;
// (14, 13, 'neigh_op_tnr_3')
// (14, 14, 'local_g2_3')
// (14, 14, 'lutff_4/in_3')
// (14, 14, 'neigh_op_rgt_3')
// (14, 15, 'neigh_op_bnr_3')
// (15, 13, 'neigh_op_top_3')
// (15, 14, 'local_g3_3')
// (15, 14, 'lutff_3/out')
// (15, 14, 'lutff_7/in_3')
// (15, 15, 'neigh_op_bot_3')
// (16, 13, 'neigh_op_tnl_3')
// (16, 14, 'neigh_op_lft_3')
// (16, 15, 'neigh_op_bnl_3')

wire n2127;
// (14, 13, 'neigh_op_tnr_7')
// (14, 14, 'neigh_op_rgt_7')
// (14, 15, 'neigh_op_bnr_7')
// (15, 13, 'local_g1_7')
// (15, 13, 'lutff_6/in_0')
// (15, 13, 'neigh_op_top_7')
// (15, 14, 'lutff_7/out')
// (15, 15, 'neigh_op_bot_7')
// (16, 13, 'neigh_op_tnl_7')
// (16, 14, 'neigh_op_lft_7')
// (16, 15, 'neigh_op_bnl_7')

reg n2128 = 0;
// (14, 13, 'sp4_r_v_b_41')
// (14, 14, 'local_g0_4')
// (14, 14, 'lutff_3/in_3')
// (14, 14, 'sp4_r_v_b_28')
// (14, 15, 'neigh_op_tnr_2')
// (14, 15, 'sp4_r_v_b_17')
// (14, 16, 'local_g3_2')
// (14, 16, 'lutff_3/in_2')
// (14, 16, 'neigh_op_rgt_2')
// (14, 16, 'sp4_r_v_b_4')
// (14, 17, 'neigh_op_bnr_2')
// (15, 12, 'sp4_v_t_41')
// (15, 13, 'sp4_v_b_41')
// (15, 14, 'sp4_r_v_b_45')
// (15, 14, 'sp4_v_b_28')
// (15, 15, 'local_g1_2')
// (15, 15, 'lutff_3/in_0')
// (15, 15, 'lutff_4/in_1')
// (15, 15, 'neigh_op_top_2')
// (15, 15, 'sp4_r_v_b_32')
// (15, 15, 'sp4_v_b_17')
// (15, 16, 'local_g2_2')
// (15, 16, 'lutff_2/in_2')
// (15, 16, 'lutff_2/out')
// (15, 16, 'sp4_r_v_b_21')
// (15, 16, 'sp4_v_b_4')
// (15, 17, 'neigh_op_bot_2')
// (15, 17, 'sp4_r_v_b_8')
// (16, 13, 'sp4_v_t_45')
// (16, 14, 'local_g2_5')
// (16, 14, 'lutff_0/in_1')
// (16, 14, 'lutff_4/in_1')
// (16, 14, 'lutff_6/in_1')
// (16, 14, 'sp4_v_b_45')
// (16, 15, 'neigh_op_tnl_2')
// (16, 15, 'sp4_v_b_32')
// (16, 16, 'neigh_op_lft_2')
// (16, 16, 'sp4_v_b_21')
// (16, 17, 'neigh_op_bnl_2')
// (16, 17, 'sp4_v_b_8')

wire n2129;
// (14, 14, 'local_g3_3')
// (14, 14, 'lutff_3/in_1')
// (14, 14, 'neigh_op_tnr_3')
// (14, 15, 'neigh_op_rgt_3')
// (14, 16, 'neigh_op_bnr_3')
// (15, 14, 'local_g1_3')
// (15, 14, 'lutff_5/in_3')
// (15, 14, 'neigh_op_top_3')
// (15, 15, 'lutff_3/out')
// (15, 16, 'neigh_op_bot_3')
// (16, 14, 'local_g2_3')
// (16, 14, 'local_g3_3')
// (16, 14, 'lutff_4/in_2')
// (16, 14, 'lutff_5/in_2')
// (16, 14, 'neigh_op_tnl_3')
// (16, 15, 'neigh_op_lft_3')
// (16, 16, 'neigh_op_bnl_3')

wire n2130;
// (14, 14, 'neigh_op_tnr_5')
// (14, 15, 'neigh_op_rgt_5')
// (14, 16, 'neigh_op_bnr_5')
// (15, 14, 'neigh_op_top_5')
// (15, 15, 'local_g3_5')
// (15, 15, 'lutff_3/in_1')
// (15, 15, 'lutff_5/out')
// (15, 16, 'neigh_op_bot_5')
// (16, 14, 'neigh_op_tnl_5')
// (16, 15, 'neigh_op_lft_5')
// (16, 16, 'neigh_op_bnl_5')

reg n2131 = 0;
// (14, 14, 'neigh_op_tnr_6')
// (14, 15, 'neigh_op_rgt_6')
// (14, 16, 'neigh_op_bnr_6')
// (15, 14, 'neigh_op_top_6')
// (15, 15, 'lutff_6/out')
// (15, 16, 'neigh_op_bot_6')
// (16, 14, 'neigh_op_tnl_6')
// (16, 15, 'local_g0_6')
// (16, 15, 'lutff_2/in_0')
// (16, 15, 'neigh_op_lft_6')
// (16, 16, 'neigh_op_bnl_6')

reg n2132 = 0;
// (14, 14, 'neigh_op_tnr_7')
// (14, 15, 'neigh_op_rgt_7')
// (14, 16, 'neigh_op_bnr_7')
// (15, 14, 'neigh_op_top_7')
// (15, 15, 'lutff_7/out')
// (15, 16, 'neigh_op_bot_7')
// (16, 14, 'neigh_op_tnl_7')
// (16, 15, 'local_g0_7')
// (16, 15, 'lutff_7/in_0')
// (16, 15, 'neigh_op_lft_7')
// (16, 16, 'neigh_op_bnl_7')

wire n2133;
// (14, 14, 'sp12_h_r_0')
// (15, 14, 'sp12_h_r_3')
// (16, 14, 'sp12_h_r_4')
// (17, 13, 'neigh_op_tnr_0')
// (17, 14, 'neigh_op_rgt_0')
// (17, 14, 'sp12_h_r_7')
// (17, 15, 'neigh_op_bnr_0')
// (18, 8, 'sp4_r_v_b_42')
// (18, 9, 'sp4_r_v_b_31')
// (18, 10, 'sp4_r_v_b_18')
// (18, 11, 'sp4_r_v_b_7')
// (18, 12, 'sp4_r_v_b_41')
// (18, 13, 'neigh_op_top_0')
// (18, 13, 'sp4_r_v_b_28')
// (18, 13, 'sp4_r_v_b_44')
// (18, 14, 'lutff_0/out')
// (18, 14, 'sp12_h_r_8')
// (18, 14, 'sp4_r_v_b_17')
// (18, 14, 'sp4_r_v_b_33')
// (18, 15, 'neigh_op_bot_0')
// (18, 15, 'sp4_r_v_b_20')
// (18, 15, 'sp4_r_v_b_4')
// (18, 16, 'sp4_r_v_b_9')
// (19, 7, 'sp4_v_t_42')
// (19, 8, 'sp4_v_b_42')
// (19, 9, 'sp4_v_b_31')
// (19, 10, 'local_g0_2')
// (19, 10, 'ram/WCLKE')
// (19, 10, 'sp4_v_b_18')
// (19, 11, 'sp4_v_b_7')
// (19, 11, 'sp4_v_t_41')
// (19, 12, 'local_g0_2')
// (19, 12, 'ram/WCLKE')
// (19, 12, 'sp4_h_r_2')
// (19, 12, 'sp4_v_b_41')
// (19, 12, 'sp4_v_t_44')
// (19, 13, 'neigh_op_tnl_0')
// (19, 13, 'sp4_v_b_28')
// (19, 13, 'sp4_v_b_44')
// (19, 14, 'local_g1_3')
// (19, 14, 'neigh_op_lft_0')
// (19, 14, 'ram/WCLKE')
// (19, 14, 'sp12_h_r_11')
// (19, 14, 'sp4_v_b_17')
// (19, 14, 'sp4_v_b_33')
// (19, 15, 'neigh_op_bnl_0')
// (19, 15, 'sp4_v_b_20')
// (19, 15, 'sp4_v_b_4')
// (19, 16, 'sp4_v_b_9')
// (20, 12, 'local_g0_7')
// (20, 12, 'lutff_3/in_0')
// (20, 12, 'sp4_h_r_15')
// (20, 14, 'sp12_h_r_12')
// (21, 12, 'sp4_h_r_26')
// (21, 14, 'sp12_h_r_15')
// (22, 12, 'sp4_h_r_39')
// (22, 14, 'sp12_h_r_16')
// (23, 12, 'sp4_h_l_39')
// (23, 14, 'sp12_h_r_19')
// (24, 14, 'sp12_h_r_20')
// (25, 14, 'sp12_h_r_23')

wire n2134;
// (14, 14, 'sp4_r_v_b_47')
// (14, 15, 'sp4_r_v_b_34')
// (14, 16, 'neigh_op_tnr_5')
// (14, 16, 'sp4_r_v_b_23')
// (14, 17, 'neigh_op_rgt_5')
// (14, 17, 'sp4_r_v_b_10')
// (14, 18, 'neigh_op_bnr_5')
// (15, 10, 'sp12_v_t_22')
// (15, 11, 'sp12_v_b_22')
// (15, 12, 'sp12_v_b_21')
// (15, 13, 'sp12_v_b_18')
// (15, 13, 'sp4_v_t_47')
// (15, 14, 'sp12_v_b_17')
// (15, 14, 'sp4_v_b_47')
// (15, 15, 'local_g2_2')
// (15, 15, 'lutff_6/in_0')
// (15, 15, 'sp12_v_b_14')
// (15, 15, 'sp4_v_b_34')
// (15, 16, 'neigh_op_top_5')
// (15, 16, 'sp12_v_b_13')
// (15, 16, 'sp4_v_b_23')
// (15, 17, 'lutff_5/out')
// (15, 17, 'sp12_v_b_10')
// (15, 17, 'sp4_v_b_10')
// (15, 18, 'neigh_op_bot_5')
// (15, 18, 'sp12_v_b_9')
// (15, 19, 'sp12_v_b_6')
// (15, 20, 'sp12_v_b_5')
// (15, 21, 'local_g2_2')
// (15, 21, 'lutff_5/in_3')
// (15, 21, 'sp12_v_b_2')
// (15, 22, 'sp12_v_b_1')
// (16, 16, 'neigh_op_tnl_5')
// (16, 17, 'neigh_op_lft_5')
// (16, 18, 'neigh_op_bnl_5')

wire n2135;
// (14, 15, 'neigh_op_tnr_3')
// (14, 16, 'neigh_op_rgt_3')
// (14, 17, 'neigh_op_bnr_3')
// (15, 15, 'local_g1_3')
// (15, 15, 'lutff_0/in_2')
// (15, 15, 'neigh_op_top_3')
// (15, 16, 'lutff_3/out')
// (15, 17, 'neigh_op_bot_3')
// (16, 15, 'neigh_op_tnl_3')
// (16, 16, 'neigh_op_lft_3')
// (16, 17, 'neigh_op_bnl_3')

wire n2136;
// (14, 15, 'neigh_op_tnr_5')
// (14, 16, 'neigh_op_rgt_5')
// (14, 17, 'neigh_op_bnr_5')
// (15, 15, 'local_g1_5')
// (15, 15, 'lutff_1/in_1')
// (15, 15, 'neigh_op_top_5')
// (15, 16, 'lutff_5/out')
// (15, 17, 'neigh_op_bot_5')
// (16, 15, 'neigh_op_tnl_5')
// (16, 16, 'neigh_op_lft_5')
// (16, 17, 'neigh_op_bnl_5')

wire n2137;
// (14, 15, 'sp4_h_r_3')
// (15, 15, 'sp4_h_r_14')
// (16, 12, 'sp4_r_v_b_43')
// (16, 13, 'sp4_r_v_b_30')
// (16, 14, 'neigh_op_tnr_3')
// (16, 14, 'sp4_r_v_b_19')
// (16, 15, 'neigh_op_rgt_3')
// (16, 15, 'sp4_h_r_27')
// (16, 15, 'sp4_r_v_b_6')
// (16, 16, 'neigh_op_bnr_3')
// (17, 11, 'sp4_h_r_6')
// (17, 11, 'sp4_v_t_43')
// (17, 12, 'local_g3_3')
// (17, 12, 'lutff_global/cen')
// (17, 12, 'sp4_r_v_b_42')
// (17, 12, 'sp4_r_v_b_46')
// (17, 12, 'sp4_v_b_43')
// (17, 13, 'sp4_r_v_b_31')
// (17, 13, 'sp4_r_v_b_35')
// (17, 13, 'sp4_r_v_b_47')
// (17, 13, 'sp4_v_b_30')
// (17, 14, 'neigh_op_top_3')
// (17, 14, 'sp4_r_v_b_18')
// (17, 14, 'sp4_r_v_b_22')
// (17, 14, 'sp4_r_v_b_34')
// (17, 14, 'sp4_v_b_19')
// (17, 15, 'lutff_3/out')
// (17, 15, 'sp4_h_r_38')
// (17, 15, 'sp4_h_r_6')
// (17, 15, 'sp4_r_v_b_11')
// (17, 15, 'sp4_r_v_b_23')
// (17, 15, 'sp4_r_v_b_7')
// (17, 15, 'sp4_v_b_6')
// (17, 16, 'neigh_op_bot_3')
// (17, 16, 'sp4_r_v_b_10')
// (18, 11, 'local_g1_3')
// (18, 11, 'lutff_global/cen')
// (18, 11, 'sp4_h_r_0')
// (18, 11, 'sp4_h_r_19')
// (18, 11, 'sp4_v_t_42')
// (18, 11, 'sp4_v_t_46')
// (18, 12, 'local_g2_2')
// (18, 12, 'lutff_global/cen')
// (18, 12, 'sp4_h_r_10')
// (18, 12, 'sp4_v_b_42')
// (18, 12, 'sp4_v_b_46')
// (18, 12, 'sp4_v_t_47')
// (18, 13, 'local_g3_3')
// (18, 13, 'lutff_global/cen')
// (18, 13, 'sp4_v_b_31')
// (18, 13, 'sp4_v_b_35')
// (18, 13, 'sp4_v_b_47')
// (18, 14, 'local_g3_3')
// (18, 14, 'lutff_global/cen')
// (18, 14, 'neigh_op_tnl_3')
// (18, 14, 'sp4_v_b_18')
// (18, 14, 'sp4_v_b_22')
// (18, 14, 'sp4_v_b_34')
// (18, 15, 'neigh_op_lft_3')
// (18, 15, 'sp4_h_l_38')
// (18, 15, 'sp4_h_r_11')
// (18, 15, 'sp4_h_r_19')
// (18, 15, 'sp4_v_b_11')
// (18, 15, 'sp4_v_b_23')
// (18, 15, 'sp4_v_b_7')
// (18, 16, 'neigh_op_bnl_3')
// (18, 16, 'sp4_v_b_10')
// (19, 11, 'sp4_h_r_13')
// (19, 11, 'sp4_h_r_30')
// (19, 12, 'sp4_h_r_23')
// (19, 15, 'sp4_h_r_22')
// (19, 15, 'sp4_h_r_30')
// (20, 11, 'local_g3_3')
// (20, 11, 'lutff_global/cen')
// (20, 11, 'sp4_h_r_24')
// (20, 11, 'sp4_h_r_43')
// (20, 12, 'sp4_h_r_34')
// (20, 12, 'sp4_r_v_b_43')
// (20, 13, 'sp4_r_v_b_30')
// (20, 14, 'local_g3_3')
// (20, 14, 'lutff_global/cen')
// (20, 14, 'sp4_r_v_b_19')
// (20, 15, 'sp4_h_r_35')
// (20, 15, 'sp4_h_r_43')
// (20, 15, 'sp4_r_v_b_6')
// (21, 8, 'sp4_r_v_b_43')
// (21, 9, 'sp4_r_v_b_30')
// (21, 10, 'local_g3_3')
// (21, 10, 'lutff_global/cen')
// (21, 10, 'sp4_r_v_b_19')
// (21, 11, 'sp4_h_l_43')
// (21, 11, 'sp4_h_r_37')
// (21, 11, 'sp4_r_v_b_6')
// (21, 11, 'sp4_v_t_43')
// (21, 12, 'sp4_h_r_47')
// (21, 12, 'sp4_v_b_43')
// (21, 13, 'sp4_v_b_30')
// (21, 14, 'sp4_v_b_19')
// (21, 15, 'sp4_h_l_43')
// (21, 15, 'sp4_h_r_46')
// (21, 15, 'sp4_v_b_6')
// (22, 7, 'sp4_v_t_43')
// (22, 8, 'sp4_v_b_43')
// (22, 9, 'sp4_v_b_30')
// (22, 10, 'sp4_v_b_19')
// (22, 11, 'sp4_h_l_37')
// (22, 11, 'sp4_v_b_6')
// (22, 12, 'local_g0_1')
// (22, 12, 'local_g0_2')
// (22, 12, 'lutff_1/in_2')
// (22, 12, 'lutff_global/cen')
// (22, 12, 'sp4_h_l_47')
// (22, 12, 'sp4_h_r_1')
// (22, 12, 'sp4_h_r_10')
// (22, 15, 'sp4_h_l_46')
// (23, 12, 'sp4_h_r_12')
// (23, 12, 'sp4_h_r_23')
// (24, 12, 'sp4_h_r_25')
// (24, 12, 'sp4_h_r_34')
// (25, 12, 'sp4_h_r_36')
// (25, 12, 'sp4_h_r_47')

wire n2138;
// (14, 15, 'sp4_h_r_8')
// (15, 15, 'sp4_h_r_21')
// (16, 14, 'neigh_op_tnr_1')
// (16, 15, 'neigh_op_rgt_1')
// (16, 15, 'sp4_h_r_32')
// (16, 16, 'neigh_op_bnr_1')
// (17, 12, 'sp4_r_v_b_38')
// (17, 13, 'sp4_r_v_b_27')
// (17, 14, 'neigh_op_top_1')
// (17, 14, 'sp4_r_v_b_14')
// (17, 15, 'local_g3_5')
// (17, 15, 'lutff_1/out')
// (17, 15, 'lutff_global/s_r')
// (17, 15, 'sp4_h_r_45')
// (17, 15, 'sp4_r_v_b_3')
// (17, 16, 'neigh_op_bot_1')
// (18, 11, 'sp4_v_t_38')
// (18, 12, 'sp4_v_b_38')
// (18, 13, 'sp4_v_b_27')
// (18, 14, 'neigh_op_tnl_1')
// (18, 14, 'sp4_v_b_14')
// (18, 15, 'neigh_op_lft_1')
// (18, 15, 'sp4_h_l_45')
// (18, 15, 'sp4_v_b_3')
// (18, 16, 'neigh_op_bnl_1')

wire n2139;
// (14, 17, 'neigh_op_tnr_2')
// (14, 18, 'local_g3_2')
// (14, 18, 'lutff_0/in_1')
// (14, 18, 'neigh_op_rgt_2')
// (14, 19, 'neigh_op_bnr_2')
// (15, 17, 'neigh_op_top_2')
// (15, 18, 'lutff_2/out')
// (15, 19, 'neigh_op_bot_2')
// (16, 17, 'neigh_op_tnl_2')
// (16, 18, 'neigh_op_lft_2')
// (16, 19, 'neigh_op_bnl_2')

wire n2140;
// (14, 17, 'neigh_op_tnr_4')
// (14, 18, 'local_g3_4')
// (14, 18, 'lutff_1/in_2')
// (14, 18, 'neigh_op_rgt_4')
// (14, 19, 'neigh_op_bnr_4')
// (15, 17, 'neigh_op_top_4')
// (15, 18, 'lutff_4/out')
// (15, 19, 'neigh_op_bot_4')
// (16, 17, 'neigh_op_tnl_4')
// (16, 18, 'neigh_op_lft_4')
// (16, 19, 'neigh_op_bnl_4')

wire n2141;
// (14, 17, 'neigh_op_tnr_6')
// (14, 18, 'local_g2_6')
// (14, 18, 'lutff_3/in_3')
// (14, 18, 'neigh_op_rgt_6')
// (14, 19, 'neigh_op_bnr_6')
// (15, 17, 'neigh_op_top_6')
// (15, 18, 'lutff_6/out')
// (15, 19, 'neigh_op_bot_6')
// (16, 17, 'neigh_op_tnl_6')
// (16, 18, 'neigh_op_lft_6')
// (16, 19, 'neigh_op_bnl_6')

reg n2142 = 0;
// (14, 18, 'local_g1_2')
// (14, 18, 'lutff_2/in_3')
// (14, 18, 'sp4_h_r_10')
// (15, 17, 'neigh_op_tnr_1')
// (15, 18, 'local_g2_1')
// (15, 18, 'lutff_1/in_2')
// (15, 18, 'neigh_op_rgt_1')
// (15, 18, 'sp4_h_r_23')
// (15, 19, 'neigh_op_bnr_1')
// (16, 17, 'neigh_op_top_1')
// (16, 18, 'local_g0_1')
// (16, 18, 'lutff_1/in_2')
// (16, 18, 'lutff_1/out')
// (16, 18, 'sp4_h_r_34')
// (16, 19, 'neigh_op_bot_1')
// (17, 17, 'neigh_op_tnl_1')
// (17, 18, 'neigh_op_lft_1')
// (17, 18, 'sp4_h_r_47')
// (17, 19, 'neigh_op_bnl_1')
// (18, 18, 'sp4_h_l_47')

wire n2143;
// (14, 18, 'local_g1_4')
// (14, 18, 'lutff_3/in_2')
// (14, 18, 'sp4_h_r_4')
// (15, 17, 'neigh_op_tnr_6')
// (15, 18, 'neigh_op_rgt_6')
// (15, 18, 'sp4_h_r_17')
// (15, 19, 'neigh_op_bnr_6')
// (16, 17, 'neigh_op_top_6')
// (16, 18, 'lutff_6/out')
// (16, 18, 'sp4_h_r_28')
// (16, 19, 'neigh_op_bot_6')
// (17, 17, 'neigh_op_tnl_6')
// (17, 18, 'neigh_op_lft_6')
// (17, 18, 'sp4_h_r_41')
// (17, 19, 'neigh_op_bnl_6')
// (18, 18, 'sp4_h_l_41')

wire n2144;
// (14, 18, 'neigh_op_tnr_0')
// (14, 19, 'neigh_op_rgt_0')
// (14, 20, 'neigh_op_bnr_0')
// (15, 18, 'neigh_op_top_0')
// (15, 19, 'lutff_0/out')
// (15, 20, 'neigh_op_bot_0')
// (16, 18, 'neigh_op_tnl_0')
// (16, 19, 'local_g0_0')
// (16, 19, 'lutff_7/in_1')
// (16, 19, 'neigh_op_lft_0')
// (16, 20, 'neigh_op_bnl_0')

wire n2145;
// (14, 18, 'neigh_op_tnr_2')
// (14, 19, 'neigh_op_rgt_2')
// (14, 20, 'neigh_op_bnr_2')
// (15, 18, 'neigh_op_top_2')
// (15, 19, 'lutff_2/out')
// (15, 20, 'neigh_op_bot_2')
// (16, 18, 'neigh_op_tnl_2')
// (16, 19, 'local_g0_2')
// (16, 19, 'lutff_6/in_2')
// (16, 19, 'neigh_op_lft_2')
// (16, 20, 'neigh_op_bnl_2')

wire n2146;
// (14, 18, 'neigh_op_tnr_4')
// (14, 19, 'neigh_op_rgt_4')
// (14, 20, 'neigh_op_bnr_4')
// (15, 18, 'neigh_op_top_4')
// (15, 19, 'lutff_4/out')
// (15, 20, 'neigh_op_bot_4')
// (16, 18, 'neigh_op_tnl_4')
// (16, 19, 'local_g0_4')
// (16, 19, 'lutff_4/in_0')
// (16, 19, 'neigh_op_lft_4')
// (16, 20, 'neigh_op_bnl_4')

wire n2147;
// (14, 19, 'lutff_0/cout')
// (14, 19, 'lutff_1/in_3')

wire n2148;
// (14, 19, 'lutff_1/cout')
// (14, 19, 'lutff_2/in_3')

wire n2149;
// (14, 19, 'lutff_2/cout')
// (14, 19, 'lutff_3/in_3')

wire n2150;
// (14, 19, 'lutff_3/cout')
// (14, 19, 'lutff_4/in_3')

wire n2151;
// (14, 19, 'lutff_4/cout')
// (14, 19, 'lutff_5/in_3')

wire n2152;
// (14, 19, 'neigh_op_tnr_0')
// (14, 20, 'neigh_op_rgt_0')
// (14, 21, 'neigh_op_bnr_0')
// (15, 19, 'neigh_op_top_0')
// (15, 20, 'local_g1_0')
// (15, 20, 'lutff_0/out')
// (15, 20, 'lutff_7/in_0')
// (15, 21, 'neigh_op_bot_0')
// (16, 19, 'neigh_op_tnl_0')
// (16, 20, 'neigh_op_lft_0')
// (16, 21, 'neigh_op_bnl_0')

wire n2153;
// (14, 19, 'neigh_op_tnr_3')
// (14, 20, 'neigh_op_rgt_3')
// (14, 21, 'neigh_op_bnr_3')
// (15, 19, 'neigh_op_top_3')
// (15, 20, 'local_g0_3')
// (15, 20, 'lutff_2/in_1')
// (15, 20, 'lutff_3/out')
// (15, 21, 'neigh_op_bot_3')
// (16, 19, 'neigh_op_tnl_3')
// (16, 20, 'neigh_op_lft_3')
// (16, 21, 'neigh_op_bnl_3')

wire n2154;
// (14, 19, 'neigh_op_tnr_5')
// (14, 20, 'neigh_op_rgt_5')
// (14, 21, 'neigh_op_bnr_5')
// (15, 19, 'neigh_op_top_5')
// (15, 20, 'local_g0_5')
// (15, 20, 'lutff_5/out')
// (15, 20, 'lutff_7/in_2')
// (15, 21, 'neigh_op_bot_5')
// (16, 19, 'neigh_op_tnl_5')
// (16, 20, 'local_g0_5')
// (16, 20, 'lutff_3/in_2')
// (16, 20, 'neigh_op_lft_5')
// (16, 21, 'neigh_op_bnl_5')

reg n2155 = 0;
// (14, 20, 'local_g3_5')
// (14, 20, 'lutff_global/s_r')
// (14, 20, 'neigh_op_tnr_5')
// (14, 21, 'local_g3_5')
// (14, 21, 'lutff_6/in_2')
// (14, 21, 'neigh_op_rgt_5')
// (14, 22, 'neigh_op_bnr_5')
// (15, 20, 'neigh_op_top_5')
// (15, 21, 'lutff_5/out')
// (15, 22, 'neigh_op_bot_5')
// (16, 20, 'local_g3_5')
// (16, 20, 'lutff_3/in_1')
// (16, 20, 'neigh_op_tnl_5')
// (16, 21, 'neigh_op_lft_5')
// (16, 22, 'neigh_op_bnl_5')

reg n2156 = 0;
// (14, 20, 'sp4_h_r_1')
// (15, 20, 'sp4_h_r_12')
// (15, 21, 'sp4_r_v_b_38')
// (15, 22, 'sp4_r_v_b_27')
// (15, 23, 'sp4_r_v_b_14')
// (15, 24, 'sp4_r_v_b_3')
// (16, 17, 'sp4_r_v_b_41')
// (16, 18, 'sp4_r_v_b_28')
// (16, 19, 'local_g2_2')
// (16, 19, 'lutff_5/in_3')
// (16, 19, 'neigh_op_tnr_2')
// (16, 19, 'sp4_r_v_b_17')
// (16, 20, 'local_g2_2')
// (16, 20, 'lutff_2/in_2')
// (16, 20, 'lutff_6/in_2')
// (16, 20, 'neigh_op_rgt_2')
// (16, 20, 'sp4_h_r_25')
// (16, 20, 'sp4_h_r_9')
// (16, 20, 'sp4_r_v_b_36')
// (16, 20, 'sp4_r_v_b_4')
// (16, 20, 'sp4_v_t_38')
// (16, 21, 'local_g0_2')
// (16, 21, 'lutff_7/in_1')
// (16, 21, 'neigh_op_bnr_2')
// (16, 21, 'sp4_r_v_b_25')
// (16, 21, 'sp4_v_b_38')
// (16, 22, 'local_g2_4')
// (16, 22, 'lutff_2/in_0')
// (16, 22, 'sp4_r_v_b_12')
// (16, 22, 'sp4_v_b_27')
// (16, 23, 'local_g1_1')
// (16, 23, 'lutff_0/in_0')
// (16, 23, 'lutff_7/in_3')
// (16, 23, 'sp4_r_v_b_1')
// (16, 23, 'sp4_v_b_14')
// (16, 24, 'local_g0_3')
// (16, 24, 'lutff_3/in_2')
// (16, 24, 'sp4_v_b_3')
// (17, 13, 'sp4_r_v_b_45')
// (17, 14, 'sp4_r_v_b_32')
// (17, 15, 'sp4_r_v_b_21')
// (17, 16, 'sp4_h_r_4')
// (17, 16, 'sp4_r_v_b_8')
// (17, 16, 'sp4_v_t_41')
// (17, 17, 'sp4_r_v_b_40')
// (17, 17, 'sp4_v_b_41')
// (17, 18, 'sp4_r_v_b_29')
// (17, 18, 'sp4_r_v_b_45')
// (17, 18, 'sp4_v_b_28')
// (17, 19, 'local_g0_2')
// (17, 19, 'lutff_5/in_1')
// (17, 19, 'neigh_op_top_2')
// (17, 19, 'sp4_r_v_b_16')
// (17, 19, 'sp4_r_v_b_32')
// (17, 19, 'sp4_v_b_17')
// (17, 19, 'sp4_v_t_36')
// (17, 20, 'local_g2_2')
// (17, 20, 'lutff_2/in_0')
// (17, 20, 'lutff_2/out')
// (17, 20, 'sp4_h_r_20')
// (17, 20, 'sp4_h_r_36')
// (17, 20, 'sp4_r_v_b_21')
// (17, 20, 'sp4_r_v_b_37')
// (17, 20, 'sp4_r_v_b_5')
// (17, 20, 'sp4_v_b_36')
// (17, 20, 'sp4_v_b_4')
// (17, 21, 'local_g1_2')
// (17, 21, 'lutff_1/in_0')
// (17, 21, 'lutff_4/in_1')
// (17, 21, 'neigh_op_bot_2')
// (17, 21, 'sp4_r_v_b_24')
// (17, 21, 'sp4_r_v_b_8')
// (17, 21, 'sp4_v_b_25')
// (17, 22, 'local_g0_4')
// (17, 22, 'lutff_6/in_2')
// (17, 22, 'sp4_r_v_b_13')
// (17, 22, 'sp4_r_v_b_46')
// (17, 22, 'sp4_v_b_12')
// (17, 23, 'local_g1_0')
// (17, 23, 'lutff_2/in_1')
// (17, 23, 'sp4_r_v_b_0')
// (17, 23, 'sp4_r_v_b_35')
// (17, 23, 'sp4_v_b_1')
// (17, 24, 'local_g3_6')
// (17, 24, 'lutff_7/in_0')
// (17, 24, 'sp4_r_v_b_22')
// (17, 25, 'sp4_r_v_b_11')
// (18, 12, 'sp4_v_t_45')
// (18, 13, 'sp4_v_b_45')
// (18, 14, 'sp4_v_b_32')
// (18, 15, 'local_g0_5')
// (18, 15, 'lutff_5/in_2')
// (18, 15, 'sp4_v_b_21')
// (18, 16, 'sp4_h_r_17')
// (18, 16, 'sp4_h_r_5')
// (18, 16, 'sp4_v_b_8')
// (18, 16, 'sp4_v_t_40')
// (18, 17, 'local_g2_0')
// (18, 17, 'lutff_3/in_3')
// (18, 17, 'sp4_h_r_1')
// (18, 17, 'sp4_v_b_40')
// (18, 17, 'sp4_v_t_45')
// (18, 18, 'local_g2_5')
// (18, 18, 'lutff_2/in_3')
// (18, 18, 'sp4_v_b_29')
// (18, 18, 'sp4_v_b_45')
// (18, 19, 'local_g3_2')
// (18, 19, 'lutff_2/in_1')
// (18, 19, 'lutff_7/in_2')
// (18, 19, 'neigh_op_tnl_2')
// (18, 19, 'sp4_h_r_5')
// (18, 19, 'sp4_v_b_16')
// (18, 19, 'sp4_v_b_32')
// (18, 19, 'sp4_v_t_37')
// (18, 20, 'local_g0_2')
// (18, 20, 'lutff_7/in_1')
// (18, 20, 'neigh_op_lft_2')
// (18, 20, 'sp4_h_l_36')
// (18, 20, 'sp4_h_r_33')
// (18, 20, 'sp4_h_r_4')
// (18, 20, 'sp4_h_r_5')
// (18, 20, 'sp4_v_b_21')
// (18, 20, 'sp4_v_b_37')
// (18, 20, 'sp4_v_b_5')
// (18, 21, 'local_g3_2')
// (18, 21, 'lutff_2/in_1')
// (18, 21, 'neigh_op_bnl_2')
// (18, 21, 'sp4_h_r_2')
// (18, 21, 'sp4_v_b_24')
// (18, 21, 'sp4_v_b_8')
// (18, 21, 'sp4_v_t_46')
// (18, 22, 'local_g1_5')
// (18, 22, 'lutff_4/in_2')
// (18, 22, 'sp4_v_b_13')
// (18, 22, 'sp4_v_b_46')
// (18, 23, 'sp4_h_r_6')
// (18, 23, 'sp4_v_b_0')
// (18, 23, 'sp4_v_b_35')
// (18, 24, 'local_g1_6')
// (18, 24, 'lutff_4/in_3')
// (18, 24, 'sp4_v_b_22')
// (18, 25, 'sp4_v_b_11')
// (19, 16, 'sp4_h_r_16')
// (19, 16, 'sp4_h_r_28')
// (19, 17, 'sp4_h_r_12')
// (19, 17, 'sp4_r_v_b_44')
// (19, 18, 'sp4_r_v_b_33')
// (19, 19, 'sp4_h_r_16')
// (19, 19, 'sp4_r_v_b_20')
// (19, 20, 'sp4_h_r_16')
// (19, 20, 'sp4_h_r_17')
// (19, 20, 'sp4_h_r_44')
// (19, 20, 'sp4_r_v_b_9')
// (19, 21, 'sp4_h_r_15')
// (19, 21, 'sp4_r_v_b_44')
// (19, 22, 'sp4_r_v_b_33')
// (19, 23, 'sp4_h_r_19')
// (19, 23, 'sp4_r_v_b_20')
// (19, 24, 'sp4_r_v_b_9')
// (20, 13, 'sp4_r_v_b_41')
// (20, 14, 'sp4_r_v_b_28')
// (20, 15, 'local_g3_1')
// (20, 15, 'lutff_5/in_3')
// (20, 15, 'sp4_r_v_b_17')
// (20, 16, 'sp4_h_r_29')
// (20, 16, 'sp4_h_r_41')
// (20, 16, 'sp4_r_v_b_4')
// (20, 16, 'sp4_v_t_44')
// (20, 17, 'local_g3_1')
// (20, 17, 'lutff_7/in_1')
// (20, 17, 'sp4_h_r_25')
// (20, 17, 'sp4_v_b_44')
// (20, 18, 'local_g3_1')
// (20, 18, 'lutff_5/in_3')
// (20, 18, 'sp4_v_b_33')
// (20, 19, 'sp4_h_r_29')
// (20, 19, 'sp4_v_b_20')
// (20, 20, 'local_g0_0')
// (20, 20, 'lutff_0/in_0')
// (20, 20, 'lutff_4/in_2')
// (20, 20, 'lutff_6/in_0')
// (20, 20, 'sp4_h_l_44')
// (20, 20, 'sp4_h_r_0')
// (20, 20, 'sp4_h_r_28')
// (20, 20, 'sp4_h_r_29')
// (20, 20, 'sp4_v_b_9')
// (20, 20, 'sp4_v_t_44')
// (20, 21, 'local_g3_2')
// (20, 21, 'lutff_6/in_3')
// (20, 21, 'sp4_h_r_26')
// (20, 21, 'sp4_v_b_44')
// (20, 22, 'local_g2_1')
// (20, 22, 'lutff_4/in_3')
// (20, 22, 'sp4_v_b_33')
// (20, 23, 'local_g0_4')
// (20, 23, 'lutff_3/in_1')
// (20, 23, 'sp4_h_r_30')
// (20, 23, 'sp4_v_b_20')
// (20, 24, 'sp4_v_b_9')
// (21, 12, 'sp4_v_t_41')
// (21, 13, 'sp4_v_b_41')
// (21, 14, 'sp4_v_b_28')
// (21, 15, 'sp4_v_b_17')
// (21, 16, 'local_g3_0')
// (21, 16, 'lutff_5/in_2')
// (21, 16, 'sp4_h_l_41')
// (21, 16, 'sp4_h_r_40')
// (21, 16, 'sp4_r_v_b_46')
// (21, 16, 'sp4_v_b_4')
// (21, 17, 'local_g3_4')
// (21, 17, 'lutff_1/in_2')
// (21, 17, 'lutff_6/in_3')
// (21, 17, 'sp4_h_r_36')
// (21, 17, 'sp4_r_v_b_35')
// (21, 17, 'sp4_r_v_b_41')
// (21, 18, 'local_g3_6')
// (21, 18, 'lutff_6/in_3')
// (21, 18, 'sp4_r_v_b_22')
// (21, 18, 'sp4_r_v_b_28')
// (21, 19, 'local_g3_0')
// (21, 19, 'lutff_7/in_0')
// (21, 19, 'sp4_h_r_40')
// (21, 19, 'sp4_r_v_b_11')
// (21, 19, 'sp4_r_v_b_17')
// (21, 20, 'local_g2_0')
// (21, 20, 'lutff_5/in_3')
// (21, 20, 'sp4_h_r_13')
// (21, 20, 'sp4_h_r_40')
// (21, 20, 'sp4_h_r_41')
// (21, 20, 'sp4_r_v_b_37')
// (21, 20, 'sp4_r_v_b_4')
// (21, 21, 'local_g3_7')
// (21, 21, 'lutff_3/in_3')
// (21, 21, 'sp4_h_r_39')
// (21, 21, 'sp4_r_v_b_24')
// (21, 21, 'sp4_r_v_b_44')
// (21, 22, 'local_g2_5')
// (21, 22, 'lutff_5/in_0')
// (21, 22, 'sp4_r_v_b_13')
// (21, 22, 'sp4_r_v_b_33')
// (21, 23, 'local_g2_3')
// (21, 23, 'local_g3_3')
// (21, 23, 'lutff_4/in_2')
// (21, 23, 'lutff_7/in_2')
// (21, 23, 'sp4_h_r_43')
// (21, 23, 'sp4_r_v_b_0')
// (21, 23, 'sp4_r_v_b_20')
// (21, 24, 'sp4_r_v_b_9')
// (22, 15, 'sp4_v_t_46')
// (22, 16, 'local_g1_5')
// (22, 16, 'lutff_4/in_2')
// (22, 16, 'lutff_5/in_3')
// (22, 16, 'lutff_6/in_2')
// (22, 16, 'lutff_7/in_3')
// (22, 16, 'sp4_h_l_40')
// (22, 16, 'sp4_h_r_5')
// (22, 16, 'sp4_v_b_46')
// (22, 16, 'sp4_v_t_41')
// (22, 17, 'local_g1_1')
// (22, 17, 'lutff_1/in_3')
// (22, 17, 'lutff_3/in_1')
// (22, 17, 'lutff_4/in_2')
// (22, 17, 'lutff_6/in_2')
// (22, 17, 'sp4_h_l_36')
// (22, 17, 'sp4_h_r_1')
// (22, 17, 'sp4_v_b_35')
// (22, 17, 'sp4_v_b_41')
// (22, 18, 'local_g0_6')
// (22, 18, 'local_g3_4')
// (22, 18, 'lutff_0/in_1')
// (22, 18, 'lutff_1/in_2')
// (22, 18, 'lutff_3/in_3')
// (22, 18, 'sp4_v_b_22')
// (22, 18, 'sp4_v_b_28')
// (22, 19, 'local_g0_0')
// (22, 19, 'local_g1_1')
// (22, 19, 'lutff_0/in_0')
// (22, 19, 'lutff_4/in_0')
// (22, 19, 'lutff_6/in_2')
// (22, 19, 'sp4_h_l_40')
// (22, 19, 'sp4_h_r_8')
// (22, 19, 'sp4_v_b_11')
// (22, 19, 'sp4_v_b_17')
// (22, 19, 'sp4_v_t_37')
// (22, 20, 'local_g2_0')
// (22, 20, 'local_g3_0')
// (22, 20, 'lutff_2/in_3')
// (22, 20, 'lutff_3/in_2')
// (22, 20, 'lutff_4/in_2')
// (22, 20, 'lutff_6/in_1')
// (22, 20, 'lutff_7/in_3')
// (22, 20, 'sp4_h_l_40')
// (22, 20, 'sp4_h_l_41')
// (22, 20, 'sp4_h_r_24')
// (22, 20, 'sp4_v_b_37')
// (22, 20, 'sp4_v_b_4')
// (22, 20, 'sp4_v_t_44')
// (22, 21, 'local_g1_5')
// (22, 21, 'lutff_7/in_1')
// (22, 21, 'sp4_h_l_39')
// (22, 21, 'sp4_h_r_5')
// (22, 21, 'sp4_v_b_24')
// (22, 21, 'sp4_v_b_44')
// (22, 22, 'local_g2_1')
// (22, 22, 'lutff_3/in_0')
// (22, 22, 'lutff_7/in_2')
// (22, 22, 'sp4_v_b_13')
// (22, 22, 'sp4_v_b_33')
// (22, 23, 'local_g0_1')
// (22, 23, 'lutff_1/in_0')
// (22, 23, 'sp4_h_l_43')
// (22, 23, 'sp4_h_r_9')
// (22, 23, 'sp4_v_b_0')
// (22, 23, 'sp4_v_b_20')
// (22, 24, 'sp4_v_b_9')
// (23, 16, 'sp4_h_r_16')
// (23, 17, 'sp4_h_r_12')
// (23, 19, 'sp4_h_r_21')
// (23, 20, 'sp4_h_r_37')
// (23, 21, 'sp4_h_r_16')
// (23, 23, 'sp4_h_r_20')
// (24, 16, 'sp4_h_r_29')
// (24, 17, 'sp4_h_r_25')
// (24, 19, 'sp4_h_r_32')
// (24, 20, 'sp4_h_l_37')
// (24, 21, 'sp4_h_r_29')
// (24, 23, 'sp4_h_r_33')
// (25, 16, 'sp4_h_r_40')
// (25, 17, 'sp4_h_r_36')
// (25, 19, 'sp4_h_r_45')
// (25, 21, 'sp4_h_r_40')
// (25, 23, 'sp4_h_r_44')

wire n2157;
// (14, 20, 'sp4_r_v_b_47')
// (14, 21, 'sp4_r_v_b_34')
// (14, 22, 'sp4_r_v_b_23')
// (14, 23, 'sp4_r_v_b_10')
// (15, 19, 'sp4_v_t_47')
// (15, 20, 'sp4_v_b_47')
// (15, 21, 'sp4_v_b_34')
// (15, 22, 'neigh_op_tnr_0')
// (15, 22, 'sp4_v_b_23')
// (15, 23, 'local_g0_2')
// (15, 23, 'lutff_global/cen')
// (15, 23, 'neigh_op_rgt_0')
// (15, 23, 'sp4_h_r_5')
// (15, 23, 'sp4_v_b_10')
// (15, 24, 'neigh_op_bnr_0')
// (16, 22, 'neigh_op_top_0')
// (16, 23, 'lutff_0/out')
// (16, 23, 'sp4_h_r_16')
// (16, 24, 'neigh_op_bot_0')
// (17, 22, 'neigh_op_tnl_0')
// (17, 23, 'neigh_op_lft_0')
// (17, 23, 'sp4_h_r_29')
// (17, 24, 'neigh_op_bnl_0')
// (18, 23, 'sp4_h_r_40')
// (19, 23, 'sp4_h_l_40')

reg n2158 = 0;
// (14, 21, 'neigh_op_tnr_4')
// (14, 22, 'neigh_op_rgt_4')
// (14, 23, 'neigh_op_bnr_4')
// (15, 21, 'neigh_op_top_4')
// (15, 22, 'lutff_4/out')
// (15, 22, 'sp4_h_r_8')
// (15, 23, 'neigh_op_bot_4')
// (16, 21, 'neigh_op_tnl_4')
// (16, 22, 'neigh_op_lft_4')
// (16, 22, 'sp4_h_r_21')
// (16, 23, 'neigh_op_bnl_4')
// (17, 22, 'sp4_h_r_32')
// (18, 22, 'local_g3_5')
// (18, 22, 'lutff_2/in_0')
// (18, 22, 'sp4_h_r_45')
// (19, 22, 'sp4_h_l_45')

reg n2159 = 0;
// (14, 22, 'neigh_op_tnr_1')
// (14, 23, 'neigh_op_rgt_1')
// (14, 24, 'neigh_op_bnr_1')
// (15, 22, 'neigh_op_top_1')
// (15, 22, 'sp4_r_v_b_46')
// (15, 23, 'lutff_1/out')
// (15, 23, 'sp4_r_v_b_35')
// (15, 24, 'neigh_op_bot_1')
// (15, 24, 'sp4_r_v_b_22')
// (15, 25, 'sp4_r_v_b_11')
// (16, 21, 'sp4_h_r_4')
// (16, 21, 'sp4_v_t_46')
// (16, 22, 'neigh_op_tnl_1')
// (16, 22, 'sp4_v_b_46')
// (16, 23, 'neigh_op_lft_1')
// (16, 23, 'sp4_v_b_35')
// (16, 24, 'neigh_op_bnl_1')
// (16, 24, 'sp4_v_b_22')
// (16, 25, 'sp4_v_b_11')
// (17, 21, 'sp4_h_r_17')
// (18, 21, 'local_g2_4')
// (18, 21, 'lutff_1/in_1')
// (18, 21, 'sp4_h_r_28')
// (19, 21, 'sp4_h_r_41')
// (20, 21, 'sp4_h_l_41')

wire n2160;
// (14, 22, 'sp4_h_r_9')
// (15, 22, 'sp4_h_r_20')
// (16, 21, 'neigh_op_tnr_6')
// (16, 22, 'neigh_op_rgt_6')
// (16, 22, 'sp4_h_r_33')
// (16, 23, 'neigh_op_bnr_6')
// (17, 19, 'sp4_r_v_b_38')
// (17, 20, 'sp4_r_v_b_27')
// (17, 21, 'neigh_op_top_6')
// (17, 21, 'sp4_r_v_b_14')
// (17, 22, 'local_g1_3')
// (17, 22, 'lutff_6/out')
// (17, 22, 'lutff_global/cen')
// (17, 22, 'sp4_h_r_44')
// (17, 22, 'sp4_r_v_b_3')
// (17, 23, 'neigh_op_bot_6')
// (18, 18, 'sp4_v_t_38')
// (18, 19, 'sp4_v_b_38')
// (18, 20, 'sp4_v_b_27')
// (18, 21, 'neigh_op_tnl_6')
// (18, 21, 'sp4_v_b_14')
// (18, 22, 'neigh_op_lft_6')
// (18, 22, 'sp4_h_l_44')
// (18, 22, 'sp4_v_b_3')
// (18, 23, 'neigh_op_bnl_6')

wire n2161;
// (14, 23, 'lutff_0/cout')
// (14, 23, 'lutff_1/in_3')

wire n2162;
// (14, 23, 'lutff_1/cout')
// (14, 23, 'lutff_2/in_3')

wire n2163;
// (14, 23, 'lutff_2/cout')
// (14, 23, 'lutff_3/in_3')

wire n2164;
// (14, 23, 'lutff_3/cout')
// (14, 23, 'lutff_4/in_3')

wire n2165;
// (14, 23, 'lutff_4/cout')
// (14, 23, 'lutff_5/in_3')

wire n2166;
// (14, 23, 'lutff_5/cout')
// (14, 23, 'lutff_6/in_3')

reg n2167 = 0;
// (15, 0, 'logic_op_tnr_5')
// (15, 1, 'neigh_op_rgt_5')
// (15, 2, 'neigh_op_bnr_5')
// (16, 0, 'logic_op_top_5')
// (16, 1, 'local_g2_5')
// (16, 1, 'lutff_1/in_2')
// (16, 1, 'lutff_5/out')
// (16, 2, 'neigh_op_bot_5')
// (17, 0, 'logic_op_tnl_5')
// (17, 1, 'neigh_op_lft_5')
// (17, 2, 'neigh_op_bnl_5')

wire io_16_0_0;
// (15, 1, 'neigh_op_bnr_0')
// (15, 1, 'neigh_op_bnr_4')
// (16, 0, 'io_0/D_IN_0')
// (16, 0, 'io_0/PAD')
// (16, 1, 'local_g0_4')
// (16, 1, 'lutff_5/in_1')
// (16, 1, 'neigh_op_bot_0')
// (16, 1, 'neigh_op_bot_4')
// (17, 1, 'neigh_op_bnl_0')
// (17, 1, 'neigh_op_bnl_4')

reg n2169 = 0;
// (15, 1, 'neigh_op_tnr_7')
// (15, 2, 'local_g2_7')
// (15, 2, 'lutff_7/in_0')
// (15, 2, 'neigh_op_rgt_7')
// (15, 2, 'sp4_r_v_b_46')
// (15, 3, 'neigh_op_bnr_7')
// (15, 3, 'sp4_r_v_b_35')
// (15, 4, 'sp4_r_v_b_22')
// (15, 5, 'sp4_r_v_b_11')
// (15, 6, 'sp4_r_v_b_42')
// (15, 7, 'sp4_r_v_b_31')
// (15, 8, 'local_g3_2')
// (15, 8, 'lutff_2/in_1')
// (15, 8, 'lutff_6/in_3')
// (15, 8, 'sp4_r_v_b_18')
// (15, 9, 'sp4_r_v_b_7')
// (16, 0, 'span12_vert_17')
// (16, 1, 'neigh_op_top_7')
// (16, 1, 'sp12_v_b_17')
// (16, 1, 'sp4_v_t_46')
// (16, 2, 'lutff_7/out')
// (16, 2, 'sp12_v_b_14')
// (16, 2, 'sp4_v_b_46')
// (16, 3, 'neigh_op_bot_7')
// (16, 3, 'sp12_v_b_13')
// (16, 3, 'sp4_v_b_35')
// (16, 4, 'sp12_v_b_10')
// (16, 4, 'sp4_v_b_22')
// (16, 5, 'sp12_v_b_9')
// (16, 5, 'sp4_v_b_11')
// (16, 5, 'sp4_v_t_42')
// (16, 6, 'sp12_v_b_6')
// (16, 6, 'sp4_v_b_42')
// (16, 7, 'sp12_v_b_5')
// (16, 7, 'sp4_v_b_31')
// (16, 8, 'local_g2_2')
// (16, 8, 'lutff_3/in_3')
// (16, 8, 'sp12_v_b_2')
// (16, 8, 'sp4_v_b_18')
// (16, 9, 'sp12_v_b_1')
// (16, 9, 'sp4_v_b_7')
// (17, 1, 'neigh_op_tnl_7')
// (17, 2, 'neigh_op_lft_7')
// (17, 3, 'neigh_op_bnl_7')

wire n2170;
// (15, 2, 'sp4_h_r_8')
// (16, 1, 'neigh_op_tnr_0')
// (16, 1, 'sp4_r_v_b_45')
// (16, 2, 'neigh_op_rgt_0')
// (16, 2, 'sp4_h_r_21')
// (16, 2, 'sp4_r_v_b_32')
// (16, 3, 'neigh_op_bnr_0')
// (16, 3, 'sp4_r_v_b_21')
// (16, 4, 'sp4_r_v_b_8')
// (17, 0, 'span4_vert_45')
// (17, 1, 'neigh_op_top_0')
// (17, 1, 'sp4_v_b_45')
// (17, 2, 'local_g2_0')
// (17, 2, 'lutff_0/out')
// (17, 2, 'lutff_2/in_2')
// (17, 2, 'sp4_h_r_32')
// (17, 2, 'sp4_v_b_32')
// (17, 3, 'neigh_op_bot_0')
// (17, 3, 'sp4_v_b_21')
// (17, 4, 'local_g0_0')
// (17, 4, 'lutff_1/in_1')
// (17, 4, 'sp4_v_b_8')
// (18, 1, 'neigh_op_tnl_0')
// (18, 2, 'neigh_op_lft_0')
// (18, 2, 'sp4_h_r_45')
// (18, 3, 'neigh_op_bnl_0')
// (19, 2, 'sp4_h_l_45')
// (19, 2, 'sp4_h_r_4')
// (20, 2, 'sp4_h_r_17')
// (21, 2, 'sp4_h_r_28')
// (22, 2, 'sp4_h_r_41')
// (22, 3, 'sp4_r_v_b_41')
// (22, 4, 'sp4_r_v_b_28')
// (22, 5, 'local_g3_1')
// (22, 5, 'lutff_5/in_3')
// (22, 5, 'sp4_r_v_b_17')
// (22, 6, 'sp4_r_v_b_4')
// (23, 2, 'sp4_h_l_41')
// (23, 2, 'sp4_v_t_41')
// (23, 3, 'sp4_v_b_41')
// (23, 4, 'sp4_v_b_28')
// (23, 5, 'sp4_v_b_17')
// (23, 6, 'sp4_v_b_4')

reg n2171 = 0;
// (15, 2, 'sp4_h_r_9')
// (16, 2, 'sp4_h_r_20')
// (17, 1, 'neigh_op_tnr_6')
// (17, 2, 'neigh_op_rgt_6')
// (17, 2, 'sp4_h_r_33')
// (17, 3, 'neigh_op_bnr_6')
// (18, 1, 'neigh_op_top_6')
// (18, 2, 'lutff_6/out')
// (18, 2, 'sp4_h_r_44')
// (18, 3, 'neigh_op_bot_6')
// (18, 3, 'sp4_r_v_b_39')
// (18, 4, 'sp4_r_v_b_26')
// (18, 5, 'sp4_r_v_b_15')
// (18, 6, 'sp4_r_v_b_2')
// (19, 1, 'neigh_op_tnl_6')
// (19, 2, 'neigh_op_lft_6')
// (19, 2, 'sp4_h_l_44')
// (19, 2, 'sp4_v_t_39')
// (19, 3, 'neigh_op_bnl_6')
// (19, 3, 'sp4_v_b_39')
// (19, 4, 'sp4_v_b_26')
// (19, 5, 'sp4_v_b_15')
// (19, 6, 'local_g0_2')
// (19, 6, 'ram/WDATA_0')
// (19, 6, 'sp4_v_b_2')

wire n2172;
// (15, 3, 'neigh_op_tnr_0')
// (15, 4, 'neigh_op_rgt_0')
// (15, 5, 'neigh_op_bnr_0')
// (16, 3, 'neigh_op_top_0')
// (16, 4, 'local_g3_0')
// (16, 4, 'lutff_0/out')
// (16, 4, 'lutff_5/in_0')
// (16, 5, 'neigh_op_bot_0')
// (17, 3, 'neigh_op_tnl_0')
// (17, 4, 'local_g1_0')
// (17, 4, 'lutff_3/in_0')
// (17, 4, 'neigh_op_lft_0')
// (17, 5, 'local_g3_0')
// (17, 5, 'lutff_6/in_3')
// (17, 5, 'neigh_op_bnl_0')

wire n2173;
// (15, 3, 'neigh_op_tnr_1')
// (15, 4, 'neigh_op_rgt_1')
// (15, 5, 'neigh_op_bnr_1')
// (16, 2, 'sp4_r_v_b_43')
// (16, 3, 'neigh_op_top_1')
// (16, 3, 'sp4_r_v_b_30')
// (16, 4, 'local_g0_1')
// (16, 4, 'lutff_1/out')
// (16, 4, 'lutff_3/in_2')
// (16, 4, 'sp4_h_r_2')
// (16, 4, 'sp4_r_v_b_19')
// (16, 5, 'neigh_op_bot_1')
// (16, 5, 'sp4_r_v_b_6')
// (17, 1, 'sp4_v_t_43')
// (17, 2, 'sp4_v_b_43')
// (17, 3, 'neigh_op_tnl_1')
// (17, 3, 'sp4_v_b_30')
// (17, 4, 'local_g1_1')
// (17, 4, 'lutff_0/in_2')
// (17, 4, 'neigh_op_lft_1')
// (17, 4, 'sp4_h_r_15')
// (17, 4, 'sp4_v_b_19')
// (17, 5, 'neigh_op_bnl_1')
// (17, 5, 'sp4_h_r_0')
// (17, 5, 'sp4_v_b_6')
// (18, 4, 'local_g2_2')
// (18, 4, 'lutff_0/in_0')
// (18, 4, 'sp4_h_r_26')
// (18, 5, 'local_g1_5')
// (18, 5, 'lutff_7/in_1')
// (18, 5, 'sp4_h_r_13')
// (19, 4, 'sp4_h_r_39')
// (19, 5, 'sp4_h_r_24')
// (20, 4, 'sp4_h_l_39')
// (20, 5, 'sp4_h_r_37')
// (21, 5, 'sp4_h_l_37')

reg n2174 = 0;
// (15, 3, 'neigh_op_tnr_2')
// (15, 4, 'neigh_op_rgt_2')
// (15, 5, 'neigh_op_bnr_2')
// (16, 3, 'neigh_op_top_2')
// (16, 4, 'local_g3_2')
// (16, 4, 'lutff_0/in_3')
// (16, 4, 'lutff_2/out')
// (16, 5, 'neigh_op_bot_2')
// (17, 3, 'neigh_op_tnl_2')
// (17, 4, 'neigh_op_lft_2')
// (17, 5, 'neigh_op_bnl_2')

reg n2175 = 0;
// (15, 3, 'neigh_op_tnr_3')
// (15, 4, 'neigh_op_rgt_3')
// (15, 5, 'neigh_op_bnr_3')
// (16, 3, 'neigh_op_top_3')
// (16, 4, 'local_g0_3')
// (16, 4, 'lutff_1/in_2')
// (16, 4, 'lutff_3/out')
// (16, 5, 'neigh_op_bot_3')
// (17, 3, 'neigh_op_tnl_3')
// (17, 4, 'neigh_op_lft_3')
// (17, 5, 'neigh_op_bnl_3')

reg n2176 = 0;
// (15, 3, 'neigh_op_tnr_5')
// (15, 4, 'neigh_op_rgt_5')
// (15, 5, 'neigh_op_bnr_5')
// (16, 3, 'neigh_op_top_5')
// (16, 4, 'local_g2_5')
// (16, 4, 'lutff_0/in_1')
// (16, 4, 'lutff_5/out')
// (16, 5, 'neigh_op_bot_5')
// (17, 3, 'neigh_op_tnl_5')
// (17, 4, 'neigh_op_lft_5')
// (17, 5, 'neigh_op_bnl_5')

reg n2177 = 0;
// (15, 3, 'neigh_op_tnr_7')
// (15, 4, 'neigh_op_rgt_7')
// (15, 5, 'neigh_op_bnr_7')
// (16, 3, 'neigh_op_top_7')
// (16, 4, 'local_g3_7')
// (16, 4, 'lutff_1/in_3')
// (16, 4, 'lutff_7/out')
// (16, 5, 'neigh_op_bot_7')
// (17, 3, 'neigh_op_tnl_7')
// (17, 4, 'neigh_op_lft_7')
// (17, 5, 'neigh_op_bnl_7')

reg n2178 = 0;
// (15, 3, 'sp4_h_r_11')
// (15, 5, 'sp4_h_r_7')
// (16, 3, 'local_g1_6')
// (16, 3, 'lutff_3/in_2')
// (16, 3, 'sp4_h_r_22')
// (16, 4, 'sp4_r_v_b_44')
// (16, 5, 'local_g1_2')
// (16, 5, 'lutff_4/in_3')
// (16, 5, 'sp4_h_r_18')
// (16, 5, 'sp4_r_v_b_33')
// (16, 6, 'sp4_r_v_b_20')
// (16, 7, 'sp4_r_v_b_9')
// (17, 2, 'neigh_op_tnr_7')
// (17, 3, 'neigh_op_rgt_7')
// (17, 3, 'sp4_h_r_3')
// (17, 3, 'sp4_h_r_35')
// (17, 3, 'sp4_v_t_44')
// (17, 4, 'neigh_op_bnr_7')
// (17, 4, 'sp4_v_b_44')
// (17, 5, 'sp4_h_r_31')
// (17, 5, 'sp4_v_b_33')
// (17, 6, 'sp4_v_b_20')
// (17, 7, 'local_g1_1')
// (17, 7, 'lutff_4/in_2')
// (17, 7, 'sp4_v_b_9')
// (18, 2, 'neigh_op_top_7')
// (18, 2, 'sp4_r_v_b_42')
// (18, 3, 'local_g0_7')
// (18, 3, 'lutff_7/in_0')
// (18, 3, 'lutff_7/out')
// (18, 3, 'sp4_h_r_14')
// (18, 3, 'sp4_h_r_46')
// (18, 3, 'sp4_r_v_b_31')
// (18, 4, 'neigh_op_bot_7')
// (18, 4, 'sp4_r_v_b_18')
// (18, 5, 'sp4_h_r_42')
// (18, 5, 'sp4_r_v_b_7')
// (19, 1, 'sp4_v_t_42')
// (19, 2, 'neigh_op_tnl_7')
// (19, 2, 'sp4_v_b_42')
// (19, 3, 'neigh_op_lft_7')
// (19, 3, 'sp4_h_l_46')
// (19, 3, 'sp4_h_r_27')
// (19, 3, 'sp4_v_b_31')
// (19, 4, 'neigh_op_bnl_7')
// (19, 4, 'sp4_v_b_18')
// (19, 5, 'sp4_h_l_42')
// (19, 5, 'sp4_v_b_7')
// (20, 3, 'sp4_h_r_38')
// (21, 3, 'sp4_h_l_38')

reg n2179 = 0;
// (15, 4, 'local_g2_2')
// (15, 4, 'lutff_6/in_0')
// (15, 4, 'neigh_op_tnr_2')
// (15, 5, 'neigh_op_rgt_2')
// (15, 5, 'sp4_r_v_b_36')
// (15, 6, 'neigh_op_bnr_2')
// (15, 6, 'sp4_r_v_b_25')
// (15, 7, 'sp4_r_v_b_12')
// (15, 8, 'local_g1_1')
// (15, 8, 'lutff_2/in_2')
// (15, 8, 'lutff_6/in_2')
// (15, 8, 'sp4_r_v_b_1')
// (16, 4, 'neigh_op_top_2')
// (16, 4, 'sp4_v_t_36')
// (16, 5, 'lutff_2/out')
// (16, 5, 'sp4_v_b_36')
// (16, 6, 'neigh_op_bot_2')
// (16, 6, 'sp4_v_b_25')
// (16, 7, 'sp4_v_b_12')
// (16, 8, 'local_g0_1')
// (16, 8, 'lutff_3/in_2')
// (16, 8, 'sp4_v_b_1')
// (17, 4, 'neigh_op_tnl_2')
// (17, 5, 'neigh_op_lft_2')
// (17, 6, 'neigh_op_bnl_2')

wire n2180;
// (15, 4, 'neigh_op_tnr_6')
// (15, 5, 'neigh_op_rgt_6')
// (15, 6, 'neigh_op_bnr_6')
// (16, 4, 'neigh_op_top_6')
// (16, 5, 'local_g2_6')
// (16, 5, 'lutff_1/in_3')
// (16, 5, 'lutff_6/out')
// (16, 6, 'neigh_op_bot_6')
// (17, 4, 'neigh_op_tnl_6')
// (17, 5, 'neigh_op_lft_6')
// (17, 6, 'neigh_op_bnl_6')

wire n2181;
// (15, 4, 'neigh_op_tnr_7')
// (15, 5, 'neigh_op_rgt_7')
// (15, 6, 'neigh_op_bnr_7')
// (16, 4, 'neigh_op_top_7')
// (16, 5, 'local_g1_7')
// (16, 5, 'lutff_1/in_1')
// (16, 5, 'lutff_7/out')
// (16, 6, 'neigh_op_bot_7')
// (17, 4, 'neigh_op_tnl_7')
// (17, 5, 'neigh_op_lft_7')
// (17, 6, 'neigh_op_bnl_7')

wire n2182;
// (15, 4, 'sp4_h_r_7')
// (16, 4, 'local_g1_2')
// (16, 4, 'lutff_3/in_0')
// (16, 4, 'lutff_7/in_0')
// (16, 4, 'sp4_h_r_18')
// (17, 1, 'neigh_op_tnr_7')
// (17, 2, 'local_g3_7')
// (17, 2, 'lutff_1/in_3')
// (17, 2, 'lutff_3/in_3')
// (17, 2, 'lutff_4/in_2')
// (17, 2, 'lutff_7/in_3')
// (17, 2, 'neigh_op_rgt_7')
// (17, 3, 'local_g1_7')
// (17, 3, 'lutff_0/in_0')
// (17, 3, 'lutff_6/in_0')
// (17, 3, 'neigh_op_bnr_7')
// (17, 4, 'sp4_h_r_31')
// (18, 1, 'neigh_op_top_7')
// (18, 1, 'sp4_r_v_b_42')
// (18, 2, 'lutff_7/out')
// (18, 2, 'sp4_r_v_b_31')
// (18, 3, 'neigh_op_bot_7')
// (18, 3, 'sp4_r_v_b_18')
// (18, 4, 'sp4_h_r_42')
// (18, 4, 'sp4_r_v_b_7')
// (19, 0, 'span4_vert_42')
// (19, 1, 'neigh_op_tnl_7')
// (19, 1, 'sp4_v_b_42')
// (19, 2, 'neigh_op_lft_7')
// (19, 2, 'sp4_v_b_31')
// (19, 3, 'neigh_op_bnl_7')
// (19, 3, 'sp4_v_b_18')
// (19, 4, 'sp4_h_l_42')
// (19, 4, 'sp4_v_b_7')

wire io_19_0_1;
// (15, 4, 'sp4_h_r_9')
// (16, 1, 'sp4_r_v_b_13')
// (16, 2, 'sp4_r_v_b_0')
// (16, 4, 'local_g1_4')
// (16, 4, 'lutff_2/in_3')
// (16, 4, 'lutff_7/in_2')
// (16, 4, 'sp4_h_r_20')
// (17, 0, 'span4_horz_r_2')
// (17, 0, 'span4_vert_13')
// (17, 1, 'sp4_r_v_b_37')
// (17, 1, 'sp4_v_b_13')
// (17, 2, 'local_g0_0')
// (17, 2, 'lutff_3/in_1')
// (17, 2, 'lutff_7/in_1')
// (17, 2, 'sp4_r_v_b_24')
// (17, 2, 'sp4_v_b_0')
// (17, 3, 'local_g2_5')
// (17, 3, 'lutff_4/in_3')
// (17, 3, 'lutff_6/in_3')
// (17, 3, 'lutff_7/in_0')
// (17, 3, 'sp4_r_v_b_13')
// (17, 4, 'sp4_h_r_33')
// (17, 4, 'sp4_r_v_b_0')
// (18, 0, 'span4_horz_r_2')
// (18, 0, 'span4_horz_r_6')
// (18, 0, 'span4_vert_37')
// (18, 1, 'neigh_op_bnr_2')
// (18, 1, 'neigh_op_bnr_6')
// (18, 1, 'sp4_r_v_b_12')
// (18, 1, 'sp4_r_v_b_44')
// (18, 1, 'sp4_v_b_37')
// (18, 2, 'sp4_r_v_b_1')
// (18, 2, 'sp4_r_v_b_33')
// (18, 2, 'sp4_v_b_24')
// (18, 3, 'sp4_r_v_b_20')
// (18, 3, 'sp4_v_b_13')
// (18, 4, 'sp4_h_r_44')
// (18, 4, 'sp4_r_v_b_9')
// (18, 4, 'sp4_v_b_0')
// (19, 0, 'io_1/D_IN_0')
// (19, 0, 'io_1/PAD')
// (19, 0, 'span4_horz_r_10')
// (19, 0, 'span4_horz_r_6')
// (19, 0, 'span4_vert_12')
// (19, 0, 'span4_vert_44')
// (19, 1, 'neigh_op_bot_2')
// (19, 1, 'neigh_op_bot_6')
// (19, 1, 'sp4_v_b_12')
// (19, 1, 'sp4_v_b_44')
// (19, 2, 'sp4_h_r_1')
// (19, 2, 'sp4_h_r_7')
// (19, 2, 'sp4_v_b_1')
// (19, 2, 'sp4_v_b_33')
// (19, 3, 'sp4_v_b_20')
// (19, 4, 'sp4_h_l_44')
// (19, 4, 'sp4_v_b_9')
// (20, 0, 'span4_horz_r_10')
// (20, 0, 'span4_horz_r_14')
// (20, 1, 'neigh_op_bnl_2')
// (20, 1, 'neigh_op_bnl_6')
// (20, 2, 'local_g1_2')
// (20, 2, 'lutff_6/in_3')
// (20, 2, 'sp4_h_r_12')
// (20, 2, 'sp4_h_r_18')
// (21, 0, 'span4_horz_l_14')
// (21, 0, 'span4_horz_r_14')
// (21, 2, 'local_g3_1')
// (21, 2, 'lutff_1/in_3')
// (21, 2, 'lutff_4/in_0')
// (21, 2, 'sp4_h_r_25')
// (21, 2, 'sp4_h_r_31')
// (22, 0, 'span4_horz_l_14')
// (22, 2, 'local_g2_2')
// (22, 2, 'local_g3_4')
// (22, 2, 'lutff_0/in_1')
// (22, 2, 'lutff_1/in_0')
// (22, 2, 'lutff_6/in_0')
// (22, 2, 'sp4_h_r_36')
// (22, 2, 'sp4_h_r_42')
// (23, 2, 'sp4_h_l_36')
// (23, 2, 'sp4_h_l_42')

wire n2184;
// (15, 5, 'neigh_op_tnr_0')
// (15, 6, 'neigh_op_rgt_0')
// (15, 7, 'neigh_op_bnr_0')
// (16, 5, 'neigh_op_top_0')
// (16, 6, 'local_g2_0')
// (16, 6, 'lutff_0/out')
// (16, 6, 'lutff_1/in_3')
// (16, 7, 'neigh_op_bot_0')
// (17, 5, 'neigh_op_tnl_0')
// (17, 6, 'neigh_op_lft_0')
// (17, 7, 'neigh_op_bnl_0')

wire n2185;
// (15, 5, 'neigh_op_tnr_1')
// (15, 6, 'neigh_op_rgt_1')
// (15, 7, 'local_g0_1')
// (15, 7, 'lutff_0/in_1')
// (15, 7, 'neigh_op_bnr_1')
// (16, 5, 'neigh_op_top_1')
// (16, 6, 'lutff_1/out')
// (16, 7, 'neigh_op_bot_1')
// (17, 5, 'neigh_op_tnl_1')
// (17, 6, 'neigh_op_lft_1')
// (17, 7, 'neigh_op_bnl_1')

wire n2186;
// (15, 5, 'neigh_op_tnr_2')
// (15, 6, 'neigh_op_rgt_2')
// (15, 7, 'neigh_op_bnr_2')
// (16, 5, 'neigh_op_top_2')
// (16, 6, 'local_g3_2')
// (16, 6, 'lutff_1/in_2')
// (16, 6, 'lutff_2/out')
// (16, 7, 'neigh_op_bot_2')
// (17, 5, 'neigh_op_tnl_2')
// (17, 6, 'neigh_op_lft_2')
// (17, 7, 'neigh_op_bnl_2')

wire n2187;
// (15, 5, 'neigh_op_tnr_4')
// (15, 6, 'neigh_op_rgt_4')
// (15, 7, 'neigh_op_bnr_4')
// (16, 5, 'neigh_op_top_4')
// (16, 6, 'local_g3_4')
// (16, 6, 'lutff_1/in_0')
// (16, 6, 'lutff_4/out')
// (16, 7, 'neigh_op_bot_4')
// (17, 5, 'neigh_op_tnl_4')
// (17, 6, 'neigh_op_lft_4')
// (17, 7, 'neigh_op_bnl_4')

wire n2188;
// (15, 5, 'neigh_op_tnr_6')
// (15, 6, 'neigh_op_rgt_6')
// (15, 7, 'neigh_op_bnr_6')
// (16, 5, 'local_g1_6')
// (16, 5, 'lutff_1/in_2')
// (16, 5, 'neigh_op_top_6')
// (16, 6, 'lutff_6/out')
// (16, 7, 'neigh_op_bot_6')
// (17, 5, 'neigh_op_tnl_6')
// (17, 6, 'neigh_op_lft_6')
// (17, 7, 'neigh_op_bnl_6')

wire n2189;
// (15, 5, 'neigh_op_tnr_7')
// (15, 6, 'neigh_op_rgt_7')
// (15, 7, 'neigh_op_bnr_7')
// (16, 5, 'neigh_op_top_7')
// (16, 6, 'local_g3_7')
// (16, 6, 'lutff_1/in_1')
// (16, 6, 'lutff_7/out')
// (16, 7, 'neigh_op_bot_7')
// (17, 5, 'neigh_op_tnl_7')
// (17, 6, 'neigh_op_lft_7')
// (17, 7, 'neigh_op_bnl_7')

reg n2190 = 0;
// (15, 5, 'sp4_h_r_6')
// (16, 4, 'neigh_op_tnr_7')
// (16, 5, 'neigh_op_rgt_7')
// (16, 5, 'sp4_h_r_19')
// (16, 6, 'neigh_op_bnr_7')
// (17, 4, 'neigh_op_top_7')
// (17, 5, 'lutff_7/out')
// (17, 5, 'sp4_h_r_30')
// (17, 6, 'neigh_op_bot_7')
// (18, 4, 'neigh_op_tnl_7')
// (18, 5, 'neigh_op_lft_7')
// (18, 5, 'sp4_h_r_43')
// (18, 6, 'neigh_op_bnl_7')
// (19, 5, 'local_g1_6')
// (19, 5, 'ram/WDATA_15')
// (19, 5, 'sp4_h_l_43')
// (19, 5, 'sp4_h_r_6')
// (20, 5, 'sp4_h_r_19')
// (21, 5, 'sp4_h_r_30')
// (22, 5, 'sp4_h_r_43')
// (23, 5, 'sp4_h_l_43')

wire n2191;
// (15, 5, 'sp4_r_v_b_47')
// (15, 6, 'local_g2_2')
// (15, 6, 'lutff_global/cen')
// (15, 6, 'sp4_r_v_b_34')
// (15, 7, 'sp4_r_v_b_23')
// (15, 8, 'sp4_r_v_b_10')
// (15, 9, 'sp4_r_v_b_42')
// (15, 10, 'sp4_r_v_b_31')
// (15, 11, 'sp4_r_v_b_18')
// (15, 12, 'sp4_r_v_b_7')
// (16, 4, 'sp4_v_t_47')
// (16, 5, 'sp4_v_b_47')
// (16, 6, 'sp4_r_v_b_38')
// (16, 6, 'sp4_v_b_34')
// (16, 7, 'sp4_r_v_b_27')
// (16, 7, 'sp4_v_b_23')
// (16, 8, 'sp4_r_v_b_14')
// (16, 8, 'sp4_v_b_10')
// (16, 8, 'sp4_v_t_42')
// (16, 9, 'sp4_r_v_b_3')
// (16, 9, 'sp4_v_b_42')
// (16, 10, 'sp4_r_v_b_42')
// (16, 10, 'sp4_v_b_31')
// (16, 11, 'neigh_op_tnr_1')
// (16, 11, 'sp4_r_v_b_31')
// (16, 11, 'sp4_v_b_18')
// (16, 12, 'neigh_op_rgt_1')
// (16, 12, 'sp4_h_r_7')
// (16, 12, 'sp4_r_v_b_18')
// (16, 12, 'sp4_v_b_7')
// (16, 13, 'neigh_op_bnr_1')
// (16, 13, 'sp4_r_v_b_7')
// (17, 2, 'sp4_r_v_b_39')
// (17, 3, 'sp4_r_v_b_26')
// (17, 4, 'sp4_r_v_b_15')
// (17, 5, 'sp4_r_v_b_2')
// (17, 5, 'sp4_v_t_38')
// (17, 6, 'sp4_r_v_b_43')
// (17, 6, 'sp4_v_b_38')
// (17, 7, 'local_g3_3')
// (17, 7, 'lutff_global/cen')
// (17, 7, 'sp4_r_v_b_30')
// (17, 7, 'sp4_v_b_27')
// (17, 8, 'sp4_r_v_b_19')
// (17, 8, 'sp4_v_b_14')
// (17, 9, 'sp4_r_v_b_6')
// (17, 9, 'sp4_v_b_3')
// (17, 9, 'sp4_v_t_42')
// (17, 10, 'sp4_r_v_b_43')
// (17, 10, 'sp4_v_b_42')
// (17, 11, 'neigh_op_top_1')
// (17, 11, 'sp4_r_v_b_30')
// (17, 11, 'sp4_v_b_31')
// (17, 12, 'lutff_1/out')
// (17, 12, 'sp4_h_r_18')
// (17, 12, 'sp4_r_v_b_19')
// (17, 12, 'sp4_v_b_18')
// (17, 13, 'neigh_op_bot_1')
// (17, 13, 'sp4_r_v_b_6')
// (17, 13, 'sp4_v_b_7')
// (18, 1, 'sp4_v_t_39')
// (18, 2, 'sp4_v_b_39')
// (18, 3, 'local_g2_2')
// (18, 3, 'lutff_global/cen')
// (18, 3, 'sp4_v_b_26')
// (18, 4, 'sp4_v_b_15')
// (18, 5, 'sp4_v_b_2')
// (18, 5, 'sp4_v_t_43')
// (18, 6, 'sp4_v_b_43')
// (18, 7, 'sp4_v_b_30')
// (18, 8, 'sp4_v_b_19')
// (18, 9, 'sp4_v_b_6')
// (18, 9, 'sp4_v_t_43')
// (18, 10, 'sp4_v_b_43')
// (18, 11, 'neigh_op_tnl_1')
// (18, 11, 'sp4_v_b_30')
// (18, 12, 'neigh_op_lft_1')
// (18, 12, 'sp4_h_r_31')
// (18, 12, 'sp4_v_b_19')
// (18, 13, 'neigh_op_bnl_1')
// (18, 13, 'sp4_v_b_6')
// (19, 12, 'sp4_h_r_42')
// (20, 12, 'sp4_h_l_42')

reg n2192 = 0;
// (15, 6, 'local_g0_1')
// (15, 6, 'lutff_5/in_0')
// (15, 6, 'sp4_h_r_9')
// (16, 6, 'sp4_h_r_20')
// (17, 6, 'sp4_h_r_33')
// (18, 6, 'sp4_h_r_44')
// (19, 6, 'sp4_h_l_44')
// (19, 6, 'sp4_h_r_6')
// (20, 5, 'neigh_op_tnr_7')
// (20, 6, 'neigh_op_rgt_7')
// (20, 6, 'sp4_h_r_19')
// (20, 6, 'sp4_r_v_b_46')
// (20, 7, 'neigh_op_bnr_7')
// (20, 7, 'sp4_r_v_b_35')
// (20, 8, 'sp4_r_v_b_22')
// (20, 9, 'sp4_r_v_b_11')
// (21, 5, 'neigh_op_top_7')
// (21, 5, 'sp4_v_t_46')
// (21, 6, 'lutff_7/out')
// (21, 6, 'sp4_h_r_30')
// (21, 6, 'sp4_v_b_46')
// (21, 7, 'neigh_op_bot_7')
// (21, 7, 'sp4_v_b_35')
// (21, 8, 'sp4_v_b_22')
// (21, 9, 'local_g0_3')
// (21, 9, 'lutff_7/in_2')
// (21, 9, 'sp4_v_b_11')
// (22, 5, 'neigh_op_tnl_7')
// (22, 6, 'neigh_op_lft_7')
// (22, 6, 'sp4_h_r_43')
// (22, 7, 'neigh_op_bnl_7')
// (23, 6, 'sp4_h_l_43')

wire n2193;
// (15, 6, 'local_g0_2')
// (15, 6, 'lutff_3/in_3')
// (15, 6, 'sp4_h_r_2')
// (16, 5, 'neigh_op_tnr_5')
// (16, 6, 'neigh_op_rgt_5')
// (16, 6, 'sp4_h_r_15')
// (16, 7, 'neigh_op_bnr_5')
// (17, 5, 'neigh_op_top_5')
// (17, 6, 'lutff_5/out')
// (17, 6, 'sp4_h_r_26')
// (17, 7, 'neigh_op_bot_5')
// (18, 5, 'neigh_op_tnl_5')
// (18, 6, 'neigh_op_lft_5')
// (18, 6, 'sp4_h_r_39')
// (18, 7, 'neigh_op_bnl_5')
// (19, 6, 'sp4_h_l_39')

reg n2194 = 0;
// (15, 6, 'local_g0_5')
// (15, 6, 'lutff_0/in_1')
// (15, 6, 'sp4_h_r_5')
// (16, 1, 'sp4_r_v_b_17')
// (16, 2, 'sp4_r_v_b_4')
// (16, 6, 'sp4_h_r_16')
// (17, 0, 'span4_vert_17')
// (17, 1, 'local_g0_1')
// (17, 1, 'lutff_5/in_0')
// (17, 1, 'sp4_v_b_17')
// (17, 2, 'sp4_h_r_4')
// (17, 2, 'sp4_v_b_4')
// (17, 6, 'sp4_h_r_29')
// (18, 2, 'sp4_h_r_17')
// (18, 6, 'sp4_h_r_40')
// (19, 2, 'sp4_h_r_28')
// (19, 6, 'sp4_h_l_40')
// (19, 6, 'sp4_h_r_2')
// (20, 2, 'sp4_h_r_41')
// (20, 3, 'sp4_r_v_b_47')
// (20, 4, 'sp4_r_v_b_34')
// (20, 5, 'neigh_op_tnr_5')
// (20, 5, 'sp4_r_v_b_23')
// (20, 6, 'neigh_op_rgt_5')
// (20, 6, 'sp4_h_r_15')
// (20, 6, 'sp4_r_v_b_10')
// (20, 7, 'neigh_op_bnr_5')
// (21, 2, 'sp4_h_l_41')
// (21, 2, 'sp4_v_t_47')
// (21, 3, 'sp4_v_b_47')
// (21, 4, 'sp4_v_b_34')
// (21, 5, 'neigh_op_top_5')
// (21, 5, 'sp4_v_b_23')
// (21, 6, 'lutff_5/out')
// (21, 6, 'sp4_h_r_26')
// (21, 6, 'sp4_v_b_10')
// (21, 7, 'neigh_op_bot_5')
// (22, 5, 'neigh_op_tnl_5')
// (22, 6, 'neigh_op_lft_5')
// (22, 6, 'sp4_h_r_39')
// (22, 7, 'neigh_op_bnl_5')
// (23, 6, 'sp4_h_l_39')

reg n2195 = 0;
// (15, 6, 'local_g1_0')
// (15, 6, 'lutff_4/in_1')
// (15, 6, 'sp12_h_r_0')
// (16, 6, 'sp12_h_r_3')
// (17, 6, 'sp12_h_r_4')
// (18, 6, 'sp12_h_r_7')
// (19, 6, 'sp12_h_r_8')
// (20, 5, 'neigh_op_tnr_2')
// (20, 6, 'neigh_op_rgt_2')
// (20, 6, 'sp12_h_r_11')
// (20, 7, 'neigh_op_bnr_2')
// (21, 5, 'neigh_op_top_2')
// (21, 6, 'lutff_2/out')
// (21, 6, 'sp12_h_r_12')
// (21, 7, 'neigh_op_bot_2')
// (22, 5, 'neigh_op_tnl_2')
// (22, 6, 'local_g1_2')
// (22, 6, 'lutff_7/in_2')
// (22, 6, 'neigh_op_lft_2')
// (22, 6, 'sp12_h_r_15')
// (22, 7, 'neigh_op_bnl_2')
// (23, 6, 'sp12_h_r_16')
// (24, 6, 'sp12_h_r_19')
// (25, 6, 'sp12_h_r_20')

reg n2196 = 0;
// (15, 6, 'local_g1_1')
// (15, 6, 'lutff_5/in_3')
// (15, 6, 'sp4_h_r_1')
// (16, 6, 'sp4_h_r_12')
// (17, 3, 'sp4_r_v_b_44')
// (17, 4, 'sp4_r_v_b_33')
// (17, 5, 'sp4_r_v_b_20')
// (17, 6, 'local_g2_1')
// (17, 6, 'lutff_0/in_1')
// (17, 6, 'sp4_h_r_25')
// (17, 6, 'sp4_r_v_b_9')
// (18, 2, 'sp4_v_t_44')
// (18, 3, 'sp4_v_b_44')
// (18, 4, 'sp4_v_b_33')
// (18, 5, 'sp4_v_b_20')
// (18, 6, 'sp4_h_r_36')
// (18, 6, 'sp4_h_r_4')
// (18, 6, 'sp4_v_b_9')
// (19, 6, 'sp4_h_l_36')
// (19, 6, 'sp4_h_r_17')
// (19, 6, 'sp4_h_r_5')
// (20, 6, 'sp4_h_r_16')
// (20, 6, 'sp4_h_r_28')
// (21, 6, 'sp4_h_r_29')
// (21, 6, 'sp4_h_r_41')
// (21, 7, 'sp4_r_v_b_47')
// (21, 8, 'sp4_r_v_b_34')
// (21, 9, 'neigh_op_tnr_5')
// (21, 9, 'sp4_r_v_b_23')
// (21, 10, 'neigh_op_rgt_5')
// (21, 10, 'sp4_r_v_b_10')
// (21, 11, 'neigh_op_bnr_5')
// (22, 6, 'sp4_h_l_41')
// (22, 6, 'sp4_h_r_40')
// (22, 6, 'sp4_v_t_47')
// (22, 7, 'sp4_r_v_b_46')
// (22, 7, 'sp4_v_b_47')
// (22, 8, 'sp4_r_v_b_35')
// (22, 8, 'sp4_v_b_34')
// (22, 9, 'neigh_op_top_5')
// (22, 9, 'sp4_r_v_b_22')
// (22, 9, 'sp4_v_b_23')
// (22, 10, 'lutff_5/out')
// (22, 10, 'sp4_r_v_b_11')
// (22, 10, 'sp4_v_b_10')
// (22, 11, 'neigh_op_bot_5')
// (23, 6, 'sp4_h_l_40')
// (23, 6, 'sp4_v_t_46')
// (23, 7, 'sp4_v_b_46')
// (23, 8, 'sp4_v_b_35')
// (23, 9, 'neigh_op_tnl_5')
// (23, 9, 'sp4_v_b_22')
// (23, 10, 'neigh_op_lft_5')
// (23, 10, 'sp4_v_b_11')
// (23, 11, 'neigh_op_bnl_5')

reg n2197 = 0;
// (15, 6, 'local_g1_4')
// (15, 6, 'lutff_3/in_0')
// (15, 6, 'sp4_h_r_4')
// (16, 6, 'sp4_h_r_17')
// (17, 6, 'sp4_h_r_28')
// (18, 6, 'sp4_h_r_41')
// (19, 6, 'sp4_h_l_41')
// (19, 6, 'sp4_h_r_8')
// (20, 5, 'neigh_op_tnr_0')
// (20, 5, 'sp4_r_v_b_45')
// (20, 6, 'neigh_op_rgt_0')
// (20, 6, 'sp4_h_r_21')
// (20, 6, 'sp4_r_v_b_32')
// (20, 7, 'neigh_op_bnr_0')
// (20, 7, 'sp4_r_v_b_21')
// (20, 8, 'local_g2_0')
// (20, 8, 'lutff_6/in_2')
// (20, 8, 'sp4_r_v_b_8')
// (21, 4, 'sp4_v_t_45')
// (21, 5, 'neigh_op_top_0')
// (21, 5, 'sp4_v_b_45')
// (21, 6, 'lutff_0/out')
// (21, 6, 'sp4_h_r_32')
// (21, 6, 'sp4_v_b_32')
// (21, 7, 'neigh_op_bot_0')
// (21, 7, 'sp4_v_b_21')
// (21, 8, 'sp4_v_b_8')
// (22, 5, 'neigh_op_tnl_0')
// (22, 6, 'neigh_op_lft_0')
// (22, 6, 'sp4_h_r_45')
// (22, 7, 'neigh_op_bnl_0')
// (23, 6, 'sp4_h_l_45')

wire n2198;
// (15, 6, 'neigh_op_tnr_0')
// (15, 7, 'neigh_op_rgt_0')
// (15, 8, 'neigh_op_bnr_0')
// (16, 6, 'neigh_op_top_0')
// (16, 7, 'lutff_0/out')
// (16, 8, 'local_g1_0')
// (16, 8, 'lutff_5/in_2')
// (16, 8, 'neigh_op_bot_0')
// (17, 6, 'neigh_op_tnl_0')
// (17, 7, 'neigh_op_lft_0')
// (17, 8, 'neigh_op_bnl_0')

reg n2199 = 0;
// (15, 6, 'neigh_op_tnr_2')
// (15, 7, 'neigh_op_rgt_2')
// (15, 7, 'sp4_r_v_b_36')
// (15, 8, 'neigh_op_bnr_2')
// (15, 8, 'sp4_r_v_b_25')
// (15, 9, 'sp4_r_v_b_12')
// (15, 10, 'sp4_r_v_b_1')
// (16, 6, 'neigh_op_top_2')
// (16, 6, 'sp4_v_t_36')
// (16, 7, 'lutff_2/out')
// (16, 7, 'sp4_v_b_36')
// (16, 8, 'neigh_op_bot_2')
// (16, 8, 'sp4_v_b_25')
// (16, 9, 'local_g0_4')
// (16, 9, 'lutff_1/in_1')
// (16, 9, 'sp4_v_b_12')
// (16, 10, 'sp4_v_b_1')
// (17, 6, 'neigh_op_tnl_2')
// (17, 7, 'neigh_op_lft_2')
// (17, 8, 'neigh_op_bnl_2')

wire n2200;
// (15, 6, 'neigh_op_tnr_4')
// (15, 7, 'neigh_op_rgt_4')
// (15, 8, 'neigh_op_bnr_4')
// (16, 6, 'neigh_op_top_4')
// (16, 7, 'lutff_4/out')
// (16, 8, 'local_g1_4')
// (16, 8, 'lutff_0/in_1')
// (16, 8, 'neigh_op_bot_4')
// (17, 6, 'neigh_op_tnl_4')
// (17, 7, 'neigh_op_lft_4')
// (17, 8, 'neigh_op_bnl_4')

wire n2201;
// (15, 6, 'neigh_op_tnr_5')
// (15, 7, 'neigh_op_rgt_5')
// (15, 8, 'neigh_op_bnr_5')
// (16, 6, 'neigh_op_top_5')
// (16, 7, 'local_g2_5')
// (16, 7, 'lutff_0/in_1')
// (16, 7, 'lutff_5/out')
// (16, 8, 'neigh_op_bot_5')
// (17, 6, 'neigh_op_tnl_5')
// (17, 7, 'neigh_op_lft_5')
// (17, 8, 'neigh_op_bnl_5')

reg n2202 = 0;
// (15, 6, 'neigh_op_tnr_6')
// (15, 7, 'neigh_op_rgt_6')
// (15, 8, 'neigh_op_bnr_6')
// (16, 6, 'neigh_op_top_6')
// (16, 6, 'sp4_r_v_b_40')
// (16, 7, 'lutff_6/out')
// (16, 7, 'sp4_r_v_b_29')
// (16, 8, 'neigh_op_bot_6')
// (16, 8, 'sp4_r_v_b_16')
// (16, 9, 'sp4_r_v_b_5')
// (17, 5, 'sp4_v_t_40')
// (17, 6, 'neigh_op_tnl_6')
// (17, 6, 'sp4_v_b_40')
// (17, 7, 'neigh_op_lft_6')
// (17, 7, 'sp4_v_b_29')
// (17, 8, 'neigh_op_bnl_6')
// (17, 8, 'sp4_v_b_16')
// (17, 9, 'local_g1_5')
// (17, 9, 'lutff_4/in_0')
// (17, 9, 'sp4_v_b_5')

wire n2203;
// (15, 6, 'neigh_op_tnr_7')
// (15, 7, 'neigh_op_rgt_7')
// (15, 8, 'neigh_op_bnr_7')
// (16, 6, 'neigh_op_top_7')
// (16, 7, 'lutff_7/out')
// (16, 8, 'local_g1_7')
// (16, 8, 'lutff_6/in_0')
// (16, 8, 'neigh_op_bot_7')
// (17, 6, 'neigh_op_tnl_7')
// (17, 7, 'neigh_op_lft_7')
// (17, 8, 'neigh_op_bnl_7')

reg n2204 = 0;
// (15, 6, 'sp4_r_v_b_47')
// (15, 7, 'local_g2_2')
// (15, 7, 'lutff_5/in_3')
// (15, 7, 'sp4_r_v_b_34')
// (15, 8, 'local_g3_7')
// (15, 8, 'lutff_4/in_0')
// (15, 8, 'sp4_r_v_b_23')
// (15, 9, 'sp4_r_v_b_10')
// (15, 9, 'sp4_r_v_b_38')
// (15, 10, 'sp4_r_v_b_27')
// (15, 10, 'sp4_r_v_b_47')
// (15, 11, 'sp4_r_v_b_14')
// (15, 11, 'sp4_r_v_b_34')
// (15, 12, 'local_g3_5')
// (15, 12, 'lutff_6/in_0')
// (15, 12, 'neigh_op_tnr_5')
// (15, 12, 'sp4_r_v_b_23')
// (15, 12, 'sp4_r_v_b_3')
// (15, 13, 'neigh_op_rgt_5')
// (15, 13, 'sp4_r_v_b_10')
// (15, 13, 'sp4_r_v_b_42')
// (15, 14, 'neigh_op_bnr_5')
// (15, 14, 'sp4_r_v_b_31')
// (15, 15, 'sp4_r_v_b_18')
// (15, 16, 'sp4_r_v_b_7')
// (16, 5, 'sp4_v_t_47')
// (16, 6, 'sp4_v_b_47')
// (16, 7, 'local_g3_2')
// (16, 7, 'lutff_6/in_3')
// (16, 7, 'sp4_v_b_34')
// (16, 8, 'sp4_h_r_3')
// (16, 8, 'sp4_r_v_b_43')
// (16, 8, 'sp4_v_b_23')
// (16, 8, 'sp4_v_t_38')
// (16, 9, 'sp4_r_v_b_30')
// (16, 9, 'sp4_v_b_10')
// (16, 9, 'sp4_v_b_38')
// (16, 9, 'sp4_v_t_47')
// (16, 10, 'local_g2_7')
// (16, 10, 'lutff_0/in_3')
// (16, 10, 'sp4_r_v_b_19')
// (16, 10, 'sp4_v_b_27')
// (16, 10, 'sp4_v_b_47')
// (16, 11, 'sp4_r_v_b_6')
// (16, 11, 'sp4_v_b_14')
// (16, 11, 'sp4_v_b_34')
// (16, 12, 'neigh_op_top_5')
// (16, 12, 'sp4_r_v_b_38')
// (16, 12, 'sp4_v_b_23')
// (16, 12, 'sp4_v_b_3')
// (16, 12, 'sp4_v_t_42')
// (16, 13, 'lutff_5/out')
// (16, 13, 'sp4_r_v_b_27')
// (16, 13, 'sp4_v_b_10')
// (16, 13, 'sp4_v_b_42')
// (16, 14, 'neigh_op_bot_5')
// (16, 14, 'sp4_r_v_b_14')
// (16, 14, 'sp4_v_b_31')
// (16, 15, 'sp4_r_v_b_3')
// (16, 15, 'sp4_v_b_18')
// (16, 16, 'sp4_v_b_7')
// (17, 7, 'sp4_h_r_6')
// (17, 7, 'sp4_v_t_43')
// (17, 8, 'local_g2_3')
// (17, 8, 'lutff_0/in_1')
// (17, 8, 'sp4_h_r_14')
// (17, 8, 'sp4_v_b_43')
// (17, 9, 'sp4_v_b_30')
// (17, 10, 'local_g0_3')
// (17, 10, 'lutff_7/in_0')
// (17, 10, 'sp4_v_b_19')
// (17, 11, 'sp4_v_b_6')
// (17, 11, 'sp4_v_t_38')
// (17, 12, 'neigh_op_tnl_5')
// (17, 12, 'sp4_v_b_38')
// (17, 13, 'neigh_op_lft_5')
// (17, 13, 'sp4_v_b_27')
// (17, 14, 'neigh_op_bnl_5')
// (17, 14, 'sp4_v_b_14')
// (17, 15, 'sp4_v_b_3')
// (18, 7, 'local_g0_3')
// (18, 7, 'lutff_2/in_3')
// (18, 7, 'sp4_h_r_19')
// (18, 8, 'local_g2_3')
// (18, 8, 'lutff_7/in_0')
// (18, 8, 'sp4_h_r_27')
// (19, 7, 'sp4_h_r_30')
// (19, 8, 'sp4_h_r_38')
// (20, 7, 'sp4_h_r_43')
// (20, 8, 'sp4_h_l_38')
// (21, 7, 'sp4_h_l_43')

wire n2205;
// (15, 7, 'neigh_op_tnr_0')
// (15, 8, 'neigh_op_rgt_0')
// (15, 9, 'neigh_op_bnr_0')
// (16, 7, 'neigh_op_top_0')
// (16, 8, 'local_g0_0')
// (16, 8, 'lutff_0/out')
// (16, 8, 'lutff_5/in_1')
// (16, 9, 'neigh_op_bot_0')
// (17, 7, 'neigh_op_tnl_0')
// (17, 8, 'neigh_op_lft_0')
// (17, 9, 'neigh_op_bnl_0')

wire n2206;
// (15, 7, 'neigh_op_tnr_1')
// (15, 8, 'neigh_op_rgt_1')
// (15, 9, 'neigh_op_bnr_1')
// (16, 7, 'neigh_op_top_1')
// (16, 8, 'local_g1_1')
// (16, 8, 'lutff_1/out')
// (16, 8, 'lutff_5/in_3')
// (16, 9, 'neigh_op_bot_1')
// (17, 7, 'neigh_op_tnl_1')
// (17, 8, 'neigh_op_lft_1')
// (17, 9, 'neigh_op_bnl_1')

reg n2207 = 0;
// (15, 7, 'neigh_op_tnr_2')
// (15, 8, 'neigh_op_rgt_2')
// (15, 9, 'neigh_op_bnr_2')
// (16, 7, 'neigh_op_top_2')
// (16, 8, 'lutff_2/out')
// (16, 9, 'local_g1_2')
// (16, 9, 'lutff_1/in_0')
// (16, 9, 'neigh_op_bot_2')
// (17, 7, 'neigh_op_tnl_2')
// (17, 8, 'neigh_op_lft_2')
// (17, 9, 'neigh_op_bnl_2')

wire n2208;
// (15, 7, 'neigh_op_tnr_3')
// (15, 8, 'neigh_op_rgt_3')
// (15, 9, 'neigh_op_bnr_3')
// (16, 7, 'neigh_op_top_3')
// (16, 8, 'local_g2_3')
// (16, 8, 'lutff_3/out')
// (16, 8, 'lutff_5/in_0')
// (16, 9, 'neigh_op_bot_3')
// (17, 7, 'neigh_op_tnl_3')
// (17, 8, 'neigh_op_lft_3')
// (17, 9, 'neigh_op_bnl_3')

wire n2209;
// (15, 7, 'neigh_op_tnr_4')
// (15, 8, 'neigh_op_rgt_4')
// (15, 9, 'local_g0_4')
// (15, 9, 'lutff_4/in_0')
// (15, 9, 'neigh_op_bnr_4')
// (16, 7, 'neigh_op_top_4')
// (16, 8, 'lutff_4/out')
// (16, 9, 'neigh_op_bot_4')
// (17, 7, 'neigh_op_tnl_4')
// (17, 8, 'neigh_op_lft_4')
// (17, 9, 'neigh_op_bnl_4')

wire n2210;
// (15, 7, 'neigh_op_tnr_5')
// (15, 7, 'sp4_r_v_b_39')
// (15, 8, 'neigh_op_rgt_5')
// (15, 8, 'sp4_r_v_b_26')
// (15, 9, 'neigh_op_bnr_5')
// (15, 9, 'sp4_r_v_b_15')
// (15, 10, 'local_g1_2')
// (15, 10, 'lutff_4/in_1')
// (15, 10, 'sp4_r_v_b_2')
// (16, 6, 'sp4_v_t_39')
// (16, 7, 'neigh_op_top_5')
// (16, 7, 'sp4_v_b_39')
// (16, 8, 'lutff_5/out')
// (16, 8, 'sp4_v_b_26')
// (16, 9, 'neigh_op_bot_5')
// (16, 9, 'sp4_v_b_15')
// (16, 10, 'sp4_v_b_2')
// (17, 7, 'neigh_op_tnl_5')
// (17, 8, 'neigh_op_lft_5')
// (17, 9, 'neigh_op_bnl_5')

wire n2211;
// (15, 7, 'neigh_op_tnr_6')
// (15, 8, 'neigh_op_rgt_6')
// (15, 9, 'local_g1_6')
// (15, 9, 'lutff_6/in_1')
// (15, 9, 'neigh_op_bnr_6')
// (16, 7, 'neigh_op_top_6')
// (16, 8, 'lutff_6/out')
// (16, 9, 'neigh_op_bot_6')
// (17, 7, 'neigh_op_tnl_6')
// (17, 8, 'neigh_op_lft_6')
// (17, 9, 'neigh_op_bnl_6')

reg n2212 = 0;
// (15, 7, 'neigh_op_tnr_7')
// (15, 8, 'neigh_op_rgt_7')
// (15, 9, 'neigh_op_bnr_7')
// (16, 7, 'neigh_op_top_7')
// (16, 8, 'lutff_7/out')
// (16, 9, 'local_g0_7')
// (16, 9, 'lutff_2/in_3')
// (16, 9, 'neigh_op_bot_7')
// (17, 7, 'neigh_op_tnl_7')
// (17, 8, 'neigh_op_lft_7')
// (17, 9, 'neigh_op_bnl_7')

wire n2213;
// (15, 7, 'sp4_r_v_b_43')
// (15, 8, 'sp4_r_v_b_30')
// (15, 9, 'local_g3_3')
// (15, 9, 'lutff_global/cen')
// (15, 9, 'sp4_r_v_b_19')
// (15, 10, 'sp4_r_v_b_6')
// (16, 6, 'sp4_h_r_6')
// (16, 6, 'sp4_v_t_43')
// (16, 7, 'sp4_v_b_43')
// (16, 8, 'sp4_v_b_30')
// (16, 9, 'sp4_v_b_19')
// (16, 10, 'sp12_h_r_0')
// (16, 10, 'sp4_v_b_6')
// (17, 6, 'sp4_h_r_19')
// (17, 10, 'local_g1_3')
// (17, 10, 'lutff_global/cen')
// (17, 10, 'sp12_h_r_3')
// (18, 6, 'sp4_h_r_30')
// (18, 10, 'sp12_h_r_4')
// (19, 6, 'sp4_h_r_43')
// (19, 7, 'sp4_r_v_b_37')
// (19, 8, 'sp4_r_v_b_24')
// (19, 9, 'neigh_op_tnr_0')
// (19, 9, 'sp4_r_v_b_13')
// (19, 10, 'neigh_op_rgt_0')
// (19, 10, 'sp12_h_r_7')
// (19, 10, 'sp4_r_v_b_0')
// (19, 11, 'neigh_op_bnr_0')
// (20, 6, 'sp4_h_l_43')
// (20, 6, 'sp4_v_t_37')
// (20, 7, 'sp4_v_b_37')
// (20, 8, 'sp4_r_v_b_41')
// (20, 8, 'sp4_v_b_24')
// (20, 9, 'neigh_op_top_0')
// (20, 9, 'sp4_r_v_b_28')
// (20, 9, 'sp4_v_b_13')
// (20, 10, 'lutff_0/out')
// (20, 10, 'sp12_h_r_8')
// (20, 10, 'sp4_r_v_b_17')
// (20, 10, 'sp4_v_b_0')
// (20, 11, 'neigh_op_bot_0')
// (20, 11, 'sp4_r_v_b_4')
// (21, 7, 'sp4_v_t_41')
// (21, 8, 'sp4_v_b_41')
// (21, 9, 'neigh_op_tnl_0')
// (21, 9, 'sp4_v_b_28')
// (21, 10, 'neigh_op_lft_0')
// (21, 10, 'sp12_h_r_11')
// (21, 10, 'sp4_v_b_17')
// (21, 11, 'local_g0_2')
// (21, 11, 'lutff_global/cen')
// (21, 11, 'neigh_op_bnl_0')
// (21, 11, 'sp4_h_r_10')
// (21, 11, 'sp4_v_b_4')
// (22, 10, 'sp12_h_r_12')
// (22, 11, 'sp4_h_r_23')
// (23, 10, 'sp12_h_r_15')
// (23, 11, 'sp4_h_r_34')
// (24, 10, 'sp12_h_r_16')
// (24, 11, 'sp4_h_r_47')
// (25, 10, 'sp12_h_r_19')
// (25, 11, 'sp4_h_l_47')

wire n2214;
// (15, 8, 'neigh_op_tnr_0')
// (15, 9, 'neigh_op_rgt_0')
// (15, 10, 'neigh_op_bnr_0')
// (16, 8, 'neigh_op_top_0')
// (16, 9, 'lutff_0/out')
// (16, 10, 'local_g1_0')
// (16, 10, 'lutff_6/in_1')
// (16, 10, 'neigh_op_bot_0')
// (17, 8, 'neigh_op_tnl_0')
// (17, 9, 'neigh_op_lft_0')
// (17, 10, 'neigh_op_bnl_0')

wire n2215;
// (15, 8, 'neigh_op_tnr_1')
// (15, 9, 'neigh_op_rgt_1')
// (15, 10, 'neigh_op_bnr_1')
// (16, 8, 'neigh_op_top_1')
// (16, 9, 'lutff_1/out')
// (16, 10, 'neigh_op_bot_1')
// (17, 8, 'neigh_op_tnl_1')
// (17, 9, 'local_g0_1')
// (17, 9, 'lutff_7/in_0')
// (17, 9, 'neigh_op_lft_1')
// (17, 10, 'neigh_op_bnl_1')

wire n2216;
// (15, 8, 'neigh_op_tnr_2')
// (15, 9, 'neigh_op_rgt_2')
// (15, 10, 'neigh_op_bnr_2')
// (16, 8, 'neigh_op_top_2')
// (16, 9, 'lutff_2/out')
// (16, 10, 'local_g1_2')
// (16, 10, 'lutff_1/in_0')
// (16, 10, 'neigh_op_bot_2')
// (17, 8, 'neigh_op_tnl_2')
// (17, 9, 'neigh_op_lft_2')
// (17, 10, 'neigh_op_bnl_2')

wire n2217;
// (15, 8, 'neigh_op_tnr_3')
// (15, 9, 'neigh_op_rgt_3')
// (15, 10, 'neigh_op_bnr_3')
// (16, 8, 'neigh_op_top_3')
// (16, 9, 'lutff_3/out')
// (16, 10, 'local_g1_3')
// (16, 10, 'lutff_3/in_3')
// (16, 10, 'neigh_op_bot_3')
// (17, 8, 'neigh_op_tnl_3')
// (17, 9, 'neigh_op_lft_3')
// (17, 10, 'neigh_op_bnl_3')

wire n2218;
// (15, 8, 'neigh_op_tnr_5')
// (15, 9, 'neigh_op_rgt_5')
// (15, 10, 'neigh_op_bnr_5')
// (16, 8, 'neigh_op_top_5')
// (16, 9, 'local_g1_5')
// (16, 9, 'lutff_5/out')
// (16, 9, 'lutff_7/in_1')
// (16, 10, 'neigh_op_bot_5')
// (17, 8, 'neigh_op_tnl_5')
// (17, 9, 'neigh_op_lft_5')
// (17, 10, 'neigh_op_bnl_5')

wire n2219;
// (15, 8, 'neigh_op_tnr_6')
// (15, 9, 'neigh_op_rgt_6')
// (15, 10, 'neigh_op_bnr_6')
// (16, 8, 'neigh_op_top_6')
// (16, 9, 'lutff_6/out')
// (16, 10, 'local_g1_6')
// (16, 10, 'lutff_3/in_2')
// (16, 10, 'neigh_op_bot_6')
// (17, 8, 'neigh_op_tnl_6')
// (17, 9, 'neigh_op_lft_6')
// (17, 10, 'neigh_op_bnl_6')

wire n2220;
// (15, 8, 'neigh_op_tnr_7')
// (15, 8, 'sp4_r_v_b_43')
// (15, 9, 'neigh_op_rgt_7')
// (15, 9, 'sp4_r_v_b_30')
// (15, 10, 'neigh_op_bnr_7')
// (15, 10, 'sp4_r_v_b_19')
// (15, 11, 'sp4_r_v_b_6')
// (16, 7, 'sp4_v_t_43')
// (16, 8, 'neigh_op_top_7')
// (16, 8, 'sp4_v_b_43')
// (16, 9, 'lutff_7/out')
// (16, 9, 'sp4_v_b_30')
// (16, 10, 'neigh_op_bot_7')
// (16, 10, 'sp4_v_b_19')
// (16, 11, 'local_g0_6')
// (16, 11, 'lutff_0/in_0')
// (16, 11, 'sp4_v_b_6')
// (17, 8, 'neigh_op_tnl_7')
// (17, 9, 'neigh_op_lft_7')
// (17, 10, 'neigh_op_bnl_7')

reg n2221 = 0;
// (15, 9, 'neigh_op_tnr_0')
// (15, 10, 'neigh_op_rgt_0')
// (15, 10, 'sp4_h_r_5')
// (15, 11, 'neigh_op_bnr_0')
// (16, 9, 'neigh_op_top_0')
// (16, 10, 'lutff_0/out')
// (16, 10, 'sp4_h_r_16')
// (16, 11, 'neigh_op_bot_0')
// (17, 9, 'neigh_op_tnl_0')
// (17, 10, 'neigh_op_lft_0')
// (17, 10, 'sp4_h_r_29')
// (17, 11, 'neigh_op_bnl_0')
// (18, 7, 'sp4_r_v_b_40')
// (18, 8, 'sp4_r_v_b_29')
// (18, 9, 'local_g3_0')
// (18, 9, 'lutff_7/in_0')
// (18, 9, 'sp4_r_v_b_16')
// (18, 10, 'sp4_h_r_40')
// (18, 10, 'sp4_r_v_b_5')
// (19, 6, 'sp4_v_t_40')
// (19, 7, 'sp4_v_b_40')
// (19, 8, 'sp4_v_b_29')
// (19, 9, 'sp4_v_b_16')
// (19, 10, 'sp4_h_l_40')
// (19, 10, 'sp4_v_b_5')

wire n2222;
// (15, 9, 'neigh_op_tnr_1')
// (15, 10, 'neigh_op_rgt_1')
// (15, 11, 'neigh_op_bnr_1')
// (16, 9, 'neigh_op_top_1')
// (16, 10, 'lutff_1/out')
// (16, 11, 'local_g1_1')
// (16, 11, 'lutff_4/in_0')
// (16, 11, 'neigh_op_bot_1')
// (17, 9, 'neigh_op_tnl_1')
// (17, 10, 'neigh_op_lft_1')
// (17, 11, 'neigh_op_bnl_1')

wire n2223;
// (15, 9, 'neigh_op_tnr_2')
// (15, 10, 'neigh_op_rgt_2')
// (15, 11, 'neigh_op_bnr_2')
// (16, 9, 'neigh_op_top_2')
// (16, 10, 'lutff_2/out')
// (16, 11, 'neigh_op_bot_2')
// (17, 9, 'neigh_op_tnl_2')
// (17, 10, 'neigh_op_lft_2')
// (17, 11, 'local_g3_2')
// (17, 11, 'lutff_7/in_0')
// (17, 11, 'neigh_op_bnl_2')

wire n2224;
// (15, 9, 'neigh_op_tnr_3')
// (15, 10, 'neigh_op_rgt_3')
// (15, 11, 'local_g0_3')
// (15, 11, 'lutff_0/in_3')
// (15, 11, 'neigh_op_bnr_3')
// (16, 9, 'neigh_op_top_3')
// (16, 10, 'lutff_3/out')
// (16, 11, 'neigh_op_bot_3')
// (17, 9, 'neigh_op_tnl_3')
// (17, 10, 'neigh_op_lft_3')
// (17, 11, 'neigh_op_bnl_3')

wire n2225;
// (15, 9, 'neigh_op_tnr_4')
// (15, 10, 'neigh_op_rgt_4')
// (15, 11, 'neigh_op_bnr_4')
// (16, 9, 'neigh_op_top_4')
// (16, 10, 'local_g1_4')
// (16, 10, 'lutff_3/in_0')
// (16, 10, 'lutff_4/out')
// (16, 11, 'neigh_op_bot_4')
// (17, 9, 'neigh_op_tnl_4')
// (17, 10, 'neigh_op_lft_4')
// (17, 11, 'neigh_op_bnl_4')

reg n2226 = 0;
// (15, 9, 'neigh_op_tnr_5')
// (15, 10, 'neigh_op_rgt_5')
// (15, 11, 'neigh_op_bnr_5')
// (16, 9, 'neigh_op_top_5')
// (16, 10, 'local_g2_5')
// (16, 10, 'lutff_4/in_1')
// (16, 10, 'lutff_5/out')
// (16, 11, 'neigh_op_bot_5')
// (17, 9, 'neigh_op_tnl_5')
// (17, 10, 'neigh_op_lft_5')
// (17, 11, 'neigh_op_bnl_5')

wire n2227;
// (15, 9, 'neigh_op_tnr_6')
// (15, 10, 'neigh_op_rgt_6')
// (15, 11, 'local_g0_6')
// (15, 11, 'lutff_2/in_0')
// (15, 11, 'neigh_op_bnr_6')
// (16, 9, 'neigh_op_top_6')
// (16, 10, 'lutff_6/out')
// (16, 11, 'neigh_op_bot_6')
// (17, 9, 'neigh_op_tnl_6')
// (17, 10, 'neigh_op_lft_6')
// (17, 11, 'neigh_op_bnl_6')

wire n2228;
// (15, 9, 'neigh_op_tnr_7')
// (15, 10, 'neigh_op_rgt_7')
// (15, 11, 'neigh_op_bnr_7')
// (16, 9, 'neigh_op_top_7')
// (16, 10, 'local_g3_7')
// (16, 10, 'lutff_1/in_3')
// (16, 10, 'lutff_7/out')
// (16, 11, 'neigh_op_bot_7')
// (17, 9, 'neigh_op_tnl_7')
// (17, 10, 'neigh_op_lft_7')
// (17, 11, 'neigh_op_bnl_7')

reg n2229 = 0;
// (15, 9, 'sp4_h_r_10')
// (16, 9, 'local_g1_7')
// (16, 9, 'lutff_2/in_0')
// (16, 9, 'sp4_h_r_23')
// (17, 9, 'sp4_h_r_34')
// (18, 9, 'sp4_h_r_47')
// (19, 8, 'neigh_op_tnr_1')
// (19, 9, 'neigh_op_rgt_1')
// (19, 9, 'sp4_h_l_47')
// (19, 9, 'sp4_h_r_7')
// (19, 10, 'neigh_op_bnr_1')
// (20, 8, 'neigh_op_top_1')
// (20, 9, 'lutff_1/out')
// (20, 9, 'sp4_h_r_18')
// (20, 10, 'neigh_op_bot_1')
// (21, 8, 'neigh_op_tnl_1')
// (21, 9, 'neigh_op_lft_1')
// (21, 9, 'sp4_h_r_31')
// (21, 10, 'neigh_op_bnl_1')
// (22, 9, 'sp4_h_r_42')
// (23, 9, 'sp4_h_l_42')

reg n2230 = 0;
// (15, 10, 'neigh_op_tnr_1')
// (15, 11, 'neigh_op_rgt_1')
// (15, 12, 'neigh_op_bnr_1')
// (16, 10, 'neigh_op_top_1')
// (16, 11, 'lutff_1/out')
// (16, 12, 'neigh_op_bot_1')
// (17, 10, 'local_g2_1')
// (17, 10, 'lutff_5/in_2')
// (17, 10, 'neigh_op_tnl_1')
// (17, 11, 'neigh_op_lft_1')
// (17, 12, 'neigh_op_bnl_1')

reg n2231 = 0;
// (15, 10, 'neigh_op_tnr_2')
// (15, 11, 'neigh_op_rgt_2')
// (15, 12, 'neigh_op_bnr_2')
// (16, 10, 'neigh_op_top_2')
// (16, 11, 'local_g2_2')
// (16, 11, 'lutff_2/out')
// (16, 11, 'lutff_5/in_3')
// (16, 12, 'neigh_op_bot_2')
// (17, 10, 'neigh_op_tnl_2')
// (17, 11, 'neigh_op_lft_2')
// (17, 12, 'neigh_op_bnl_2')

wire n2232;
// (15, 10, 'neigh_op_tnr_3')
// (15, 11, 'neigh_op_rgt_3')
// (15, 12, 'neigh_op_bnr_3')
// (16, 10, 'neigh_op_top_3')
// (16, 11, 'local_g3_3')
// (16, 11, 'lutff_0/in_2')
// (16, 11, 'lutff_3/out')
// (16, 12, 'neigh_op_bot_3')
// (17, 10, 'neigh_op_tnl_3')
// (17, 11, 'neigh_op_lft_3')
// (17, 12, 'neigh_op_bnl_3')

wire n2233;
// (15, 10, 'neigh_op_tnr_4')
// (15, 11, 'local_g2_4')
// (15, 11, 'lutff_1/in_1')
// (15, 11, 'neigh_op_rgt_4')
// (15, 12, 'neigh_op_bnr_4')
// (16, 10, 'neigh_op_top_4')
// (16, 11, 'lutff_4/out')
// (16, 12, 'neigh_op_bot_4')
// (17, 10, 'neigh_op_tnl_4')
// (17, 11, 'neigh_op_lft_4')
// (17, 12, 'neigh_op_bnl_4')

wire n2234;
// (15, 10, 'neigh_op_tnr_5')
// (15, 11, 'neigh_op_rgt_5')
// (15, 12, 'neigh_op_bnr_5')
// (16, 10, 'neigh_op_top_5')
// (16, 11, 'local_g0_5')
// (16, 11, 'lutff_3/in_0')
// (16, 11, 'lutff_5/out')
// (16, 12, 'neigh_op_bot_5')
// (17, 10, 'neigh_op_tnl_5')
// (17, 11, 'neigh_op_lft_5')
// (17, 12, 'neigh_op_bnl_5')

wire n2235;
// (15, 10, 'neigh_op_tnr_6')
// (15, 11, 'neigh_op_rgt_6')
// (15, 12, 'neigh_op_bnr_6')
// (16, 10, 'neigh_op_top_6')
// (16, 11, 'local_g3_6')
// (16, 11, 'lutff_4/in_1')
// (16, 11, 'lutff_6/out')
// (16, 12, 'neigh_op_bot_6')
// (17, 10, 'neigh_op_tnl_6')
// (17, 11, 'neigh_op_lft_6')
// (17, 12, 'neigh_op_bnl_6')

reg n2236 = 0;
// (15, 10, 'neigh_op_tnr_7')
// (15, 11, 'neigh_op_rgt_7')
// (15, 12, 'neigh_op_bnr_7')
// (16, 10, 'neigh_op_top_7')
// (16, 11, 'local_g3_7')
// (16, 11, 'lutff_6/in_2')
// (16, 11, 'lutff_7/out')
// (16, 12, 'neigh_op_bot_7')
// (17, 10, 'neigh_op_tnl_7')
// (17, 11, 'neigh_op_lft_7')
// (17, 12, 'neigh_op_bnl_7')

wire n2237;
// (15, 11, 'local_g2_6')
// (15, 11, 'local_g3_6')
// (15, 11, 'lutff_0/in_1')
// (15, 11, 'lutff_2/in_2')
// (15, 11, 'neigh_op_tnr_6')
// (15, 12, 'neigh_op_rgt_6')
// (15, 13, 'local_g1_6')
// (15, 13, 'lutff_1/in_2')
// (15, 13, 'neigh_op_bnr_6')
// (16, 11, 'neigh_op_top_6')
// (16, 12, 'local_g2_6')
// (16, 12, 'lutff_2/in_2')
// (16, 12, 'lutff_4/in_0')
// (16, 12, 'lutff_6/out')
// (16, 13, 'neigh_op_bot_6')
// (17, 11, 'neigh_op_tnl_6')
// (17, 12, 'local_g0_6')
// (17, 12, 'lutff_5/in_1')
// (17, 12, 'neigh_op_lft_6')
// (17, 13, 'neigh_op_bnl_6')

wire n2238;
// (15, 11, 'local_g3_0')
// (15, 11, 'lutff_1/in_2')
// (15, 11, 'lutff_3/in_2')
// (15, 11, 'lutff_6/in_3')
// (15, 11, 'neigh_op_tnr_0')
// (15, 12, 'local_g2_0')
// (15, 12, 'lutff_1/in_3')
// (15, 12, 'lutff_5/in_1')
// (15, 12, 'lutff_7/in_3')
// (15, 12, 'neigh_op_rgt_0')
// (15, 13, 'neigh_op_bnr_0')
// (16, 11, 'neigh_op_top_0')
// (16, 12, 'local_g1_0')
// (16, 12, 'lutff_0/out')
// (16, 12, 'lutff_3/in_0')
// (16, 12, 'lutff_4/in_1')
// (16, 12, 'lutff_5/in_0')
// (16, 13, 'local_g1_0')
// (16, 13, 'lutff_0/in_3')
// (16, 13, 'neigh_op_bot_0')
// (17, 11, 'neigh_op_tnl_0')
// (17, 12, 'neigh_op_lft_0')
// (17, 13, 'neigh_op_bnl_0')

wire n2239;
// (15, 11, 'local_g3_2')
// (15, 11, 'lutff_1/in_0')
// (15, 11, 'neigh_op_tnr_2')
// (15, 12, 'neigh_op_rgt_2')
// (15, 13, 'neigh_op_bnr_2')
// (16, 11, 'local_g1_2')
// (16, 11, 'lutff_0/in_3')
// (16, 11, 'neigh_op_top_2')
// (16, 12, 'local_g3_2')
// (16, 12, 'lutff_2/out')
// (16, 12, 'lutff_3/in_2')
// (16, 13, 'neigh_op_bot_2')
// (17, 11, 'neigh_op_tnl_2')
// (17, 12, 'local_g0_2')
// (17, 12, 'lutff_4/in_0')
// (17, 12, 'neigh_op_lft_2')
// (17, 13, 'neigh_op_bnl_2')

reg n2240 = 0;
// (15, 11, 'neigh_op_tnr_1')
// (15, 12, 'neigh_op_rgt_1')
// (15, 13, 'neigh_op_bnr_1')
// (16, 11, 'neigh_op_top_1')
// (16, 12, 'lutff_1/out')
// (16, 13, 'neigh_op_bot_1')
// (17, 11, 'local_g2_1')
// (17, 11, 'lutff_6/in_1')
// (17, 11, 'neigh_op_tnl_1')
// (17, 12, 'neigh_op_lft_1')
// (17, 13, 'neigh_op_bnl_1')

wire n2241;
// (15, 11, 'neigh_op_tnr_3')
// (15, 12, 'local_g2_3')
// (15, 12, 'lutff_0/in_3')
// (15, 12, 'neigh_op_rgt_3')
// (15, 13, 'neigh_op_bnr_3')
// (16, 11, 'neigh_op_top_3')
// (16, 12, 'lutff_3/out')
// (16, 13, 'neigh_op_bot_3')
// (17, 11, 'neigh_op_tnl_3')
// (17, 12, 'neigh_op_lft_3')
// (17, 13, 'neigh_op_bnl_3')

wire n2242;
// (15, 11, 'neigh_op_tnr_4')
// (15, 12, 'neigh_op_rgt_4')
// (15, 13, 'local_g1_4')
// (15, 13, 'lutff_5/in_0')
// (15, 13, 'neigh_op_bnr_4')
// (16, 11, 'neigh_op_top_4')
// (16, 12, 'lutff_4/out')
// (16, 13, 'neigh_op_bot_4')
// (17, 11, 'neigh_op_tnl_4')
// (17, 12, 'neigh_op_lft_4')
// (17, 13, 'neigh_op_bnl_4')

wire n2243;
// (15, 11, 'neigh_op_tnr_5')
// (15, 12, 'local_g2_5')
// (15, 12, 'lutff_4/in_3')
// (15, 12, 'neigh_op_rgt_5')
// (15, 13, 'neigh_op_bnr_5')
// (16, 11, 'neigh_op_top_5')
// (16, 12, 'lutff_5/out')
// (16, 13, 'neigh_op_bot_5')
// (17, 11, 'neigh_op_tnl_5')
// (17, 12, 'neigh_op_lft_5')
// (17, 13, 'neigh_op_bnl_5')

reg n2244 = 0;
// (15, 11, 'neigh_op_tnr_7')
// (15, 12, 'neigh_op_rgt_7')
// (15, 13, 'neigh_op_bnr_7')
// (16, 11, 'neigh_op_top_7')
// (16, 12, 'lutff_7/out')
// (16, 13, 'neigh_op_bot_7')
// (17, 11, 'local_g2_7')
// (17, 11, 'lutff_3/in_0')
// (17, 11, 'neigh_op_tnl_7')
// (17, 12, 'neigh_op_lft_7')
// (17, 13, 'neigh_op_bnl_7')

wire n2245;
// (15, 11, 'sp4_r_v_b_45')
// (15, 12, 'sp4_r_v_b_32')
// (15, 13, 'neigh_op_tnr_4')
// (15, 13, 'sp4_r_v_b_21')
// (15, 14, 'neigh_op_rgt_4')
// (15, 14, 'sp4_r_v_b_8')
// (15, 15, 'neigh_op_bnr_4')
// (16, 10, 'sp4_v_t_45')
// (16, 11, 'sp4_v_b_45')
// (16, 12, 'local_g2_0')
// (16, 12, 'lutff_0/in_2')
// (16, 12, 'lutff_6/in_2')
// (16, 12, 'sp4_v_b_32')
// (16, 13, 'neigh_op_top_4')
// (16, 13, 'sp4_v_b_21')
// (16, 14, 'lutff_4/out')
// (16, 14, 'sp4_v_b_8')
// (16, 15, 'neigh_op_bot_4')
// (17, 13, 'neigh_op_tnl_4')
// (17, 14, 'neigh_op_lft_4')
// (17, 15, 'neigh_op_bnl_4')

wire n2246;
// (15, 12, 'neigh_op_tnr_0')
// (15, 13, 'neigh_op_rgt_0')
// (15, 14, 'local_g1_0')
// (15, 14, 'lutff_0/in_3')
// (15, 14, 'neigh_op_bnr_0')
// (16, 12, 'neigh_op_top_0')
// (16, 13, 'lutff_0/out')
// (16, 14, 'neigh_op_bot_0')
// (17, 12, 'neigh_op_tnl_0')
// (17, 13, 'neigh_op_lft_0')
// (17, 14, 'neigh_op_bnl_0')

wire n2247;
// (15, 12, 'neigh_op_tnr_1')
// (15, 13, 'neigh_op_rgt_1')
// (15, 14, 'neigh_op_bnr_1')
// (16, 12, 'local_g0_1')
// (16, 12, 'lutff_0/in_1')
// (16, 12, 'neigh_op_top_1')
// (16, 13, 'lutff_1/out')
// (16, 14, 'neigh_op_bot_1')
// (17, 12, 'neigh_op_tnl_1')
// (17, 13, 'neigh_op_lft_1')
// (17, 14, 'neigh_op_bnl_1')

wire n2248;
// (15, 12, 'sp4_h_r_0')
// (16, 12, 'sp4_h_r_13')
// (17, 12, 'local_g2_0')
// (17, 12, 'lutff_0/in_0')
// (17, 12, 'sp4_h_r_24')
// (18, 9, 'sp4_r_v_b_42')
// (18, 10, 'neigh_op_tnr_1')
// (18, 10, 'sp4_r_v_b_31')
// (18, 11, 'neigh_op_rgt_1')
// (18, 11, 'sp4_r_v_b_18')
// (18, 12, 'neigh_op_bnr_1')
// (18, 12, 'sp4_h_r_37')
// (18, 12, 'sp4_r_v_b_7')
// (19, 8, 'sp4_v_t_42')
// (19, 9, 'sp4_v_b_42')
// (19, 10, 'neigh_op_top_1')
// (19, 10, 'sp4_v_b_31')
// (19, 11, 'ram/RDATA_14')
// (19, 11, 'sp4_v_b_18')
// (19, 12, 'neigh_op_bot_1')
// (19, 12, 'sp4_h_l_37')
// (19, 12, 'sp4_v_b_7')
// (20, 10, 'neigh_op_tnl_1')
// (20, 11, 'neigh_op_lft_1')
// (20, 12, 'neigh_op_bnl_1')

reg n2249 = 0;
// (15, 12, 'sp4_r_v_b_41')
// (15, 13, 'sp4_r_v_b_28')
// (15, 14, 'neigh_op_tnr_2')
// (15, 14, 'sp4_r_v_b_17')
// (15, 15, 'neigh_op_rgt_2')
// (15, 15, 'sp4_r_v_b_4')
// (15, 16, 'neigh_op_bnr_2')
// (16, 11, 'sp4_h_r_4')
// (16, 11, 'sp4_v_t_41')
// (16, 12, 'sp4_v_b_41')
// (16, 13, 'sp4_v_b_28')
// (16, 14, 'neigh_op_top_2')
// (16, 14, 'sp4_v_b_17')
// (16, 15, 'lutff_2/out')
// (16, 15, 'sp4_v_b_4')
// (16, 16, 'neigh_op_bot_2')
// (17, 11, 'sp4_h_r_17')
// (17, 14, 'neigh_op_tnl_2')
// (17, 15, 'neigh_op_lft_2')
// (17, 16, 'neigh_op_bnl_2')
// (18, 11, 'sp4_h_r_28')
// (19, 8, 'sp4_r_v_b_41')
// (19, 9, 'sp4_r_v_b_28')
// (19, 10, 'local_g3_1')
// (19, 10, 'ram/WDATA_2')
// (19, 10, 'sp4_r_v_b_17')
// (19, 11, 'sp4_h_r_41')
// (19, 11, 'sp4_r_v_b_4')
// (20, 7, 'sp4_v_t_41')
// (20, 8, 'sp4_v_b_41')
// (20, 9, 'sp4_v_b_28')
// (20, 10, 'sp4_v_b_17')
// (20, 11, 'sp4_h_l_41')
// (20, 11, 'sp4_v_b_4')

wire n2250;
// (15, 12, 'sp4_r_v_b_43')
// (15, 13, 'sp4_r_v_b_30')
// (15, 14, 'sp4_r_v_b_19')
// (15, 15, 'sp4_r_v_b_6')
// (15, 17, 'sp4_h_r_11')
// (16, 11, 'sp4_h_r_0')
// (16, 11, 'sp4_v_t_43')
// (16, 12, 'sp4_v_b_43')
// (16, 13, 'sp4_v_b_30')
// (16, 14, 'local_g1_3')
// (16, 14, 'lutff_2/in_2')
// (16, 14, 'sp4_v_b_19')
// (16, 15, 'sp4_v_b_6')
// (16, 17, 'local_g1_6')
// (16, 17, 'lutff_1/in_0')
// (16, 17, 'sp4_h_r_22')
// (17, 11, 'sp4_h_r_13')
// (17, 17, 'sp4_h_r_35')
// (18, 11, 'sp4_h_r_24')
// (18, 14, 'sp4_r_v_b_43')
// (18, 15, 'sp4_r_v_b_30')
// (18, 16, 'sp4_r_v_b_19')
// (18, 17, 'sp4_h_r_46')
// (18, 17, 'sp4_r_v_b_6')
// (19, 11, 'sp4_h_r_37')
// (19, 13, 'sp4_h_r_6')
// (19, 13, 'sp4_v_t_43')
// (19, 14, 'sp4_v_b_43')
// (19, 15, 'sp4_v_b_30')
// (19, 16, 'sp4_v_b_19')
// (19, 17, 'sp4_h_l_46')
// (19, 17, 'sp4_v_b_6')
// (20, 11, 'sp4_h_l_37')
// (20, 11, 'sp4_h_r_0')
// (20, 13, 'sp4_h_r_19')
// (21, 10, 'neigh_op_tnr_4')
// (21, 11, 'neigh_op_rgt_4')
// (21, 11, 'sp4_h_r_13')
// (21, 12, 'neigh_op_bnr_4')
// (21, 13, 'sp4_h_r_30')
// (22, 10, 'neigh_op_top_4')
// (22, 10, 'sp4_r_v_b_36')
// (22, 11, 'lutff_4/out')
// (22, 11, 'sp4_h_r_24')
// (22, 11, 'sp4_r_v_b_25')
// (22, 12, 'neigh_op_bot_4')
// (22, 12, 'sp4_r_v_b_12')
// (22, 13, 'sp4_h_r_43')
// (22, 13, 'sp4_r_v_b_1')
// (23, 9, 'sp4_v_t_36')
// (23, 10, 'neigh_op_tnl_4')
// (23, 10, 'sp4_v_b_36')
// (23, 11, 'neigh_op_lft_4')
// (23, 11, 'sp4_h_r_37')
// (23, 11, 'sp4_v_b_25')
// (23, 12, 'neigh_op_bnl_4')
// (23, 12, 'sp4_v_b_12')
// (23, 13, 'sp4_h_l_43')
// (23, 13, 'sp4_v_b_1')
// (24, 11, 'sp4_h_l_37')

wire n2251;
// (15, 13, 'local_g2_5')
// (15, 13, 'lutff_4/in_3')
// (15, 13, 'neigh_op_tnr_5')
// (15, 14, 'neigh_op_rgt_5')
// (15, 14, 'sp4_r_v_b_42')
// (15, 15, 'neigh_op_bnr_5')
// (15, 15, 'sp4_r_v_b_31')
// (15, 16, 'local_g3_2')
// (15, 16, 'lutff_6/in_1')
// (15, 16, 'sp4_r_v_b_18')
// (15, 17, 'sp4_r_v_b_7')
// (16, 13, 'local_g0_5')
// (16, 13, 'lutff_1/in_2')
// (16, 13, 'lutff_7/in_0')
// (16, 13, 'neigh_op_top_5')
// (16, 13, 'sp4_v_t_42')
// (16, 14, 'lutff_5/out')
// (16, 14, 'sp4_v_b_42')
// (16, 15, 'neigh_op_bot_5')
// (16, 15, 'sp4_v_b_31')
// (16, 16, 'sp4_v_b_18')
// (16, 17, 'sp4_v_b_7')
// (17, 13, 'neigh_op_tnl_5')
// (17, 14, 'neigh_op_lft_5')
// (17, 15, 'neigh_op_bnl_5')

wire n2252;
// (15, 13, 'neigh_op_tnr_0')
// (15, 14, 'local_g2_0')
// (15, 14, 'lutff_5/in_1')
// (15, 14, 'neigh_op_rgt_0')
// (15, 15, 'neigh_op_bnr_0')
// (16, 13, 'neigh_op_top_0')
// (16, 14, 'local_g3_0')
// (16, 14, 'lutff_0/out')
// (16, 14, 'lutff_5/in_0')
// (16, 15, 'neigh_op_bot_0')
// (17, 13, 'neigh_op_tnl_0')
// (17, 14, 'neigh_op_lft_0')
// (17, 15, 'neigh_op_bnl_0')

wire n2253;
// (15, 13, 'neigh_op_tnr_1')
// (15, 14, 'neigh_op_rgt_1')
// (15, 14, 'sp4_h_r_1')
// (15, 14, 'sp4_h_r_7')
// (15, 15, 'neigh_op_bnr_1')
// (16, 13, 'neigh_op_top_1')
// (16, 14, 'local_g0_4')
// (16, 14, 'lutff_1/out')
// (16, 14, 'lutff_global/s_r')
// (16, 14, 'sp4_h_r_12')
// (16, 14, 'sp4_h_r_18')
// (16, 15, 'neigh_op_bot_1')
// (17, 13, 'neigh_op_tnl_1')
// (17, 14, 'neigh_op_lft_1')
// (17, 14, 'sp4_h_r_25')
// (17, 14, 'sp4_h_r_31')
// (17, 15, 'neigh_op_bnl_1')
// (18, 14, 'sp4_h_r_36')
// (18, 14, 'sp4_h_r_42')
// (19, 14, 'sp4_h_l_36')
// (19, 14, 'sp4_h_l_42')
// (19, 14, 'sp4_h_r_10')
// (20, 14, 'sp4_h_r_23')
// (21, 14, 'sp4_h_r_34')
// (22, 14, 'sp4_h_r_47')
// (23, 14, 'sp4_h_l_47')

wire n2254;
// (15, 13, 'neigh_op_tnr_6')
// (15, 14, 'neigh_op_rgt_6')
// (15, 15, 'neigh_op_bnr_6')
// (16, 13, 'local_g0_6')
// (16, 13, 'lutff_1/in_1')
// (16, 13, 'lutff_7/in_1')
// (16, 13, 'neigh_op_top_6')
// (16, 14, 'lutff_6/out')
// (16, 15, 'neigh_op_bot_6')
// (17, 13, 'neigh_op_tnl_6')
// (17, 14, 'neigh_op_lft_6')
// (17, 15, 'neigh_op_bnl_6')

reg n2255 = 0;
// (15, 13, 'sp4_h_r_0')
// (16, 12, 'neigh_op_tnr_4')
// (16, 13, 'neigh_op_rgt_4')
// (16, 13, 'sp4_h_r_13')
// (16, 14, 'neigh_op_bnr_4')
// (17, 12, 'neigh_op_top_4')
// (17, 13, 'local_g2_4')
// (17, 13, 'lutff_4/in_2')
// (17, 13, 'lutff_4/out')
// (17, 13, 'sp4_h_r_24')
// (17, 14, 'neigh_op_bot_4')
// (18, 10, 'sp4_r_v_b_37')
// (18, 11, 'sp4_r_v_b_24')
// (18, 12, 'neigh_op_tnl_4')
// (18, 12, 'sp4_r_v_b_13')
// (18, 13, 'neigh_op_lft_4')
// (18, 13, 'sp4_h_r_37')
// (18, 13, 'sp4_r_v_b_0')
// (18, 14, 'neigh_op_bnl_4')
// (18, 14, 'sp4_r_v_b_40')
// (18, 15, 'sp4_r_v_b_29')
// (18, 16, 'sp4_r_v_b_16')
// (18, 17, 'sp4_r_v_b_5')
// (19, 9, 'sp4_v_t_37')
// (19, 10, 'local_g2_5')
// (19, 10, 'ram/WADDR_4')
// (19, 10, 'sp4_v_b_37')
// (19, 11, 'sp4_v_b_24')
// (19, 12, 'local_g0_5')
// (19, 12, 'ram/WADDR_4')
// (19, 12, 'sp4_v_b_13')
// (19, 13, 'sp4_h_l_37')
// (19, 13, 'sp4_v_b_0')
// (19, 13, 'sp4_v_t_40')
// (19, 14, 'local_g3_0')
// (19, 14, 'ram/WADDR_4')
// (19, 14, 'sp4_v_b_40')
// (19, 15, 'sp4_v_b_29')
// (19, 16, 'sp4_v_b_16')
// (19, 17, 'sp4_v_b_5')

reg n2256 = 0;
// (15, 13, 'sp4_h_r_2')
// (16, 12, 'neigh_op_tnr_5')
// (16, 13, 'neigh_op_rgt_5')
// (16, 13, 'sp4_h_r_15')
// (16, 14, 'neigh_op_bnr_5')
// (17, 12, 'neigh_op_top_5')
// (17, 13, 'local_g1_5')
// (17, 13, 'lutff_5/in_1')
// (17, 13, 'lutff_5/out')
// (17, 13, 'sp4_h_r_26')
// (17, 14, 'neigh_op_bot_5')
// (18, 10, 'sp4_r_v_b_39')
// (18, 11, 'sp4_r_v_b_26')
// (18, 12, 'neigh_op_tnl_5')
// (18, 12, 'sp4_r_v_b_15')
// (18, 13, 'neigh_op_lft_5')
// (18, 13, 'sp4_h_r_39')
// (18, 13, 'sp4_r_v_b_2')
// (18, 14, 'neigh_op_bnl_5')
// (18, 14, 'sp4_r_v_b_39')
// (18, 15, 'sp4_r_v_b_26')
// (18, 16, 'sp4_r_v_b_15')
// (18, 17, 'sp4_r_v_b_2')
// (19, 9, 'sp4_v_t_39')
// (19, 10, 'local_g3_7')
// (19, 10, 'ram/WADDR_5')
// (19, 10, 'sp4_v_b_39')
// (19, 11, 'sp4_v_b_26')
// (19, 12, 'local_g1_7')
// (19, 12, 'ram/WADDR_5')
// (19, 12, 'sp4_v_b_15')
// (19, 13, 'sp4_h_l_39')
// (19, 13, 'sp4_v_b_2')
// (19, 13, 'sp4_v_t_39')
// (19, 14, 'local_g3_7')
// (19, 14, 'ram/WADDR_5')
// (19, 14, 'sp4_v_b_39')
// (19, 15, 'sp4_v_b_26')
// (19, 16, 'sp4_v_b_15')
// (19, 17, 'sp4_v_b_2')

reg n2257 = 0;
// (15, 13, 'sp4_h_r_6')
// (16, 12, 'neigh_op_tnr_7')
// (16, 13, 'neigh_op_rgt_7')
// (16, 13, 'sp4_h_r_19')
// (16, 14, 'neigh_op_bnr_7')
// (17, 11, 'sp4_r_v_b_39')
// (17, 12, 'neigh_op_top_7')
// (17, 12, 'sp4_r_v_b_26')
// (17, 13, 'local_g1_7')
// (17, 13, 'lutff_0/in_2')
// (17, 13, 'lutff_1/in_3')
// (17, 13, 'lutff_7/in_1')
// (17, 13, 'lutff_7/out')
// (17, 13, 'sp4_h_r_30')
// (17, 13, 'sp4_r_v_b_15')
// (17, 14, 'neigh_op_bot_7')
// (17, 14, 'sp4_r_v_b_2')
// (18, 10, 'sp4_h_r_7')
// (18, 10, 'sp4_r_v_b_43')
// (18, 10, 'sp4_v_t_39')
// (18, 11, 'sp4_r_v_b_30')
// (18, 11, 'sp4_v_b_39')
// (18, 12, 'neigh_op_tnl_7')
// (18, 12, 'sp4_r_v_b_19')
// (18, 12, 'sp4_v_b_26')
// (18, 13, 'neigh_op_lft_7')
// (18, 13, 'sp4_h_r_43')
// (18, 13, 'sp4_r_v_b_6')
// (18, 13, 'sp4_v_b_15')
// (18, 14, 'neigh_op_bnl_7')
// (18, 14, 'sp4_h_r_2')
// (18, 14, 'sp4_v_b_2')
// (19, 9, 'sp4_v_t_43')
// (19, 10, 'local_g1_2')
// (19, 10, 'ram/WADDR_0')
// (19, 10, 'sp4_h_r_18')
// (19, 10, 'sp4_v_b_43')
// (19, 11, 'sp4_v_b_30')
// (19, 12, 'local_g0_3')
// (19, 12, 'ram/WADDR_0')
// (19, 12, 'sp4_v_b_19')
// (19, 13, 'sp4_h_l_43')
// (19, 13, 'sp4_v_b_6')
// (19, 14, 'local_g0_7')
// (19, 14, 'ram/WADDR_0')
// (19, 14, 'sp4_h_r_15')
// (20, 10, 'sp4_h_r_31')
// (20, 14, 'sp4_h_r_26')
// (21, 10, 'sp4_h_r_42')
// (21, 14, 'sp4_h_r_39')
// (22, 10, 'sp4_h_l_42')
// (22, 14, 'sp4_h_l_39')

reg n2258 = 0;
// (15, 14, 'neigh_op_tnr_0')
// (15, 15, 'neigh_op_rgt_0')
// (15, 16, 'neigh_op_bnr_0')
// (16, 14, 'neigh_op_top_0')
// (16, 15, 'lutff_0/out')
// (16, 15, 'sp4_h_r_0')
// (16, 16, 'neigh_op_bot_0')
// (17, 14, 'neigh_op_tnl_0')
// (17, 15, 'neigh_op_lft_0')
// (17, 15, 'sp4_h_r_13')
// (17, 16, 'neigh_op_bnl_0')
// (18, 15, 'sp4_h_r_24')
// (19, 12, 'sp4_r_v_b_43')
// (19, 13, 'sp4_r_v_b_30')
// (19, 14, 'local_g3_3')
// (19, 14, 'ram/WDATA_6')
// (19, 14, 'sp4_r_v_b_19')
// (19, 15, 'sp4_h_r_37')
// (19, 15, 'sp4_r_v_b_6')
// (20, 11, 'sp4_v_t_43')
// (20, 12, 'sp4_v_b_43')
// (20, 13, 'sp4_v_b_30')
// (20, 14, 'sp4_v_b_19')
// (20, 15, 'sp4_h_l_37')
// (20, 15, 'sp4_v_b_6')

reg n2259 = 0;
// (15, 14, 'neigh_op_tnr_1')
// (15, 15, 'neigh_op_rgt_1')
// (15, 15, 'sp4_h_r_7')
// (15, 16, 'neigh_op_bnr_1')
// (16, 14, 'neigh_op_top_1')
// (16, 15, 'lutff_1/out')
// (16, 15, 'sp4_h_r_18')
// (16, 16, 'neigh_op_bot_1')
// (17, 14, 'neigh_op_tnl_1')
// (17, 15, 'neigh_op_lft_1')
// (17, 15, 'sp4_h_r_31')
// (17, 16, 'neigh_op_bnl_1')
// (18, 12, 'sp4_r_v_b_42')
// (18, 13, 'sp4_r_v_b_31')
// (18, 14, 'sp4_r_v_b_18')
// (18, 15, 'sp4_h_r_42')
// (18, 15, 'sp4_r_v_b_7')
// (19, 11, 'sp4_v_t_42')
// (19, 12, 'sp4_v_b_42')
// (19, 13, 'sp4_v_b_31')
// (19, 14, 'local_g0_2')
// (19, 14, 'ram/WDATA_0')
// (19, 14, 'sp4_v_b_18')
// (19, 15, 'sp4_h_l_42')
// (19, 15, 'sp4_v_b_7')

reg n2260 = 0;
// (15, 14, 'neigh_op_tnr_3')
// (15, 15, 'neigh_op_rgt_3')
// (15, 16, 'neigh_op_bnr_3')
// (16, 14, 'neigh_op_top_3')
// (16, 15, 'lutff_3/out')
// (16, 15, 'sp4_r_v_b_39')
// (16, 16, 'neigh_op_bot_3')
// (16, 16, 'sp4_r_v_b_26')
// (16, 17, 'sp4_r_v_b_15')
// (16, 18, 'sp4_r_v_b_2')
// (17, 14, 'neigh_op_tnl_3')
// (17, 14, 'sp4_h_r_2')
// (17, 14, 'sp4_v_t_39')
// (17, 15, 'neigh_op_lft_3')
// (17, 15, 'sp4_v_b_39')
// (17, 16, 'neigh_op_bnl_3')
// (17, 16, 'sp4_v_b_26')
// (17, 17, 'sp4_v_b_15')
// (17, 18, 'sp4_v_b_2')
// (18, 14, 'sp4_h_r_15')
// (19, 14, 'local_g3_2')
// (19, 14, 'ram/WDATA_3')
// (19, 14, 'sp4_h_r_26')
// (20, 14, 'sp4_h_r_39')
// (21, 14, 'sp4_h_l_39')

reg n2261 = 0;
// (15, 14, 'neigh_op_tnr_4')
// (15, 15, 'neigh_op_rgt_4')
// (15, 15, 'sp4_r_v_b_40')
// (15, 16, 'neigh_op_bnr_4')
// (15, 16, 'sp4_r_v_b_29')
// (15, 17, 'sp4_r_v_b_16')
// (15, 18, 'sp4_r_v_b_5')
// (16, 14, 'neigh_op_top_4')
// (16, 14, 'sp4_h_r_5')
// (16, 14, 'sp4_v_t_40')
// (16, 15, 'lutff_4/out')
// (16, 15, 'sp4_v_b_40')
// (16, 16, 'neigh_op_bot_4')
// (16, 16, 'sp4_v_b_29')
// (16, 17, 'sp4_v_b_16')
// (16, 18, 'sp4_v_b_5')
// (17, 14, 'neigh_op_tnl_4')
// (17, 14, 'sp4_h_r_16')
// (17, 15, 'neigh_op_lft_4')
// (17, 16, 'neigh_op_bnl_4')
// (18, 14, 'sp4_h_r_29')
// (19, 14, 'local_g2_0')
// (19, 14, 'ram/WDATA_4')
// (19, 14, 'sp4_h_r_40')
// (20, 14, 'sp4_h_l_40')

reg n2262 = 0;
// (15, 14, 'neigh_op_tnr_5')
// (15, 15, 'neigh_op_rgt_5')
// (15, 16, 'neigh_op_bnr_5')
// (16, 14, 'neigh_op_top_5')
// (16, 15, 'lutff_5/out')
// (16, 15, 'sp4_r_v_b_43')
// (16, 16, 'neigh_op_bot_5')
// (16, 16, 'sp4_r_v_b_30')
// (16, 17, 'sp4_r_v_b_19')
// (16, 18, 'sp4_r_v_b_6')
// (17, 14, 'neigh_op_tnl_5')
// (17, 14, 'sp4_h_r_6')
// (17, 14, 'sp4_v_t_43')
// (17, 15, 'neigh_op_lft_5')
// (17, 15, 'sp4_v_b_43')
// (17, 16, 'neigh_op_bnl_5')
// (17, 16, 'sp4_v_b_30')
// (17, 17, 'sp4_v_b_19')
// (17, 18, 'sp4_v_b_6')
// (18, 14, 'sp4_h_r_19')
// (19, 14, 'local_g3_6')
// (19, 14, 'ram/WDATA_1')
// (19, 14, 'sp4_h_r_30')
// (20, 14, 'sp4_h_r_43')
// (21, 14, 'sp4_h_l_43')

reg n2263 = 0;
// (15, 14, 'neigh_op_tnr_6')
// (15, 15, 'neigh_op_rgt_6')
// (15, 16, 'neigh_op_bnr_6')
// (16, 14, 'neigh_op_top_6')
// (16, 15, 'lutff_6/out')
// (16, 15, 'sp4_r_v_b_45')
// (16, 16, 'neigh_op_bot_6')
// (16, 16, 'sp4_r_v_b_32')
// (16, 17, 'sp4_r_v_b_21')
// (16, 18, 'sp4_r_v_b_8')
// (17, 14, 'neigh_op_tnl_6')
// (17, 14, 'sp4_h_r_1')
// (17, 14, 'sp4_v_t_45')
// (17, 15, 'neigh_op_lft_6')
// (17, 15, 'sp4_v_b_45')
// (17, 16, 'neigh_op_bnl_6')
// (17, 16, 'sp4_v_b_32')
// (17, 17, 'sp4_v_b_21')
// (17, 18, 'sp4_v_b_8')
// (18, 14, 'sp4_h_r_12')
// (19, 14, 'local_g3_1')
// (19, 14, 'ram/WDATA_2')
// (19, 14, 'sp4_h_r_25')
// (20, 14, 'sp4_h_r_36')
// (21, 14, 'sp4_h_l_36')

reg n2264 = 0;
// (15, 14, 'neigh_op_tnr_7')
// (15, 15, 'neigh_op_rgt_7')
// (15, 15, 'sp4_h_r_3')
// (15, 16, 'neigh_op_bnr_7')
// (16, 14, 'neigh_op_top_7')
// (16, 15, 'lutff_7/out')
// (16, 15, 'sp4_h_r_14')
// (16, 16, 'neigh_op_bot_7')
// (17, 14, 'neigh_op_tnl_7')
// (17, 15, 'neigh_op_lft_7')
// (17, 15, 'sp4_h_r_27')
// (17, 16, 'neigh_op_bnl_7')
// (18, 8, 'sp4_r_v_b_43')
// (18, 9, 'sp4_r_v_b_30')
// (18, 10, 'sp4_r_v_b_19')
// (18, 11, 'sp4_r_v_b_6')
// (18, 12, 'sp4_r_v_b_38')
// (18, 13, 'sp4_r_v_b_27')
// (18, 14, 'sp4_r_v_b_14')
// (18, 15, 'sp4_h_r_38')
// (18, 15, 'sp4_r_v_b_3')
// (19, 7, 'sp4_v_t_43')
// (19, 8, 'sp4_v_b_43')
// (19, 9, 'sp4_v_b_30')
// (19, 10, 'local_g1_3')
// (19, 10, 'ram/WDATA_0')
// (19, 10, 'sp4_v_b_19')
// (19, 11, 'sp4_v_b_6')
// (19, 11, 'sp4_v_t_38')
// (19, 12, 'sp4_v_b_38')
// (19, 13, 'sp4_v_b_27')
// (19, 14, 'sp4_v_b_14')
// (19, 15, 'sp4_h_l_38')
// (19, 15, 'sp4_v_b_3')

reg n2265 = 0;
// (15, 14, 'sp4_h_r_0')
// (16, 13, 'neigh_op_tnr_4')
// (16, 14, 'neigh_op_rgt_4')
// (16, 14, 'sp4_h_r_13')
// (16, 15, 'neigh_op_bnr_4')
// (17, 13, 'neigh_op_top_4')
// (17, 14, 'local_g3_4')
// (17, 14, 'lutff_4/in_1')
// (17, 14, 'lutff_4/out')
// (17, 14, 'sp4_h_r_24')
// (17, 15, 'neigh_op_bot_4')
// (18, 7, 'sp4_r_v_b_45')
// (18, 8, 'sp4_r_v_b_32')
// (18, 9, 'sp4_r_v_b_21')
// (18, 10, 'sp4_r_v_b_8')
// (18, 11, 'sp4_r_v_b_37')
// (18, 12, 'sp4_r_v_b_24')
// (18, 13, 'neigh_op_tnl_4')
// (18, 13, 'sp4_r_v_b_13')
// (18, 14, 'neigh_op_lft_4')
// (18, 14, 'sp4_h_r_37')
// (18, 14, 'sp4_r_v_b_0')
// (18, 15, 'neigh_op_bnl_4')
// (19, 6, 'sp4_v_t_45')
// (19, 7, 'sp4_v_b_45')
// (19, 8, 'sp4_v_b_32')
// (19, 9, 'local_g0_5')
// (19, 9, 'ram/RADDR_4')
// (19, 9, 'sp4_v_b_21')
// (19, 10, 'sp4_v_b_8')
// (19, 10, 'sp4_v_t_37')
// (19, 11, 'local_g2_5')
// (19, 11, 'ram/RADDR_4')
// (19, 11, 'sp4_v_b_37')
// (19, 12, 'sp4_v_b_24')
// (19, 13, 'local_g0_5')
// (19, 13, 'ram/RADDR_4')
// (19, 13, 'sp4_v_b_13')
// (19, 14, 'sp4_h_l_37')
// (19, 14, 'sp4_v_b_0')

reg n2266 = 0;
// (15, 14, 'sp4_h_r_10')
// (16, 13, 'neigh_op_tnr_1')
// (16, 14, 'neigh_op_rgt_1')
// (16, 14, 'sp4_h_r_23')
// (16, 14, 'sp4_h_r_7')
// (16, 15, 'neigh_op_bnr_1')
// (17, 13, 'neigh_op_top_1')
// (17, 14, 'local_g1_1')
// (17, 14, 'lutff_1/in_1')
// (17, 14, 'lutff_1/out')
// (17, 14, 'sp4_h_r_18')
// (17, 14, 'sp4_h_r_34')
// (17, 15, 'neigh_op_bot_1')
// (18, 7, 'sp4_r_v_b_42')
// (18, 8, 'sp4_r_v_b_31')
// (18, 9, 'sp4_r_v_b_18')
// (18, 10, 'sp4_r_v_b_7')
// (18, 11, 'sp4_r_v_b_41')
// (18, 12, 'sp4_r_v_b_28')
// (18, 13, 'neigh_op_tnl_1')
// (18, 13, 'sp4_r_v_b_17')
// (18, 14, 'neigh_op_lft_1')
// (18, 14, 'sp4_h_r_31')
// (18, 14, 'sp4_h_r_47')
// (18, 14, 'sp4_r_v_b_4')
// (18, 15, 'neigh_op_bnl_1')
// (19, 6, 'sp4_v_t_42')
// (19, 7, 'sp4_v_b_42')
// (19, 8, 'sp4_v_b_31')
// (19, 9, 'local_g0_2')
// (19, 9, 'ram/RADDR_1')
// (19, 9, 'sp4_v_b_18')
// (19, 10, 'sp4_v_b_7')
// (19, 10, 'sp4_v_t_41')
// (19, 11, 'local_g3_1')
// (19, 11, 'ram/RADDR_1')
// (19, 11, 'sp4_r_v_b_36')
// (19, 11, 'sp4_v_b_41')
// (19, 12, 'sp4_r_v_b_25')
// (19, 12, 'sp4_v_b_28')
// (19, 13, 'local_g2_4')
// (19, 13, 'ram/RADDR_1')
// (19, 13, 'sp4_r_v_b_12')
// (19, 13, 'sp4_v_b_17')
// (19, 14, 'sp4_h_l_47')
// (19, 14, 'sp4_h_r_42')
// (19, 14, 'sp4_r_v_b_1')
// (19, 14, 'sp4_v_b_4')
// (20, 10, 'sp4_v_t_36')
// (20, 11, 'sp4_v_b_36')
// (20, 12, 'sp4_v_b_25')
// (20, 13, 'sp4_v_b_12')
// (20, 14, 'sp4_h_l_42')
// (20, 14, 'sp4_v_b_1')

reg n2267 = 0;
// (15, 14, 'sp4_h_r_2')
// (16, 13, 'neigh_op_tnr_5')
// (16, 14, 'neigh_op_rgt_5')
// (16, 14, 'sp4_h_r_15')
// (16, 15, 'neigh_op_bnr_5')
// (17, 13, 'neigh_op_top_5')
// (17, 14, 'local_g1_5')
// (17, 14, 'lutff_5/in_1')
// (17, 14, 'lutff_5/out')
// (17, 14, 'sp4_h_r_26')
// (17, 15, 'neigh_op_bot_5')
// (18, 7, 'sp4_r_v_b_41')
// (18, 8, 'sp4_r_v_b_28')
// (18, 9, 'sp4_r_v_b_17')
// (18, 10, 'sp4_r_v_b_4')
// (18, 11, 'sp4_r_v_b_45')
// (18, 12, 'sp4_r_v_b_32')
// (18, 13, 'neigh_op_tnl_5')
// (18, 13, 'sp4_r_v_b_21')
// (18, 14, 'neigh_op_lft_5')
// (18, 14, 'sp4_h_r_39')
// (18, 14, 'sp4_r_v_b_8')
// (18, 15, 'neigh_op_bnl_5')
// (19, 6, 'sp4_v_t_41')
// (19, 7, 'sp4_v_b_41')
// (19, 8, 'sp4_v_b_28')
// (19, 9, 'local_g1_1')
// (19, 9, 'ram/RADDR_5')
// (19, 9, 'sp4_v_b_17')
// (19, 10, 'sp4_v_b_4')
// (19, 10, 'sp4_v_t_45')
// (19, 11, 'local_g3_5')
// (19, 11, 'ram/RADDR_5')
// (19, 11, 'sp4_v_b_45')
// (19, 12, 'sp4_v_b_32')
// (19, 13, 'local_g1_5')
// (19, 13, 'ram/RADDR_5')
// (19, 13, 'sp4_v_b_21')
// (19, 14, 'sp4_h_l_39')
// (19, 14, 'sp4_v_b_8')

wire n2268;
// (15, 14, 'sp4_r_v_b_38')
// (15, 15, 'neigh_op_tnr_7')
// (15, 15, 'sp4_r_v_b_27')
// (15, 16, 'neigh_op_rgt_7')
// (15, 16, 'sp4_h_r_3')
// (15, 16, 'sp4_r_v_b_14')
// (15, 17, 'neigh_op_bnr_7')
// (15, 17, 'sp4_r_v_b_3')
// (16, 13, 'sp4_v_t_38')
// (16, 14, 'sp4_v_b_38')
// (16, 15, 'local_g3_3')
// (16, 15, 'lutff_global/cen')
// (16, 15, 'neigh_op_top_7')
// (16, 15, 'sp4_v_b_27')
// (16, 16, 'local_g1_7')
// (16, 16, 'lutff_6/in_2')
// (16, 16, 'lutff_7/out')
// (16, 16, 'sp4_h_r_14')
// (16, 16, 'sp4_v_b_14')
// (16, 17, 'neigh_op_bot_7')
// (16, 17, 'sp4_v_b_3')
// (17, 15, 'neigh_op_tnl_7')
// (17, 16, 'local_g3_3')
// (17, 16, 'lutff_global/cen')
// (17, 16, 'neigh_op_lft_7')
// (17, 16, 'sp4_h_r_27')
// (17, 17, 'neigh_op_bnl_7')
// (18, 16, 'sp4_h_r_38')
// (19, 16, 'sp4_h_l_38')

wire n2269;
// (15, 15, 'lutff_2/cout')
// (15, 15, 'lutff_3/in_3')

reg n2270 = 0;
// (15, 15, 'neigh_op_tnr_0')
// (15, 16, 'neigh_op_rgt_0')
// (15, 17, 'neigh_op_bnr_0')
// (16, 15, 'neigh_op_top_0')
// (16, 16, 'local_g2_0')
// (16, 16, 'lutff_0/in_0')
// (16, 16, 'lutff_0/out')
// (16, 16, 'lutff_2/in_2')
// (16, 17, 'neigh_op_bot_0')
// (17, 15, 'local_g3_0')
// (17, 15, 'lutff_3/in_2')
// (17, 15, 'neigh_op_tnl_0')
// (17, 16, 'neigh_op_lft_0')
// (17, 17, 'neigh_op_bnl_0')

wire n2271;
// (15, 15, 'neigh_op_tnr_1')
// (15, 16, 'neigh_op_rgt_1')
// (15, 17, 'neigh_op_bnr_1')
// (16, 15, 'neigh_op_top_1')
// (16, 16, 'lutff_1/out')
// (16, 17, 'local_g1_1')
// (16, 17, 'lutff_5/in_1')
// (16, 17, 'neigh_op_bot_1')
// (17, 15, 'neigh_op_tnl_1')
// (17, 16, 'neigh_op_lft_1')
// (17, 17, 'neigh_op_bnl_1')

reg n2272 = 0;
// (15, 15, 'neigh_op_tnr_2')
// (15, 16, 'neigh_op_rgt_2')
// (15, 17, 'neigh_op_bnr_2')
// (16, 15, 'neigh_op_top_2')
// (16, 16, 'local_g2_2')
// (16, 16, 'local_g3_2')
// (16, 16, 'lutff_0/in_2')
// (16, 16, 'lutff_1/in_3')
// (16, 16, 'lutff_2/in_1')
// (16, 16, 'lutff_2/out')
// (16, 16, 'lutff_4/in_1')
// (16, 17, 'neigh_op_bot_2')
// (17, 15, 'local_g3_2')
// (17, 15, 'lutff_2/in_1')
// (17, 15, 'lutff_3/in_0')
// (17, 15, 'lutff_7/in_0')
// (17, 15, 'neigh_op_tnl_2')
// (17, 16, 'neigh_op_lft_2')
// (17, 17, 'neigh_op_bnl_2')

wire n2273;
// (15, 15, 'neigh_op_tnr_3')
// (15, 16, 'neigh_op_rgt_3')
// (15, 17, 'neigh_op_bnr_3')
// (16, 15, 'neigh_op_top_3')
// (16, 16, 'lutff_3/out')
// (16, 17, 'local_g1_3')
// (16, 17, 'lutff_global/cen')
// (16, 17, 'neigh_op_bot_3')
// (17, 15, 'neigh_op_tnl_3')
// (17, 16, 'neigh_op_lft_3')
// (17, 17, 'neigh_op_bnl_3')

reg n2274 = 0;
// (15, 15, 'neigh_op_tnr_6')
// (15, 16, 'neigh_op_rgt_6')
// (15, 17, 'neigh_op_bnr_6')
// (16, 15, 'neigh_op_top_6')
// (16, 15, 'sp4_r_v_b_40')
// (16, 16, 'local_g3_6')
// (16, 16, 'lutff_1/in_2')
// (16, 16, 'lutff_4/in_3')
// (16, 16, 'lutff_6/out')
// (16, 16, 'sp4_r_v_b_29')
// (16, 17, 'neigh_op_bot_6')
// (16, 17, 'sp4_r_v_b_16')
// (16, 18, 'sp4_r_v_b_5')
// (17, 14, 'sp4_h_r_10')
// (17, 14, 'sp4_v_t_40')
// (17, 15, 'neigh_op_tnl_6')
// (17, 15, 'sp4_v_b_40')
// (17, 16, 'neigh_op_lft_6')
// (17, 16, 'sp4_v_b_29')
// (17, 17, 'neigh_op_bnl_6')
// (17, 17, 'sp4_v_b_16')
// (17, 18, 'sp4_v_b_5')
// (18, 14, 'local_g0_7')
// (18, 14, 'lutff_0/in_3')
// (18, 14, 'lutff_3/in_0')
// (18, 14, 'sp4_h_r_23')
// (19, 14, 'sp4_h_r_34')
// (20, 14, 'sp4_h_r_47')
// (21, 14, 'sp4_h_l_47')

wire n2275;
// (15, 15, 'sp4_h_r_6')
// (16, 14, 'neigh_op_tnr_7')
// (16, 15, 'neigh_op_rgt_7')
// (16, 15, 'sp4_h_r_19')
// (16, 16, 'neigh_op_bnr_7')
// (17, 14, 'neigh_op_top_7')
// (17, 14, 'sp4_r_v_b_42')
// (17, 15, 'local_g3_7')
// (17, 15, 'lutff_1/in_1')
// (17, 15, 'lutff_7/out')
// (17, 15, 'sp4_h_r_30')
// (17, 15, 'sp4_r_v_b_31')
// (17, 16, 'neigh_op_bot_7')
// (17, 16, 'sp4_r_v_b_18')
// (17, 17, 'sp4_r_v_b_7')
// (18, 8, 'sp4_r_v_b_39')
// (18, 9, 'sp4_r_v_b_26')
// (18, 10, 'sp4_r_v_b_15')
// (18, 11, 'sp4_r_v_b_2')
// (18, 12, 'sp4_r_v_b_43')
// (18, 13, 'sp4_h_r_7')
// (18, 13, 'sp4_r_v_b_30')
// (18, 13, 'sp4_v_t_42')
// (18, 14, 'neigh_op_tnl_7')
// (18, 14, 'sp4_r_v_b_19')
// (18, 14, 'sp4_v_b_42')
// (18, 15, 'neigh_op_lft_7')
// (18, 15, 'sp4_h_r_43')
// (18, 15, 'sp4_r_v_b_6')
// (18, 15, 'sp4_v_b_31')
// (18, 16, 'neigh_op_bnl_7')
// (18, 16, 'sp4_v_b_18')
// (18, 17, 'sp4_v_b_7')
// (19, 7, 'sp4_v_t_39')
// (19, 8, 'sp4_v_b_39')
// (19, 9, 'local_g2_2')
// (19, 9, 'ram/RCLKE')
// (19, 9, 'sp4_v_b_26')
// (19, 10, 'sp4_v_b_15')
// (19, 11, 'local_g1_3')
// (19, 11, 'ram/RCLKE')
// (19, 11, 'sp4_h_r_11')
// (19, 11, 'sp4_v_b_2')
// (19, 11, 'sp4_v_t_43')
// (19, 12, 'sp4_v_b_43')
// (19, 13, 'local_g0_2')
// (19, 13, 'ram/RCLKE')
// (19, 13, 'sp4_h_r_18')
// (19, 13, 'sp4_v_b_30')
// (19, 14, 'sp4_v_b_19')
// (19, 15, 'sp4_h_l_43')
// (19, 15, 'sp4_v_b_6')
// (20, 11, 'sp4_h_r_22')
// (20, 13, 'sp4_h_r_31')
// (21, 11, 'sp4_h_r_35')
// (21, 13, 'sp4_h_r_42')
// (22, 11, 'sp4_h_r_46')
// (22, 13, 'sp4_h_l_42')
// (23, 11, 'sp4_h_l_46')

wire n2276;
// (15, 16, 'lutff_1/cout')
// (15, 16, 'lutff_2/in_3')

wire n2277;
// (15, 16, 'neigh_op_tnr_0')
// (15, 17, 'neigh_op_rgt_0')
// (15, 18, 'neigh_op_bnr_0')
// (16, 14, 'sp4_r_v_b_36')
// (16, 15, 'sp4_r_v_b_25')
// (16, 16, 'local_g0_0')
// (16, 16, 'lutff_2/in_0')
// (16, 16, 'lutff_4/in_2')
// (16, 16, 'neigh_op_top_0')
// (16, 16, 'sp4_r_v_b_12')
// (16, 17, 'lutff_0/out')
// (16, 17, 'sp4_r_v_b_1')
// (16, 18, 'neigh_op_bot_0')
// (17, 13, 'sp4_v_t_36')
// (17, 14, 'sp4_v_b_36')
// (17, 15, 'local_g2_1')
// (17, 15, 'lutff_4/in_3')
// (17, 15, 'sp4_v_b_25')
// (17, 16, 'neigh_op_tnl_0')
// (17, 16, 'sp4_v_b_12')
// (17, 17, 'neigh_op_lft_0')
// (17, 17, 'sp4_v_b_1')
// (17, 18, 'neigh_op_bnl_0')

wire n2278;
// (15, 16, 'neigh_op_tnr_3')
// (15, 17, 'neigh_op_rgt_3')
// (15, 18, 'neigh_op_bnr_3')
// (16, 16, 'local_g1_3')
// (16, 16, 'lutff_1/in_1')
// (16, 16, 'lutff_7/in_3')
// (16, 16, 'neigh_op_top_3')
// (16, 17, 'lutff_3/out')
// (16, 18, 'neigh_op_bot_3')
// (17, 16, 'neigh_op_tnl_3')
// (17, 17, 'neigh_op_lft_3')
// (17, 18, 'neigh_op_bnl_3')

reg n2279 = 0;
// (15, 16, 'sp4_r_v_b_45')
// (15, 17, 'sp4_r_v_b_32')
// (15, 18, 'neigh_op_tnr_4')
// (15, 18, 'sp4_r_v_b_21')
// (15, 19, 'neigh_op_rgt_4')
// (15, 19, 'sp4_r_v_b_8')
// (15, 20, 'neigh_op_bnr_4')
// (16, 15, 'sp4_v_t_45')
// (16, 16, 'sp4_v_b_45')
// (16, 17, 'local_g3_0')
// (16, 17, 'lutff_0/in_3')
// (16, 17, 'lutff_3/in_2')
// (16, 17, 'sp4_v_b_32')
// (16, 18, 'neigh_op_top_4')
// (16, 18, 'sp4_v_b_21')
// (16, 19, 'local_g2_4')
// (16, 19, 'lutff_4/in_2')
// (16, 19, 'lutff_4/out')
// (16, 19, 'sp4_v_b_8')
// (16, 20, 'neigh_op_bot_4')
// (17, 18, 'neigh_op_tnl_4')
// (17, 19, 'neigh_op_lft_4')
// (17, 20, 'neigh_op_bnl_4')

reg n2280 = 0;
// (15, 17, 'sp4_r_v_b_36')
// (15, 18, 'neigh_op_tnr_6')
// (15, 18, 'sp4_r_v_b_25')
// (15, 19, 'local_g3_6')
// (15, 19, 'lutff_3/in_2')
// (15, 19, 'neigh_op_rgt_6')
// (15, 19, 'sp4_r_v_b_12')
// (15, 20, 'neigh_op_bnr_6')
// (15, 20, 'sp4_r_v_b_1')
// (16, 16, 'sp4_v_t_36')
// (16, 17, 'local_g3_4')
// (16, 17, 'lutff_0/in_1')
// (16, 17, 'lutff_3/in_0')
// (16, 17, 'sp4_v_b_36')
// (16, 18, 'neigh_op_top_6')
// (16, 18, 'sp4_v_b_25')
// (16, 19, 'local_g2_6')
// (16, 19, 'lutff_3/in_1')
// (16, 19, 'lutff_6/in_0')
// (16, 19, 'lutff_6/out')
// (16, 19, 'sp4_v_b_12')
// (16, 20, 'neigh_op_bot_6')
// (16, 20, 'sp4_v_b_1')
// (17, 18, 'neigh_op_tnl_6')
// (17, 19, 'neigh_op_lft_6')
// (17, 20, 'neigh_op_bnl_6')

wire n2281;
// (15, 18, 'lutff_1/cout')
// (15, 18, 'lutff_2/in_3')

wire n2282;
// (15, 18, 'lutff_3/cout')
// (15, 18, 'lutff_4/in_3')

wire n2283;
// (15, 18, 'lutff_5/cout')
// (15, 18, 'lutff_6/in_3')

wire n2284;
// (15, 18, 'lutff_7/cout')
// (15, 19, 'carry_in')
// (15, 19, 'carry_in_mux')
// (15, 19, 'lutff_0/in_3')

wire n2285;
// (15, 18, 'neigh_op_tnr_0')
// (15, 19, 'neigh_op_rgt_0')
// (15, 20, 'neigh_op_bnr_0')
// (16, 18, 'neigh_op_top_0')
// (16, 19, 'local_g1_0')
// (16, 19, 'lutff_0/out')
// (16, 19, 'lutff_7/in_2')
// (16, 20, 'neigh_op_bot_0')
// (17, 18, 'neigh_op_tnl_0')
// (17, 19, 'neigh_op_lft_0')
// (17, 20, 'neigh_op_bnl_0')

wire n2286;
// (15, 18, 'neigh_op_tnr_2')
// (15, 19, 'neigh_op_rgt_2')
// (15, 20, 'neigh_op_bnr_2')
// (16, 18, 'neigh_op_top_2')
// (16, 19, 'local_g3_2')
// (16, 19, 'lutff_2/out')
// (16, 19, 'lutff_6/in_3')
// (16, 20, 'neigh_op_bot_2')
// (17, 18, 'neigh_op_tnl_2')
// (17, 19, 'neigh_op_lft_2')
// (17, 20, 'neigh_op_bnl_2')

wire n2287;
// (15, 18, 'neigh_op_tnr_5')
// (15, 18, 'sp4_r_v_b_39')
// (15, 19, 'local_g0_2')
// (15, 19, 'lutff_global/cen')
// (15, 19, 'neigh_op_rgt_5')
// (15, 19, 'sp4_r_v_b_26')
// (15, 20, 'neigh_op_bnr_5')
// (15, 20, 'sp4_r_v_b_15')
// (15, 21, 'sp4_r_v_b_2')
// (16, 17, 'sp4_v_t_39')
// (16, 18, 'neigh_op_top_5')
// (16, 18, 'sp4_v_b_39')
// (16, 19, 'lutff_5/out')
// (16, 19, 'sp4_v_b_26')
// (16, 20, 'neigh_op_bot_5')
// (16, 20, 'sp4_v_b_15')
// (16, 21, 'sp4_v_b_2')
// (17, 18, 'neigh_op_tnl_5')
// (17, 19, 'neigh_op_lft_5')
// (17, 20, 'neigh_op_bnl_5')

wire n2288;
// (15, 19, 'lutff_1/cout')
// (15, 19, 'lutff_2/in_3')

wire n2289;
// (15, 19, 'lutff_3/cout')
// (15, 19, 'lutff_4/in_3')

reg n2290 = 0;
// (15, 19, 'neigh_op_tnr_4')
// (15, 20, 'neigh_op_rgt_4')
// (15, 21, 'neigh_op_bnr_4')
// (16, 19, 'neigh_op_top_4')
// (16, 20, 'lutff_4/out')
// (16, 20, 'sp4_h_r_8')
// (16, 21, 'neigh_op_bot_4')
// (17, 19, 'neigh_op_tnl_4')
// (17, 20, 'neigh_op_lft_4')
// (17, 20, 'sp4_h_r_21')
// (17, 21, 'neigh_op_bnl_4')
// (18, 20, 'sp4_h_r_32')
// (19, 17, 'sp4_r_v_b_39')
// (19, 18, 'sp4_r_v_b_26')
// (19, 19, 'sp4_r_v_b_15')
// (19, 20, 'sp4_h_r_45')
// (19, 20, 'sp4_r_v_b_2')
// (20, 16, 'sp4_v_t_39')
// (20, 17, 'sp4_v_b_39')
// (20, 18, 'sp4_v_b_26')
// (20, 19, 'sp4_v_b_15')
// (20, 20, 'local_g1_2')
// (20, 20, 'lutff_5/in_2')
// (20, 20, 'sp4_h_l_45')
// (20, 20, 'sp4_v_b_2')

reg n2291 = 0;
// (15, 20, 'neigh_op_tnr_6')
// (15, 21, 'neigh_op_rgt_6')
// (15, 21, 'sp4_h_r_1')
// (15, 22, 'neigh_op_bnr_6')
// (16, 20, 'neigh_op_top_6')
// (16, 21, 'lutff_6/out')
// (16, 21, 'sp4_h_r_12')
// (16, 22, 'neigh_op_bot_6')
// (17, 20, 'neigh_op_tnl_6')
// (17, 21, 'neigh_op_lft_6')
// (17, 21, 'sp4_h_r_25')
// (17, 22, 'neigh_op_bnl_6')
// (18, 21, 'sp4_h_r_36')
// (19, 21, 'sp4_h_l_36')
// (19, 21, 'sp4_h_r_9')
// (20, 21, 'local_g0_4')
// (20, 21, 'lutff_3/in_3')
// (20, 21, 'sp4_h_r_20')
// (21, 21, 'sp4_h_r_33')
// (22, 21, 'sp4_h_r_44')
// (23, 21, 'sp4_h_l_44')

reg n2292 = 0;
// (15, 20, 'sp4_h_r_10')
// (16, 19, 'neigh_op_tnr_1')
// (16, 20, 'neigh_op_rgt_1')
// (16, 20, 'sp4_h_r_23')
// (16, 21, 'neigh_op_bnr_1')
// (17, 18, 'sp4_r_v_b_43')
// (17, 19, 'local_g0_1')
// (17, 19, 'lutff_1/in_2')
// (17, 19, 'neigh_op_top_1')
// (17, 19, 'sp4_r_v_b_30')
// (17, 20, 'local_g0_1')
// (17, 20, 'local_g3_1')
// (17, 20, 'lutff_1/in_3')
// (17, 20, 'lutff_1/out')
// (17, 20, 'lutff_6/in_1')
// (17, 20, 'sp4_h_r_2')
// (17, 20, 'sp4_h_r_34')
// (17, 20, 'sp4_r_v_b_19')
// (17, 21, 'local_g1_1')
// (17, 21, 'lutff_0/in_2')
// (17, 21, 'lutff_2/in_2')
// (17, 21, 'lutff_5/in_1')
// (17, 21, 'lutff_7/in_1')
// (17, 21, 'neigh_op_bot_1')
// (17, 21, 'sp4_r_v_b_6')
// (18, 17, 'sp4_v_t_43')
// (18, 18, 'sp4_v_b_43')
// (18, 19, 'neigh_op_tnl_1')
// (18, 19, 'sp4_v_b_30')
// (18, 20, 'neigh_op_lft_1')
// (18, 20, 'sp4_h_r_15')
// (18, 20, 'sp4_h_r_47')
// (18, 20, 'sp4_v_b_19')
// (18, 21, 'neigh_op_bnl_1')
// (18, 21, 'sp4_h_r_6')
// (18, 21, 'sp4_v_b_6')
// (19, 20, 'sp4_h_l_47')
// (19, 20, 'sp4_h_r_1')
// (19, 20, 'sp4_h_r_26')
// (19, 21, 'sp4_h_r_19')
// (20, 17, 'sp4_r_v_b_39')
// (20, 18, 'sp4_r_v_b_26')
// (20, 19, 'sp4_r_v_b_15')
// (20, 20, 'sp4_h_r_12')
// (20, 20, 'sp4_h_r_39')
// (20, 20, 'sp4_r_v_b_2')
// (20, 21, 'sp4_h_r_30')
// (21, 16, 'sp4_v_t_39')
// (21, 17, 'sp4_v_b_39')
// (21, 18, 'sp4_v_b_26')
// (21, 19, 'local_g0_7')
// (21, 19, 'lutff_3/in_2')
// (21, 19, 'sp4_v_b_15')
// (21, 20, 'sp4_h_l_39')
// (21, 20, 'sp4_h_r_25')
// (21, 20, 'sp4_v_b_2')
// (21, 21, 'local_g3_3')
// (21, 21, 'lutff_6/in_2')
// (21, 21, 'sp4_h_r_43')
// (22, 17, 'sp4_r_v_b_42')
// (22, 18, 'sp4_r_v_b_31')
// (22, 19, 'local_g3_2')
// (22, 19, 'lutff_5/in_0')
// (22, 19, 'lutff_7/in_0')
// (22, 19, 'sp4_r_v_b_18')
// (22, 20, 'sp4_h_r_36')
// (22, 20, 'sp4_r_v_b_7')
// (22, 21, 'sp4_h_l_43')
// (23, 16, 'sp4_v_t_42')
// (23, 17, 'sp4_v_b_42')
// (23, 18, 'sp4_v_b_31')
// (23, 19, 'sp4_v_b_18')
// (23, 20, 'sp4_h_l_36')
// (23, 20, 'sp4_v_b_7')

reg n2293 = 0;
// (15, 20, 'sp4_h_r_6')
// (15, 21, 'sp4_r_v_b_44')
// (15, 22, 'sp4_r_v_b_33')
// (15, 23, 'sp4_r_v_b_20')
// (15, 24, 'sp4_r_v_b_9')
// (16, 19, 'local_g2_7')
// (16, 19, 'lutff_5/in_2')
// (16, 19, 'neigh_op_tnr_7')
// (16, 20, 'local_g2_7')
// (16, 20, 'lutff_2/in_1')
// (16, 20, 'lutff_6/in_1')
// (16, 20, 'neigh_op_rgt_7')
// (16, 20, 'sp4_h_r_19')
// (16, 20, 'sp4_h_r_3')
// (16, 20, 'sp4_r_v_b_46')
// (16, 20, 'sp4_v_t_44')
// (16, 21, 'local_g1_7')
// (16, 21, 'lutff_7/in_3')
// (16, 21, 'neigh_op_bnr_7')
// (16, 21, 'sp4_r_v_b_35')
// (16, 21, 'sp4_v_b_44')
// (16, 22, 'local_g3_6')
// (16, 22, 'lutff_2/in_3')
// (16, 22, 'sp4_r_v_b_22')
// (16, 22, 'sp4_v_b_33')
// (16, 23, 'local_g2_3')
// (16, 23, 'lutff_0/in_3')
// (16, 23, 'lutff_7/in_2')
// (16, 23, 'sp4_r_v_b_11')
// (16, 23, 'sp4_v_b_20')
// (16, 24, 'local_g0_1')
// (16, 24, 'lutff_3/in_0')
// (16, 24, 'sp4_v_b_9')
// (17, 14, 'sp4_r_v_b_47')
// (17, 15, 'sp4_r_v_b_34')
// (17, 16, 'sp4_r_v_b_23')
// (17, 17, 'sp4_r_v_b_10')
// (17, 18, 'sp4_r_v_b_39')
// (17, 19, 'local_g1_7')
// (17, 19, 'lutff_7/in_1')
// (17, 19, 'neigh_op_top_7')
// (17, 19, 'sp4_r_v_b_26')
// (17, 19, 'sp4_r_v_b_42')
// (17, 19, 'sp4_v_t_46')
// (17, 20, 'local_g3_7')
// (17, 20, 'lutff_7/in_3')
// (17, 20, 'lutff_7/out')
// (17, 20, 'sp4_h_r_14')
// (17, 20, 'sp4_h_r_30')
// (17, 20, 'sp4_r_v_b_15')
// (17, 20, 'sp4_r_v_b_31')
// (17, 20, 'sp4_r_v_b_47')
// (17, 20, 'sp4_v_b_46')
// (17, 21, 'local_g1_7')
// (17, 21, 'lutff_1/in_3')
// (17, 21, 'lutff_4/in_2')
// (17, 21, 'neigh_op_bot_7')
// (17, 21, 'sp4_r_v_b_18')
// (17, 21, 'sp4_r_v_b_2')
// (17, 21, 'sp4_r_v_b_34')
// (17, 21, 'sp4_v_b_35')
// (17, 22, 'local_g0_6')
// (17, 22, 'lutff_6/in_0')
// (17, 22, 'sp4_r_v_b_23')
// (17, 22, 'sp4_r_v_b_39')
// (17, 22, 'sp4_r_v_b_7')
// (17, 22, 'sp4_v_b_22')
// (17, 23, 'local_g1_3')
// (17, 23, 'lutff_2/in_0')
// (17, 23, 'sp4_r_v_b_10')
// (17, 23, 'sp4_r_v_b_26')
// (17, 23, 'sp4_v_b_11')
// (17, 24, 'local_g2_7')
// (17, 24, 'lutff_7/in_2')
// (17, 24, 'sp4_r_v_b_15')
// (17, 25, 'sp4_r_v_b_2')
// (18, 13, 'sp4_v_t_47')
// (18, 14, 'sp4_v_b_47')
// (18, 15, 'local_g3_2')
// (18, 15, 'lutff_5/in_0')
// (18, 15, 'sp4_v_b_34')
// (18, 16, 'sp4_v_b_23')
// (18, 17, 'local_g1_2')
// (18, 17, 'lutff_3/in_2')
// (18, 17, 'sp4_h_r_2')
// (18, 17, 'sp4_v_b_10')
// (18, 17, 'sp4_v_t_39')
// (18, 18, 'local_g3_7')
// (18, 18, 'lutff_2/in_2')
// (18, 18, 'sp4_h_r_0')
// (18, 18, 'sp4_h_r_7')
// (18, 18, 'sp4_v_b_39')
// (18, 18, 'sp4_v_t_42')
// (18, 19, 'local_g3_7')
// (18, 19, 'lutff_2/in_0')
// (18, 19, 'lutff_7/in_3')
// (18, 19, 'neigh_op_tnl_7')
// (18, 19, 'sp4_h_r_10')
// (18, 19, 'sp4_v_b_26')
// (18, 19, 'sp4_v_b_42')
// (18, 19, 'sp4_v_t_47')
// (18, 20, 'local_g0_7')
// (18, 20, 'lutff_7/in_0')
// (18, 20, 'neigh_op_lft_7')
// (18, 20, 'sp4_h_r_27')
// (18, 20, 'sp4_h_r_43')
// (18, 20, 'sp4_v_b_15')
// (18, 20, 'sp4_v_b_31')
// (18, 20, 'sp4_v_b_47')
// (18, 21, 'local_g3_7')
// (18, 21, 'lutff_2/in_0')
// (18, 21, 'neigh_op_bnl_7')
// (18, 21, 'sp4_h_r_8')
// (18, 21, 'sp4_v_b_18')
// (18, 21, 'sp4_v_b_2')
// (18, 21, 'sp4_v_b_34')
// (18, 21, 'sp4_v_t_39')
// (18, 22, 'local_g0_7')
// (18, 22, 'lutff_4/in_3')
// (18, 22, 'sp4_h_r_7')
// (18, 22, 'sp4_v_b_23')
// (18, 22, 'sp4_v_b_39')
// (18, 22, 'sp4_v_b_7')
// (18, 23, 'sp4_h_r_10')
// (18, 23, 'sp4_v_b_10')
// (18, 23, 'sp4_v_b_26')
// (18, 24, 'local_g0_7')
// (18, 24, 'lutff_4/in_1')
// (18, 24, 'sp4_v_b_15')
// (18, 25, 'sp4_v_b_2')
// (19, 13, 'sp4_r_v_b_46')
// (19, 14, 'sp4_r_v_b_35')
// (19, 15, 'sp4_r_v_b_22')
// (19, 16, 'sp4_r_v_b_11')
// (19, 17, 'sp4_h_r_15')
// (19, 17, 'sp4_r_v_b_38')
// (19, 18, 'sp4_h_r_13')
// (19, 18, 'sp4_h_r_18')
// (19, 18, 'sp4_r_v_b_27')
// (19, 19, 'sp4_h_r_23')
// (19, 19, 'sp4_r_v_b_14')
// (19, 20, 'sp4_h_l_43')
// (19, 20, 'sp4_h_r_38')
// (19, 20, 'sp4_h_r_6')
// (19, 20, 'sp4_h_r_9')
// (19, 20, 'sp4_r_v_b_3')
// (19, 21, 'sp4_h_r_21')
// (19, 21, 'sp4_r_v_b_45')
// (19, 22, 'sp4_h_r_18')
// (19, 22, 'sp4_r_v_b_32')
// (19, 23, 'sp4_h_r_23')
// (19, 23, 'sp4_r_v_b_21')
// (19, 24, 'sp4_r_v_b_8')
// (20, 12, 'sp4_v_t_46')
// (20, 13, 'sp4_v_b_46')
// (20, 14, 'sp4_v_b_35')
// (20, 15, 'local_g1_6')
// (20, 15, 'lutff_5/in_2')
// (20, 15, 'sp4_v_b_22')
// (20, 16, 'sp4_v_b_11')
// (20, 16, 'sp4_v_t_38')
// (20, 17, 'local_g3_2')
// (20, 17, 'lutff_7/in_0')
// (20, 17, 'sp4_h_r_26')
// (20, 17, 'sp4_v_b_38')
// (20, 18, 'local_g2_0')
// (20, 18, 'lutff_5/in_1')
// (20, 18, 'sp4_h_r_24')
// (20, 18, 'sp4_h_r_31')
// (20, 18, 'sp4_v_b_27')
// (20, 19, 'sp4_h_r_34')
// (20, 19, 'sp4_v_b_14')
// (20, 20, 'local_g0_3')
// (20, 20, 'local_g0_4')
// (20, 20, 'lutff_0/in_1')
// (20, 20, 'lutff_4/in_0')
// (20, 20, 'lutff_6/in_3')
// (20, 20, 'sp4_h_l_38')
// (20, 20, 'sp4_h_r_11')
// (20, 20, 'sp4_h_r_19')
// (20, 20, 'sp4_h_r_20')
// (20, 20, 'sp4_v_b_3')
// (20, 20, 'sp4_v_t_45')
// (20, 21, 'local_g3_0')
// (20, 21, 'lutff_6/in_1')
// (20, 21, 'sp4_h_r_32')
// (20, 21, 'sp4_v_b_45')
// (20, 22, 'local_g3_0')
// (20, 22, 'lutff_4/in_1')
// (20, 22, 'sp4_h_r_31')
// (20, 22, 'sp4_v_b_32')
// (20, 23, 'local_g0_5')
// (20, 23, 'lutff_3/in_2')
// (20, 23, 'sp4_h_r_34')
// (20, 23, 'sp4_v_b_21')
// (20, 24, 'sp4_v_b_8')
// (21, 14, 'sp4_r_v_b_39')
// (21, 14, 'sp4_r_v_b_45')
// (21, 15, 'sp4_r_v_b_26')
// (21, 15, 'sp4_r_v_b_32')
// (21, 16, 'local_g3_5')
// (21, 16, 'lutff_5/in_1')
// (21, 16, 'sp4_r_v_b_15')
// (21, 16, 'sp4_r_v_b_21')
// (21, 17, 'local_g2_7')
// (21, 17, 'lutff_1/in_0')
// (21, 17, 'lutff_6/in_1')
// (21, 17, 'sp4_h_r_39')
// (21, 17, 'sp4_r_v_b_2')
// (21, 17, 'sp4_r_v_b_8')
// (21, 18, 'local_g3_2')
// (21, 18, 'lutff_6/in_1')
// (21, 18, 'sp4_h_r_37')
// (21, 18, 'sp4_h_r_42')
// (21, 19, 'local_g3_7')
// (21, 19, 'lutff_7/in_3')
// (21, 19, 'sp4_h_r_47')
// (21, 20, 'local_g0_6')
// (21, 20, 'lutff_5/in_1')
// (21, 20, 'sp4_h_r_22')
// (21, 20, 'sp4_h_r_30')
// (21, 20, 'sp4_h_r_33')
// (21, 21, 'local_g3_5')
// (21, 21, 'lutff_3/in_1')
// (21, 21, 'sp4_h_r_45')
// (21, 22, 'local_g2_2')
// (21, 22, 'lutff_5/in_1')
// (21, 22, 'sp4_h_r_42')
// (21, 23, 'local_g2_7')
// (21, 23, 'lutff_4/in_3')
// (21, 23, 'lutff_7/in_0')
// (21, 23, 'sp4_h_r_47')
// (22, 13, 'sp4_v_t_39')
// (22, 13, 'sp4_v_t_45')
// (22, 14, 'sp4_v_b_39')
// (22, 14, 'sp4_v_b_45')
// (22, 15, 'sp4_v_b_26')
// (22, 15, 'sp4_v_b_32')
// (22, 16, 'local_g0_7')
// (22, 16, 'lutff_4/in_3')
// (22, 16, 'lutff_5/in_2')
// (22, 16, 'lutff_6/in_3')
// (22, 16, 'lutff_7/in_2')
// (22, 16, 'sp4_v_b_15')
// (22, 16, 'sp4_v_b_21')
// (22, 17, 'local_g1_5')
// (22, 17, 'lutff_1/in_1')
// (22, 17, 'lutff_3/in_3')
// (22, 17, 'lutff_4/in_0')
// (22, 17, 'lutff_6/in_0')
// (22, 17, 'sp4_h_l_39')
// (22, 17, 'sp4_h_r_5')
// (22, 17, 'sp4_r_v_b_43')
// (22, 17, 'sp4_v_b_2')
// (22, 17, 'sp4_v_b_8')
// (22, 18, 'local_g0_3')
// (22, 18, 'local_g1_3')
// (22, 18, 'lutff_0/in_2')
// (22, 18, 'lutff_1/in_3')
// (22, 18, 'lutff_3/in_0')
// (22, 18, 'sp4_h_l_37')
// (22, 18, 'sp4_h_l_42')
// (22, 18, 'sp4_h_r_3')
// (22, 18, 'sp4_r_v_b_30')
// (22, 19, 'local_g3_3')
// (22, 19, 'lutff_0/in_2')
// (22, 19, 'lutff_4/in_2')
// (22, 19, 'lutff_6/in_0')
// (22, 19, 'sp4_h_l_47')
// (22, 19, 'sp4_r_v_b_19')
// (22, 20, 'local_g3_3')
// (22, 20, 'local_g3_4')
// (22, 20, 'lutff_2/in_2')
// (22, 20, 'lutff_3/in_3')
// (22, 20, 'lutff_4/in_0')
// (22, 20, 'lutff_6/in_0')
// (22, 20, 'lutff_7/in_2')
// (22, 20, 'sp4_h_r_35')
// (22, 20, 'sp4_h_r_43')
// (22, 20, 'sp4_h_r_44')
// (22, 20, 'sp4_r_v_b_6')
// (22, 21, 'local_g1_3')
// (22, 21, 'lutff_7/in_3')
// (22, 21, 'sp4_h_l_45')
// (22, 21, 'sp4_h_r_11')
// (22, 22, 'local_g1_7')
// (22, 22, 'lutff_3/in_1')
// (22, 22, 'lutff_7/in_3')
// (22, 22, 'sp4_h_l_42')
// (22, 22, 'sp4_h_r_7')
// (22, 23, 'local_g1_1')
// (22, 23, 'lutff_1/in_1')
// (22, 23, 'sp4_h_l_47')
// (22, 23, 'sp4_h_r_1')
// (23, 16, 'sp4_v_t_43')
// (23, 17, 'sp4_h_r_16')
// (23, 17, 'sp4_v_b_43')
// (23, 18, 'sp4_h_r_14')
// (23, 18, 'sp4_v_b_30')
// (23, 19, 'sp4_v_b_19')
// (23, 20, 'sp4_h_l_43')
// (23, 20, 'sp4_h_l_44')
// (23, 20, 'sp4_h_r_46')
// (23, 20, 'sp4_v_b_6')
// (23, 21, 'sp4_h_r_22')
// (23, 22, 'sp4_h_r_18')
// (23, 23, 'sp4_h_r_12')
// (24, 17, 'sp4_h_r_29')
// (24, 18, 'sp4_h_r_27')
// (24, 20, 'sp4_h_l_46')
// (24, 21, 'sp4_h_r_35')
// (24, 22, 'sp4_h_r_31')
// (24, 23, 'sp4_h_r_25')
// (25, 17, 'sp4_h_r_40')
// (25, 18, 'sp4_h_r_38')
// (25, 21, 'sp4_h_r_46')
// (25, 22, 'sp4_h_r_42')
// (25, 23, 'sp4_h_r_36')

wire n2294;
// (15, 21, 'neigh_op_tnr_2')
// (15, 22, 'neigh_op_rgt_2')
// (15, 23, 'neigh_op_bnr_2')
// (16, 21, 'neigh_op_top_2')
// (16, 22, 'local_g0_2')
// (16, 22, 'lutff_2/out')
// (16, 22, 'lutff_global/cen')
// (16, 23, 'neigh_op_bot_2')
// (17, 21, 'neigh_op_tnl_2')
// (17, 22, 'neigh_op_lft_2')
// (17, 23, 'neigh_op_bnl_2')

reg n2295 = 0;
// (15, 21, 'neigh_op_tnr_6')
// (15, 22, 'neigh_op_rgt_6')
// (15, 23, 'neigh_op_bnr_6')
// (16, 21, 'neigh_op_top_6')
// (16, 22, 'lutff_6/out')
// (16, 23, 'neigh_op_bot_6')
// (17, 21, 'neigh_op_tnl_6')
// (17, 22, 'local_g1_6')
// (17, 22, 'lutff_5/in_0')
// (17, 22, 'neigh_op_lft_6')
// (17, 23, 'neigh_op_bnl_6')

wire n2296;
// (15, 21, 'sp4_h_r_2')
// (16, 20, 'neigh_op_tnr_5')
// (16, 20, 'sp4_r_v_b_39')
// (16, 21, 'neigh_op_rgt_5')
// (16, 21, 'sp4_h_r_15')
// (16, 21, 'sp4_r_v_b_26')
// (16, 22, 'neigh_op_bnr_5')
// (16, 22, 'sp4_r_v_b_15')
// (16, 23, 'local_g1_2')
// (16, 23, 'lutff_0/in_1')
// (16, 23, 'lutff_7/in_0')
// (16, 23, 'sp4_r_v_b_2')
// (17, 19, 'sp4_v_t_39')
// (17, 20, 'neigh_op_top_5')
// (17, 20, 'sp4_r_v_b_38')
// (17, 20, 'sp4_v_b_39')
// (17, 21, 'lutff_5/out')
// (17, 21, 'sp4_h_r_10')
// (17, 21, 'sp4_h_r_26')
// (17, 21, 'sp4_r_v_b_27')
// (17, 21, 'sp4_v_b_26')
// (17, 22, 'neigh_op_bot_5')
// (17, 22, 'sp4_r_v_b_14')
// (17, 22, 'sp4_v_b_15')
// (17, 23, 'sp4_r_v_b_3')
// (17, 23, 'sp4_v_b_2')
// (18, 19, 'sp4_v_t_38')
// (18, 20, 'local_g3_5')
// (18, 20, 'lutff_7/in_3')
// (18, 20, 'neigh_op_tnl_5')
// (18, 20, 'sp4_v_b_38')
// (18, 21, 'neigh_op_lft_5')
// (18, 21, 'sp4_h_r_23')
// (18, 21, 'sp4_h_r_39')
// (18, 21, 'sp4_v_b_27')
// (18, 22, 'local_g2_5')
// (18, 22, 'lutff_4/in_1')
// (18, 22, 'neigh_op_bnl_5')
// (18, 22, 'sp4_v_b_14')
// (18, 23, 'sp4_h_r_3')
// (18, 23, 'sp4_v_b_3')
// (19, 21, 'sp4_h_l_39')
// (19, 21, 'sp4_h_r_2')
// (19, 21, 'sp4_h_r_34')
// (19, 23, 'sp4_h_r_14')
// (20, 18, 'sp4_r_v_b_47')
// (20, 19, 'sp4_r_v_b_34')
// (20, 20, 'local_g3_7')
// (20, 20, 'lutff_6/in_2')
// (20, 20, 'sp4_r_v_b_23')
// (20, 21, 'sp4_h_r_15')
// (20, 21, 'sp4_h_r_47')
// (20, 21, 'sp4_r_v_b_10')
// (20, 22, 'sp4_r_v_b_47')
// (20, 23, 'sp4_h_r_27')
// (20, 23, 'sp4_r_v_b_34')
// (20, 24, 'sp4_r_v_b_23')
// (20, 25, 'sp4_r_v_b_10')
// (21, 17, 'sp4_v_t_47')
// (21, 18, 'sp4_v_b_47')
// (21, 19, 'sp4_v_b_34')
// (21, 20, 'sp4_r_v_b_38')
// (21, 20, 'sp4_v_b_23')
// (21, 21, 'sp4_h_l_47')
// (21, 21, 'sp4_h_r_26')
// (21, 21, 'sp4_r_v_b_27')
// (21, 21, 'sp4_v_b_10')
// (21, 21, 'sp4_v_t_47')
// (21, 22, 'sp4_r_v_b_14')
// (21, 22, 'sp4_v_b_47')
// (21, 23, 'local_g2_2')
// (21, 23, 'lutff_7/in_3')
// (21, 23, 'sp4_h_r_38')
// (21, 23, 'sp4_r_v_b_3')
// (21, 23, 'sp4_v_b_34')
// (21, 24, 'sp4_v_b_23')
// (21, 25, 'sp4_v_b_10')
// (22, 18, 'sp4_r_v_b_45')
// (22, 19, 'sp4_r_v_b_32')
// (22, 19, 'sp4_v_t_38')
// (22, 20, 'local_g3_5')
// (22, 20, 'lutff_2/in_0')
// (22, 20, 'sp4_r_v_b_21')
// (22, 20, 'sp4_v_b_38')
// (22, 21, 'sp4_h_r_39')
// (22, 21, 'sp4_r_v_b_8')
// (22, 21, 'sp4_v_b_27')
// (22, 22, 'local_g0_6')
// (22, 22, 'lutff_3/in_3')
// (22, 22, 'sp4_v_b_14')
// (22, 23, 'sp4_h_l_38')
// (22, 23, 'sp4_v_b_3')
// (23, 17, 'sp4_v_t_45')
// (23, 18, 'sp4_v_b_45')
// (23, 19, 'sp4_v_b_32')
// (23, 20, 'sp4_v_b_21')
// (23, 21, 'sp4_h_l_39')
// (23, 21, 'sp4_v_b_8')

reg n2297 = 0;
// (15, 21, 'sp4_r_v_b_40')
// (15, 22, 'sp4_r_v_b_29')
// (15, 23, 'sp4_r_v_b_16')
// (15, 24, 'sp4_r_v_b_5')
// (16, 18, 'sp4_r_v_b_40')
// (16, 19, 'local_g2_0')
// (16, 19, 'lutff_5/in_1')
// (16, 19, 'neigh_op_tnr_0')
// (16, 19, 'sp4_r_v_b_29')
// (16, 19, 'sp4_r_v_b_45')
// (16, 20, 'local_g3_0')
// (16, 20, 'lutff_2/in_3')
// (16, 20, 'lutff_6/in_3')
// (16, 20, 'neigh_op_rgt_0')
// (16, 20, 'sp4_h_r_5')
// (16, 20, 'sp4_r_v_b_16')
// (16, 20, 'sp4_r_v_b_32')
// (16, 20, 'sp4_v_t_40')
// (16, 21, 'local_g1_0')
// (16, 21, 'lutff_7/in_0')
// (16, 21, 'neigh_op_bnr_0')
// (16, 21, 'sp4_r_v_b_21')
// (16, 21, 'sp4_r_v_b_43')
// (16, 21, 'sp4_r_v_b_5')
// (16, 21, 'sp4_v_b_40')
// (16, 22, 'local_g2_0')
// (16, 22, 'lutff_2/in_2')
// (16, 22, 'sp4_r_v_b_30')
// (16, 22, 'sp4_r_v_b_8')
// (16, 22, 'sp4_v_b_29')
// (16, 23, 'local_g0_0')
// (16, 23, 'lutff_0/in_2')
// (16, 23, 'lutff_7/in_1')
// (16, 23, 'sp4_r_v_b_19')
// (16, 23, 'sp4_v_b_16')
// (16, 24, 'local_g1_5')
// (16, 24, 'lutff_3/in_3')
// (16, 24, 'sp4_r_v_b_6')
// (16, 24, 'sp4_v_b_5')
// (17, 13, 'sp4_r_v_b_44')
// (17, 14, 'sp4_r_v_b_33')
// (17, 15, 'sp4_r_v_b_20')
// (17, 16, 'sp4_r_v_b_9')
// (17, 17, 'sp4_h_r_5')
// (17, 17, 'sp4_r_v_b_36')
// (17, 17, 'sp4_v_t_40')
// (17, 18, 'sp4_h_r_8')
// (17, 18, 'sp4_r_v_b_25')
// (17, 18, 'sp4_r_v_b_41')
// (17, 18, 'sp4_v_b_40')
// (17, 18, 'sp4_v_t_45')
// (17, 19, 'neigh_op_top_0')
// (17, 19, 'sp4_r_v_b_12')
// (17, 19, 'sp4_r_v_b_28')
// (17, 19, 'sp4_r_v_b_44')
// (17, 19, 'sp4_v_b_29')
// (17, 19, 'sp4_v_b_45')
// (17, 20, 'local_g2_0')
// (17, 20, 'lutff_0/in_2')
// (17, 20, 'lutff_0/out')
// (17, 20, 'sp4_h_r_0')
// (17, 20, 'sp4_h_r_16')
// (17, 20, 'sp4_r_v_b_1')
// (17, 20, 'sp4_r_v_b_17')
// (17, 20, 'sp4_r_v_b_33')
// (17, 20, 'sp4_v_b_16')
// (17, 20, 'sp4_v_b_32')
// (17, 20, 'sp4_v_t_43')
// (17, 21, 'local_g0_0')
// (17, 21, 'lutff_1/in_1')
// (17, 21, 'lutff_4/in_0')
// (17, 21, 'neigh_op_bot_0')
// (17, 21, 'sp4_r_v_b_20')
// (17, 21, 'sp4_r_v_b_4')
// (17, 21, 'sp4_v_b_21')
// (17, 21, 'sp4_v_b_43')
// (17, 21, 'sp4_v_b_5')
// (17, 22, 'local_g2_1')
// (17, 22, 'lutff_6/in_3')
// (17, 22, 'sp4_r_v_b_41')
// (17, 22, 'sp4_r_v_b_9')
// (17, 22, 'sp4_v_b_30')
// (17, 22, 'sp4_v_b_8')
// (17, 23, 'local_g0_3')
// (17, 23, 'lutff_2/in_3')
// (17, 23, 'sp4_r_v_b_28')
// (17, 23, 'sp4_v_b_19')
// (17, 24, 'local_g0_6')
// (17, 24, 'lutff_7/in_3')
// (17, 24, 'sp4_r_v_b_17')
// (17, 24, 'sp4_v_b_6')
// (17, 25, 'sp4_r_v_b_4')
// (18, 12, 'sp4_v_t_44')
// (18, 13, 'sp4_v_b_44')
// (18, 14, 'sp4_v_b_33')
// (18, 15, 'local_g0_4')
// (18, 15, 'lutff_5/in_1')
// (18, 15, 'sp4_v_b_20')
// (18, 16, 'sp4_h_r_1')
// (18, 16, 'sp4_v_b_9')
// (18, 16, 'sp4_v_t_36')
// (18, 17, 'local_g2_4')
// (18, 17, 'lutff_3/in_1')
// (18, 17, 'sp4_h_r_16')
// (18, 17, 'sp4_h_r_4')
// (18, 17, 'sp4_v_b_36')
// (18, 17, 'sp4_v_t_41')
// (18, 18, 'local_g3_1')
// (18, 18, 'lutff_2/in_0')
// (18, 18, 'sp4_h_r_21')
// (18, 18, 'sp4_v_b_25')
// (18, 18, 'sp4_v_b_41')
// (18, 18, 'sp4_v_t_44')
// (18, 19, 'local_g2_0')
// (18, 19, 'lutff_2/in_2')
// (18, 19, 'lutff_7/in_1')
// (18, 19, 'neigh_op_tnl_0')
// (18, 19, 'sp4_v_b_12')
// (18, 19, 'sp4_v_b_28')
// (18, 19, 'sp4_v_b_44')
// (18, 20, 'local_g1_0')
// (18, 20, 'lutff_7/in_2')
// (18, 20, 'neigh_op_lft_0')
// (18, 20, 'sp4_h_r_1')
// (18, 20, 'sp4_h_r_13')
// (18, 20, 'sp4_h_r_29')
// (18, 20, 'sp4_v_b_1')
// (18, 20, 'sp4_v_b_17')
// (18, 20, 'sp4_v_b_33')
// (18, 21, 'local_g3_0')
// (18, 21, 'lutff_2/in_3')
// (18, 21, 'neigh_op_bnl_0')
// (18, 21, 'sp4_h_r_10')
// (18, 21, 'sp4_v_b_20')
// (18, 21, 'sp4_v_b_4')
// (18, 21, 'sp4_v_t_41')
// (18, 22, 'local_g1_1')
// (18, 22, 'lutff_4/in_0')
// (18, 22, 'sp4_h_r_9')
// (18, 22, 'sp4_v_b_41')
// (18, 22, 'sp4_v_b_9')
// (18, 23, 'sp4_v_b_28')
// (18, 24, 'local_g1_1')
// (18, 24, 'lutff_4/in_2')
// (18, 24, 'sp4_v_b_17')
// (18, 25, 'sp4_v_b_4')
// (19, 13, 'sp4_r_v_b_36')
// (19, 14, 'sp4_r_v_b_25')
// (19, 15, 'sp4_r_v_b_12')
// (19, 16, 'sp4_h_r_12')
// (19, 16, 'sp4_r_v_b_1')
// (19, 17, 'sp4_h_r_17')
// (19, 17, 'sp4_h_r_29')
// (19, 17, 'sp4_r_v_b_40')
// (19, 18, 'sp4_h_r_32')
// (19, 18, 'sp4_r_v_b_29')
// (19, 19, 'sp4_r_v_b_16')
// (19, 20, 'sp4_h_r_12')
// (19, 20, 'sp4_h_r_24')
// (19, 20, 'sp4_h_r_40')
// (19, 20, 'sp4_r_v_b_5')
// (19, 21, 'sp4_h_r_23')
// (19, 21, 'sp4_r_v_b_47')
// (19, 22, 'sp4_h_r_20')
// (19, 22, 'sp4_r_v_b_34')
// (19, 23, 'sp4_r_v_b_23')
// (19, 24, 'sp4_r_v_b_10')
// (20, 12, 'sp4_v_t_36')
// (20, 13, 'sp4_v_b_36')
// (20, 14, 'sp4_v_b_25')
// (20, 15, 'local_g1_4')
// (20, 15, 'lutff_5/in_0')
// (20, 15, 'sp4_v_b_12')
// (20, 16, 'sp4_h_r_25')
// (20, 16, 'sp4_v_b_1')
// (20, 16, 'sp4_v_t_40')
// (20, 17, 'local_g2_0')
// (20, 17, 'lutff_7/in_3')
// (20, 17, 'sp4_h_r_28')
// (20, 17, 'sp4_h_r_40')
// (20, 17, 'sp4_r_v_b_43')
// (20, 17, 'sp4_v_b_40')
// (20, 18, 'local_g2_5')
// (20, 18, 'lutff_5/in_0')
// (20, 18, 'sp4_h_r_45')
// (20, 18, 'sp4_r_v_b_30')
// (20, 18, 'sp4_v_b_29')
// (20, 19, 'sp4_r_v_b_19')
// (20, 19, 'sp4_v_b_16')
// (20, 20, 'local_g2_5')
// (20, 20, 'lutff_0/in_3')
// (20, 20, 'lutff_4/in_1')
// (20, 20, 'lutff_6/in_1')
// (20, 20, 'sp4_h_l_40')
// (20, 20, 'sp4_h_r_25')
// (20, 20, 'sp4_h_r_37')
// (20, 20, 'sp4_r_v_b_6')
// (20, 20, 'sp4_v_b_5')
// (20, 20, 'sp4_v_t_47')
// (20, 21, 'local_g3_7')
// (20, 21, 'lutff_6/in_0')
// (20, 21, 'sp4_h_r_34')
// (20, 21, 'sp4_r_v_b_37')
// (20, 21, 'sp4_v_b_47')
// (20, 22, 'local_g2_2')
// (20, 22, 'lutff_4/in_0')
// (20, 22, 'sp4_h_r_33')
// (20, 22, 'sp4_r_v_b_24')
// (20, 22, 'sp4_v_b_34')
// (20, 23, 'local_g1_7')
// (20, 23, 'lutff_3/in_3')
// (20, 23, 'sp4_r_v_b_13')
// (20, 23, 'sp4_v_b_23')
// (20, 24, 'sp4_r_v_b_0')
// (20, 24, 'sp4_v_b_10')
// (21, 16, 'local_g2_4')
// (21, 16, 'lutff_5/in_3')
// (21, 16, 'sp4_h_r_36')
// (21, 16, 'sp4_v_t_43')
// (21, 17, 'local_g3_3')
// (21, 17, 'lutff_1/in_1')
// (21, 17, 'lutff_6/in_0')
// (21, 17, 'sp4_h_l_40')
// (21, 17, 'sp4_h_r_41')
// (21, 17, 'sp4_r_v_b_36')
// (21, 17, 'sp4_v_b_43')
// (21, 18, 'local_g2_6')
// (21, 18, 'lutff_6/in_0')
// (21, 18, 'sp4_h_l_45')
// (21, 18, 'sp4_h_r_4')
// (21, 18, 'sp4_r_v_b_25')
// (21, 18, 'sp4_v_b_30')
// (21, 19, 'local_g0_3')
// (21, 19, 'lutff_7/in_2')
// (21, 19, 'sp4_r_v_b_12')
// (21, 19, 'sp4_v_b_19')
// (21, 20, 'local_g1_0')
// (21, 20, 'lutff_5/in_0')
// (21, 20, 'sp4_h_l_37')
// (21, 20, 'sp4_h_r_3')
// (21, 20, 'sp4_h_r_36')
// (21, 20, 'sp4_h_r_8')
// (21, 20, 'sp4_r_v_b_1')
// (21, 20, 'sp4_v_b_6')
// (21, 20, 'sp4_v_t_37')
// (21, 21, 'local_g2_5')
// (21, 21, 'lutff_3/in_0')
// (21, 21, 'sp4_h_r_47')
// (21, 21, 'sp4_r_v_b_43')
// (21, 21, 'sp4_v_b_37')
// (21, 22, 'local_g3_0')
// (21, 22, 'lutff_5/in_2')
// (21, 22, 'sp4_h_r_44')
// (21, 22, 'sp4_r_v_b_30')
// (21, 22, 'sp4_v_b_24')
// (21, 23, 'local_g1_5')
// (21, 23, 'lutff_4/in_0')
// (21, 23, 'lutff_7/in_1')
// (21, 23, 'sp4_r_v_b_19')
// (21, 23, 'sp4_v_b_13')
// (21, 24, 'sp4_r_v_b_6')
// (21, 24, 'sp4_v_b_0')
// (22, 16, 'local_g0_1')
// (22, 16, 'local_g1_1')
// (22, 16, 'lutff_4/in_1')
// (22, 16, 'lutff_5/in_0')
// (22, 16, 'lutff_6/in_0')
// (22, 16, 'lutff_7/in_0')
// (22, 16, 'sp4_h_l_36')
// (22, 16, 'sp4_h_r_1')
// (22, 16, 'sp4_v_t_36')
// (22, 17, 'local_g1_4')
// (22, 17, 'lutff_1/in_0')
// (22, 17, 'lutff_3/in_0')
// (22, 17, 'lutff_4/in_3')
// (22, 17, 'lutff_6/in_3')
// (22, 17, 'sp4_h_l_41')
// (22, 17, 'sp4_h_r_4')
// (22, 17, 'sp4_v_b_36')
// (22, 18, 'local_g0_1')
// (22, 18, 'local_g1_1')
// (22, 18, 'lutff_0/in_0')
// (22, 18, 'lutff_1/in_1')
// (22, 18, 'lutff_3/in_2')
// (22, 18, 'sp4_h_r_17')
// (22, 18, 'sp4_v_b_25')
// (22, 19, 'local_g1_4')
// (22, 19, 'lutff_0/in_1')
// (22, 19, 'lutff_4/in_3')
// (22, 19, 'lutff_6/in_3')
// (22, 19, 'sp4_v_b_12')
// (22, 20, 'local_g1_6')
// (22, 20, 'lutff_2/in_1')
// (22, 20, 'lutff_3/in_0')
// (22, 20, 'lutff_4/in_1')
// (22, 20, 'lutff_6/in_3')
// (22, 20, 'lutff_7/in_0')
// (22, 20, 'sp4_h_l_36')
// (22, 20, 'sp4_h_r_14')
// (22, 20, 'sp4_h_r_21')
// (22, 20, 'sp4_v_b_1')
// (22, 20, 'sp4_v_t_43')
// (22, 21, 'local_g0_1')
// (22, 21, 'lutff_7/in_2')
// (22, 21, 'sp4_h_l_47')
// (22, 21, 'sp4_h_r_1')
// (22, 21, 'sp4_v_b_43')
// (22, 22, 'local_g0_0')
// (22, 22, 'local_g1_0')
// (22, 22, 'lutff_3/in_2')
// (22, 22, 'lutff_7/in_1')
// (22, 22, 'sp4_h_l_44')
// (22, 22, 'sp4_h_r_0')
// (22, 22, 'sp4_v_b_30')
// (22, 23, 'local_g1_3')
// (22, 23, 'lutff_1/in_3')
// (22, 23, 'sp4_v_b_19')
// (22, 24, 'sp4_v_b_6')
// (23, 16, 'sp4_h_r_12')
// (23, 17, 'sp4_h_r_17')
// (23, 18, 'sp4_h_r_28')
// (23, 20, 'sp4_h_r_27')
// (23, 20, 'sp4_h_r_32')
// (23, 21, 'sp4_h_r_12')
// (23, 22, 'sp4_h_r_13')
// (24, 16, 'sp4_h_r_25')
// (24, 17, 'sp4_h_r_28')
// (24, 18, 'sp4_h_r_41')
// (24, 20, 'sp4_h_r_38')
// (24, 20, 'sp4_h_r_45')
// (24, 21, 'sp4_h_r_25')
// (24, 22, 'sp4_h_r_24')
// (25, 16, 'sp4_h_r_36')
// (25, 17, 'sp4_h_r_41')
// (25, 18, 'sp4_h_l_41')
// (25, 20, 'sp4_h_l_38')
// (25, 20, 'sp4_h_l_45')
// (25, 21, 'sp4_h_r_36')
// (25, 22, 'sp4_h_r_37')

wire n2298;
// (15, 21, 'sp4_r_v_b_42')
// (15, 22, 'sp4_r_v_b_31')
// (15, 23, 'sp4_r_v_b_18')
// (15, 24, 'sp4_r_v_b_7')
// (16, 19, 'local_g3_6')
// (16, 19, 'lutff_5/in_0')
// (16, 19, 'neigh_op_tnr_6')
// (16, 20, 'local_g2_6')
// (16, 20, 'lutff_6/in_0')
// (16, 20, 'neigh_op_rgt_6')
// (16, 20, 'sp4_h_r_1')
// (16, 20, 'sp4_v_t_42')
// (16, 21, 'local_g1_6')
// (16, 21, 'lutff_7/in_2')
// (16, 21, 'neigh_op_bnr_6')
// (16, 21, 'sp4_v_b_42')
// (16, 22, 'sp4_v_b_31')
// (16, 23, 'sp4_v_b_18')
// (16, 24, 'local_g1_7')
// (16, 24, 'lutff_3/in_1')
// (16, 24, 'sp4_v_b_7')
// (17, 18, 'sp4_r_v_b_37')
// (17, 19, 'neigh_op_top_6')
// (17, 19, 'sp4_r_v_b_24')
// (17, 20, 'lutff_6/out')
// (17, 20, 'sp4_h_r_12')
// (17, 20, 'sp4_r_v_b_13')
// (17, 21, 'neigh_op_bot_6')
// (17, 21, 'sp4_r_v_b_0')
// (17, 22, 'sp4_r_v_b_38')
// (17, 23, 'sp4_r_v_b_27')
// (17, 24, 'local_g2_6')
// (17, 24, 'lutff_7/in_1')
// (17, 24, 'sp4_r_v_b_14')
// (17, 25, 'sp4_r_v_b_3')
// (18, 17, 'sp4_v_t_37')
// (18, 18, 'sp4_v_b_37')
// (18, 19, 'local_g3_6')
// (18, 19, 'lutff_2/in_3')
// (18, 19, 'lutff_7/in_0')
// (18, 19, 'neigh_op_tnl_6')
// (18, 19, 'sp4_v_b_24')
// (18, 20, 'neigh_op_lft_6')
// (18, 20, 'sp4_h_r_25')
// (18, 20, 'sp4_v_b_13')
// (18, 21, 'neigh_op_bnl_6')
// (18, 21, 'sp4_v_b_0')
// (18, 21, 'sp4_v_t_38')
// (18, 22, 'sp4_v_b_38')
// (18, 23, 'sp4_v_b_27')
// (18, 24, 'local_g0_6')
// (18, 24, 'lutff_4/in_0')
// (18, 24, 'sp4_v_b_14')
// (18, 25, 'sp4_v_b_3')
// (19, 20, 'sp4_h_r_36')
// (20, 20, 'sp4_h_l_36')

reg n2299 = 0;
// (15, 22, 'neigh_op_tnr_3')
// (15, 23, 'neigh_op_rgt_3')
// (15, 24, 'neigh_op_bnr_3')
// (16, 22, 'neigh_op_top_3')
// (16, 23, 'lutff_3/out')
// (16, 24, 'neigh_op_bot_3')
// (17, 22, 'local_g3_3')
// (17, 22, 'lutff_5/in_1')
// (17, 22, 'neigh_op_tnl_3')
// (17, 23, 'neigh_op_lft_3')
// (17, 24, 'neigh_op_bnl_3')

wire n2300;
// (15, 22, 'neigh_op_tnr_7')
// (15, 23, 'neigh_op_rgt_7')
// (15, 23, 'sp4_h_r_3')
// (15, 23, 'sp4_h_r_6')
// (15, 24, 'neigh_op_bnr_7')
// (16, 22, 'neigh_op_top_7')
// (16, 23, 'local_g1_3')
// (16, 23, 'lutff_7/out')
// (16, 23, 'lutff_global/cen')
// (16, 23, 'sp4_h_r_14')
// (16, 23, 'sp4_h_r_19')
// (16, 24, 'neigh_op_bot_7')
// (17, 22, 'neigh_op_tnl_7')
// (17, 23, 'neigh_op_lft_7')
// (17, 23, 'sp4_h_r_27')
// (17, 23, 'sp4_h_r_30')
// (17, 24, 'neigh_op_bnl_7')
// (18, 23, 'sp4_h_r_38')
// (18, 23, 'sp4_h_r_43')
// (19, 23, 'sp4_h_l_38')
// (19, 23, 'sp4_h_l_43')
// (19, 23, 'sp4_h_r_3')
// (20, 23, 'sp4_h_r_14')
// (21, 23, 'sp4_h_r_27')
// (22, 23, 'sp4_h_r_38')
// (23, 23, 'sp4_h_l_38')

wire n2301;
// (15, 23, 'neigh_op_tnr_3')
// (15, 24, 'neigh_op_rgt_3')
// (15, 25, 'neigh_op_bnr_3')
// (16, 23, 'neigh_op_top_3')
// (16, 24, 'local_g1_3')
// (16, 24, 'lutff_3/out')
// (16, 24, 'lutff_global/cen')
// (16, 25, 'neigh_op_bot_3')
// (17, 23, 'neigh_op_tnl_3')
// (17, 24, 'neigh_op_lft_3')
// (17, 25, 'neigh_op_bnl_3')

reg n2302 = 0;
// (15, 23, 'neigh_op_tnr_7')
// (15, 23, 'sp4_r_v_b_43')
// (15, 24, 'neigh_op_rgt_7')
// (15, 24, 'sp4_r_v_b_30')
// (15, 25, 'neigh_op_bnr_7')
// (15, 25, 'sp4_r_v_b_19')
// (15, 26, 'sp4_r_v_b_6')
// (16, 22, 'sp4_h_r_11')
// (16, 22, 'sp4_v_t_43')
// (16, 23, 'neigh_op_top_7')
// (16, 23, 'sp4_v_b_43')
// (16, 24, 'lutff_7/out')
// (16, 24, 'sp4_v_b_30')
// (16, 25, 'neigh_op_bot_7')
// (16, 25, 'sp4_v_b_19')
// (16, 26, 'sp4_v_b_6')
// (17, 22, 'sp4_h_r_22')
// (17, 23, 'neigh_op_tnl_7')
// (17, 24, 'neigh_op_lft_7')
// (17, 25, 'neigh_op_bnl_7')
// (18, 22, 'local_g3_3')
// (18, 22, 'lutff_1/in_1')
// (18, 22, 'sp4_h_r_35')
// (19, 22, 'sp4_h_r_46')
// (20, 22, 'sp4_h_l_46')

wire n2303;
// (16, 0, 'logic_op_tnr_1')
// (16, 1, 'neigh_op_rgt_1')
// (16, 2, 'neigh_op_bnr_1')
// (16, 2, 'sp4_r_v_b_45')
// (16, 3, 'sp4_r_v_b_32')
// (16, 4, 'local_g3_5')
// (16, 4, 'lutff_2/in_2')
// (16, 4, 'lutff_3/in_1')
// (16, 4, 'lutff_5/in_1')
// (16, 4, 'lutff_7/in_3')
// (16, 4, 'sp4_r_v_b_21')
// (16, 5, 'sp4_r_v_b_8')
// (17, 0, 'logic_op_top_1')
// (17, 1, 'lutff_1/out')
// (17, 1, 'sp4_h_r_2')
// (17, 1, 'sp4_v_t_45')
// (17, 2, 'neigh_op_bot_1')
// (17, 2, 'sp4_v_b_45')
// (17, 3, 'sp4_v_b_32')
// (17, 4, 'sp4_v_b_21')
// (17, 5, 'sp4_v_b_8')
// (18, 0, 'logic_op_tnl_1')
// (18, 1, 'neigh_op_lft_1')
// (18, 1, 'sp4_h_r_15')
// (18, 2, 'neigh_op_bnl_1')
// (19, 1, 'sp4_h_r_26')
// (20, 1, 'sp4_h_r_39')
// (21, 1, 'sp4_h_l_39')

wire n2304;
// (16, 0, 'logic_op_tnr_2')
// (16, 1, 'neigh_op_rgt_2')
// (16, 1, 'sp4_r_v_b_36')
// (16, 2, 'neigh_op_bnr_2')
// (16, 2, 'sp4_r_v_b_25')
// (16, 3, 'sp4_r_v_b_12')
// (16, 4, 'sp4_r_v_b_1')
// (17, 0, 'logic_op_top_2')
// (17, 0, 'span4_vert_36')
// (17, 1, 'lutff_2/out')
// (17, 1, 'sp4_v_b_36')
// (17, 2, 'local_g1_2')
// (17, 2, 'lutff_2/in_3')
// (17, 2, 'neigh_op_bot_2')
// (17, 2, 'sp4_v_b_25')
// (17, 3, 'local_g0_4')
// (17, 3, 'lutff_0/in_2')
// (17, 3, 'lutff_4/in_0')
// (17, 3, 'lutff_6/in_2')
// (17, 3, 'sp4_v_b_12')
// (17, 4, 'sp4_v_b_1')
// (18, 0, 'logic_op_tnl_2')
// (18, 1, 'neigh_op_lft_2')
// (18, 2, 'neigh_op_bnl_2')

wire n2305;
// (16, 0, 'logic_op_tnr_3')
// (16, 1, 'neigh_op_rgt_3')
// (16, 2, 'neigh_op_bnr_3')
// (17, 0, 'logic_op_top_3')
// (17, 1, 'lutff_3/out')
// (17, 1, 'sp4_r_v_b_39')
// (17, 2, 'local_g0_3')
// (17, 2, 'lutff_1/in_2')
// (17, 2, 'lutff_7/in_0')
// (17, 2, 'neigh_op_bot_3')
// (17, 2, 'sp4_r_v_b_26')
// (17, 3, 'local_g2_7')
// (17, 3, 'lutff_3/in_2')
// (17, 3, 'lutff_7/in_2')
// (17, 3, 'sp4_r_v_b_15')
// (17, 4, 'sp4_r_v_b_2')
// (18, 0, 'logic_op_tnl_3')
// (18, 0, 'span4_vert_39')
// (18, 1, 'neigh_op_lft_3')
// (18, 1, 'sp4_v_b_39')
// (18, 2, 'neigh_op_bnl_3')
// (18, 2, 'sp4_v_b_26')
// (18, 3, 'sp4_v_b_15')
// (18, 4, 'sp4_v_b_2')

reg n2306 = 0;
// (16, 1, 'neigh_op_tnr_1')
// (16, 2, 'neigh_op_rgt_1')
// (16, 3, 'neigh_op_bnr_1')
// (17, 1, 'neigh_op_top_1')
// (17, 2, 'local_g3_1')
// (17, 2, 'lutff_1/out')
// (17, 2, 'lutff_6/in_0')
// (17, 3, 'neigh_op_bot_1')
// (18, 1, 'neigh_op_tnl_1')
// (18, 2, 'neigh_op_lft_1')
// (18, 3, 'neigh_op_bnl_1')

reg n2307 = 0;
// (16, 1, 'neigh_op_tnr_2')
// (16, 2, 'neigh_op_rgt_2')
// (16, 3, 'neigh_op_bnr_2')
// (17, 1, 'neigh_op_top_2')
// (17, 2, 'local_g2_2')
// (17, 2, 'lutff_0/in_2')
// (17, 2, 'lutff_2/out')
// (17, 3, 'neigh_op_bot_2')
// (18, 1, 'neigh_op_tnl_2')
// (18, 2, 'neigh_op_lft_2')
// (18, 3, 'neigh_op_bnl_2')

reg n2308 = 0;
// (16, 1, 'neigh_op_tnr_3')
// (16, 2, 'neigh_op_rgt_3')
// (16, 3, 'neigh_op_bnr_3')
// (17, 1, 'neigh_op_top_3')
// (17, 2, 'local_g3_3')
// (17, 2, 'lutff_3/out')
// (17, 2, 'lutff_5/in_1')
// (17, 3, 'neigh_op_bot_3')
// (18, 1, 'neigh_op_tnl_3')
// (18, 2, 'neigh_op_lft_3')
// (18, 3, 'neigh_op_bnl_3')

reg n2309 = 0;
// (16, 1, 'neigh_op_tnr_4')
// (16, 2, 'neigh_op_rgt_4')
// (16, 3, 'neigh_op_bnr_4')
// (17, 1, 'neigh_op_top_4')
// (17, 2, 'local_g1_4')
// (17, 2, 'lutff_4/out')
// (17, 2, 'lutff_5/in_2')
// (17, 3, 'neigh_op_bot_4')
// (18, 1, 'neigh_op_tnl_4')
// (18, 2, 'neigh_op_lft_4')
// (18, 3, 'neigh_op_bnl_4')

wire n2310;
// (16, 1, 'neigh_op_tnr_5')
// (16, 2, 'neigh_op_rgt_5')
// (16, 3, 'neigh_op_bnr_5')
// (17, 1, 'neigh_op_top_5')
// (17, 1, 'sp4_r_v_b_38')
// (17, 2, 'local_g1_5')
// (17, 2, 'lutff_4/in_0')
// (17, 2, 'lutff_5/out')
// (17, 2, 'sp4_r_v_b_27')
// (17, 3, 'neigh_op_bot_5')
// (17, 3, 'sp4_r_v_b_14')
// (17, 4, 'local_g1_3')
// (17, 4, 'lutff_6/in_0')
// (17, 4, 'sp4_r_v_b_3')
// (18, 0, 'span4_vert_38')
// (18, 1, 'neigh_op_tnl_5')
// (18, 1, 'sp4_v_b_38')
// (18, 2, 'local_g0_5')
// (18, 2, 'lutff_5/in_2')
// (18, 2, 'neigh_op_lft_5')
// (18, 2, 'sp4_v_b_27')
// (18, 3, 'neigh_op_bnl_5')
// (18, 3, 'sp4_v_b_14')
// (18, 4, 'local_g1_3')
// (18, 4, 'lutff_2/in_0')
// (18, 4, 'sp4_v_b_3')

wire n2311;
// (16, 1, 'neigh_op_tnr_6')
// (16, 2, 'neigh_op_rgt_6')
// (16, 3, 'neigh_op_bnr_6')
// (17, 1, 'neigh_op_top_6')
// (17, 1, 'sp4_r_v_b_40')
// (17, 2, 'local_g1_6')
// (17, 2, 'lutff_1/in_0')
// (17, 2, 'lutff_6/out')
// (17, 2, 'sp4_r_v_b_29')
// (17, 3, 'neigh_op_bot_6')
// (17, 3, 'sp4_r_v_b_16')
// (17, 4, 'local_g1_5')
// (17, 4, 'lutff_2/in_2')
// (17, 4, 'sp4_r_v_b_5')
// (18, 0, 'span4_vert_40')
// (18, 1, 'neigh_op_tnl_6')
// (18, 1, 'sp4_v_b_40')
// (18, 2, 'local_g1_6')
// (18, 2, 'lutff_6/in_3')
// (18, 2, 'neigh_op_lft_6')
// (18, 2, 'sp4_v_b_29')
// (18, 3, 'neigh_op_bnl_6')
// (18, 3, 'sp4_v_b_16')
// (18, 4, 'local_g0_5')
// (18, 4, 'lutff_3/in_0')
// (18, 4, 'sp4_v_b_5')

reg n2312 = 0;
// (16, 1, 'neigh_op_tnr_7')
// (16, 2, 'neigh_op_rgt_7')
// (16, 3, 'neigh_op_bnr_7')
// (17, 1, 'neigh_op_top_7')
// (17, 2, 'local_g1_7')
// (17, 2, 'lutff_6/in_2')
// (17, 2, 'lutff_7/out')
// (17, 3, 'neigh_op_bot_7')
// (18, 1, 'neigh_op_tnl_7')
// (18, 2, 'neigh_op_lft_7')
// (18, 3, 'neigh_op_bnl_7')

wire n2313;
// (16, 1, 'sp4_h_r_2')
// (17, 0, 'logic_op_tnr_5')
// (17, 1, 'neigh_op_rgt_5')
// (17, 1, 'sp4_h_r_15')
// (17, 2, 'local_g0_5')
// (17, 2, 'lutff_3/in_2')
// (17, 2, 'lutff_4/in_1')
// (17, 2, 'neigh_op_bnr_5')
// (18, 0, 'logic_op_top_5')
// (18, 1, 'lutff_5/out')
// (18, 1, 'sp4_h_r_26')
// (18, 2, 'neigh_op_bot_5')
// (19, 0, 'logic_op_tnl_5')
// (19, 1, 'neigh_op_lft_5')
// (19, 1, 'sp4_h_r_39')
// (19, 2, 'neigh_op_bnl_5')
// (19, 2, 'sp4_r_v_b_42')
// (19, 3, 'sp4_r_v_b_31')
// (19, 4, 'sp4_r_v_b_18')
// (19, 5, 'sp4_r_v_b_7')
// (20, 1, 'sp4_h_l_39')
// (20, 1, 'sp4_v_t_42')
// (20, 2, 'local_g2_2')
// (20, 2, 'lutff_0/in_0')
// (20, 2, 'lutff_6/in_0')
// (20, 2, 'sp4_v_b_42')
// (20, 3, 'sp4_v_b_31')
// (20, 4, 'sp4_v_b_18')
// (20, 5, 'sp4_v_b_7')

reg n2314 = 0;
// (16, 1, 'sp4_h_r_3')
// (17, 1, 'local_g0_6')
// (17, 1, 'lutff_1/in_3')
// (17, 1, 'lutff_2/in_2')
// (17, 1, 'lutff_3/in_1')
// (17, 1, 'sp4_h_r_10')
// (17, 1, 'sp4_h_r_14')
// (18, 1, 'local_g0_7')
// (18, 1, 'local_g1_7')
// (18, 1, 'lutff_0/in_1')
// (18, 1, 'lutff_1/in_3')
// (18, 1, 'lutff_5/in_2')
// (18, 1, 'sp4_h_r_23')
// (18, 1, 'sp4_h_r_27')
// (19, 1, 'sp4_h_r_34')
// (19, 1, 'sp4_h_r_38')
// (20, 0, 'logic_op_tnr_1')
// (20, 1, 'local_g2_1')
// (20, 1, 'lutff_0/in_1')
// (20, 1, 'lutff_4/in_3')
// (20, 1, 'neigh_op_rgt_1')
// (20, 1, 'sp4_h_l_38')
// (20, 1, 'sp4_h_r_47')
// (20, 1, 'sp4_h_r_7')
// (20, 2, 'neigh_op_bnr_1')
// (21, 0, 'logic_op_top_1')
// (21, 1, 'local_g0_1')
// (21, 1, 'local_g2_1')
// (21, 1, 'lutff_0/in_3')
// (21, 1, 'lutff_1/in_2')
// (21, 1, 'lutff_1/out')
// (21, 1, 'lutff_5/in_2')
// (21, 1, 'sp4_h_l_47')
// (21, 1, 'sp4_h_r_18')
// (21, 1, 'sp4_h_r_2')
// (21, 2, 'neigh_op_bot_1')
// (22, 0, 'logic_op_tnl_1')
// (22, 1, 'neigh_op_lft_1')
// (22, 1, 'sp4_h_r_15')
// (22, 1, 'sp4_h_r_31')
// (22, 2, 'neigh_op_bnl_1')
// (23, 1, 'sp4_h_r_26')
// (23, 1, 'sp4_h_r_42')
// (24, 1, 'sp4_h_l_42')
// (24, 1, 'sp4_h_r_39')
// (25, 1, 'sp4_h_l_39')

reg n2315 = 0;
// (16, 1, 'sp4_r_v_b_34')
// (16, 2, 'sp4_r_v_b_23')
// (16, 3, 'local_g2_2')
// (16, 3, 'lutff_1/in_3')
// (16, 3, 'sp4_r_v_b_10')
// (16, 4, 'sp4_r_v_b_47')
// (16, 5, 'local_g0_1')
// (16, 5, 'lutff_4/in_1')
// (16, 5, 'sp4_r_v_b_34')
// (16, 6, 'neigh_op_tnr_5')
// (16, 6, 'sp4_r_v_b_23')
// (16, 7, 'neigh_op_rgt_5')
// (16, 7, 'sp4_r_v_b_10')
// (16, 8, 'neigh_op_bnr_5')
// (17, 0, 'span4_vert_34')
// (17, 1, 'sp4_v_b_34')
// (17, 2, 'sp4_v_b_23')
// (17, 3, 'sp4_v_b_10')
// (17, 3, 'sp4_v_t_47')
// (17, 4, 'sp4_v_b_47')
// (17, 5, 'sp4_v_b_34')
// (17, 6, 'neigh_op_top_5')
// (17, 6, 'sp4_v_b_23')
// (17, 7, 'local_g3_5')
// (17, 7, 'lutff_5/in_1')
// (17, 7, 'lutff_5/out')
// (17, 7, 'sp4_v_b_10')
// (17, 8, 'neigh_op_bot_5')
// (18, 6, 'neigh_op_tnl_5')
// (18, 7, 'neigh_op_lft_5')
// (18, 8, 'neigh_op_bnl_5')

wire n2316;
// (16, 1, 'sp4_r_v_b_47')
// (16, 2, 'sp4_r_v_b_34')
// (16, 3, 'sp4_r_v_b_23')
// (16, 4, 'sp4_r_v_b_10')
// (17, 0, 'span4_vert_47')
// (17, 1, 'sp4_v_b_47')
// (17, 2, 'sp4_v_b_34')
// (17, 3, 'sp4_v_b_23')
// (17, 4, 'local_g0_2')
// (17, 4, 'lutff_global/cen')
// (17, 4, 'sp4_h_r_5')
// (17, 4, 'sp4_v_b_10')
// (18, 4, 'sp4_h_r_16')
// (19, 3, 'neigh_op_tnr_4')
// (19, 4, 'neigh_op_rgt_4')
// (19, 4, 'sp4_h_r_29')
// (19, 5, 'neigh_op_bnr_4')
// (20, 3, 'neigh_op_top_4')
// (20, 4, 'lutff_4/out')
// (20, 4, 'sp4_h_r_40')
// (20, 5, 'neigh_op_bot_4')
// (21, 3, 'neigh_op_tnl_4')
// (21, 4, 'neigh_op_lft_4')
// (21, 4, 'sp4_h_l_40')
// (21, 5, 'neigh_op_bnl_4')

reg n2317 = 0;
// (16, 2, 'neigh_op_tnr_0')
// (16, 3, 'neigh_op_rgt_0')
// (16, 4, 'neigh_op_bnr_0')
// (17, 2, 'neigh_op_top_0')
// (17, 3, 'local_g0_0')
// (17, 3, 'lutff_0/out')
// (17, 3, 'lutff_5/in_1')
// (17, 4, 'neigh_op_bot_0')
// (18, 2, 'neigh_op_tnl_0')
// (18, 3, 'neigh_op_lft_0')
// (18, 4, 'neigh_op_bnl_0')

wire n2318;
// (16, 2, 'neigh_op_tnr_1')
// (16, 3, 'neigh_op_rgt_1')
// (16, 4, 'neigh_op_bnr_1')
// (17, 2, 'neigh_op_top_1')
// (17, 2, 'sp4_r_v_b_46')
// (17, 3, 'local_g3_1')
// (17, 3, 'lutff_1/out')
// (17, 3, 'lutff_3/in_3')
// (17, 3, 'sp4_r_v_b_35')
// (17, 4, 'local_g0_1')
// (17, 4, 'lutff_5/in_0')
// (17, 4, 'neigh_op_bot_1')
// (17, 4, 'sp4_r_v_b_22')
// (17, 5, 'sp4_r_v_b_11')
// (18, 1, 'sp4_v_t_46')
// (18, 2, 'neigh_op_tnl_1')
// (18, 2, 'sp4_v_b_46')
// (18, 3, 'neigh_op_lft_1')
// (18, 3, 'sp4_v_b_35')
// (18, 4, 'neigh_op_bnl_1')
// (18, 4, 'sp4_v_b_22')
// (18, 5, 'local_g1_3')
// (18, 5, 'lutff_3/in_3')
// (18, 5, 'sp4_v_b_11')

reg n2319 = 0;
// (16, 2, 'neigh_op_tnr_3')
// (16, 3, 'neigh_op_rgt_3')
// (16, 4, 'neigh_op_bnr_3')
// (17, 2, 'neigh_op_top_3')
// (17, 3, 'local_g3_3')
// (17, 3, 'lutff_1/in_3')
// (17, 3, 'lutff_3/out')
// (17, 4, 'neigh_op_bot_3')
// (18, 2, 'neigh_op_tnl_3')
// (18, 3, 'neigh_op_lft_3')
// (18, 4, 'neigh_op_bnl_3')

reg n2320 = 0;
// (16, 2, 'neigh_op_tnr_4')
// (16, 3, 'neigh_op_rgt_4')
// (16, 4, 'neigh_op_bnr_4')
// (17, 2, 'local_g0_4')
// (17, 2, 'lutff_0/in_0')
// (17, 2, 'neigh_op_top_4')
// (17, 3, 'lutff_4/out')
// (17, 4, 'neigh_op_bot_4')
// (18, 2, 'neigh_op_tnl_4')
// (18, 3, 'neigh_op_lft_4')
// (18, 4, 'neigh_op_bnl_4')

wire n2321;
// (16, 2, 'neigh_op_tnr_5')
// (16, 3, 'neigh_op_rgt_5')
// (16, 4, 'neigh_op_bnr_5')
// (17, 2, 'neigh_op_top_5')
// (17, 3, 'local_g0_5')
// (17, 3, 'lutff_0/in_1')
// (17, 3, 'lutff_5/out')
// (17, 4, 'local_g0_5')
// (17, 4, 'lutff_7/in_2')
// (17, 4, 'neigh_op_bot_5')
// (18, 2, 'local_g2_5')
// (18, 2, 'lutff_3/in_0')
// (18, 2, 'neigh_op_tnl_5')
// (18, 3, 'neigh_op_lft_5')
// (18, 4, 'local_g2_5')
// (18, 4, 'lutff_1/in_0')
// (18, 4, 'neigh_op_bnl_5')

reg n2322 = 0;
// (16, 2, 'neigh_op_tnr_6')
// (16, 3, 'neigh_op_rgt_6')
// (16, 4, 'neigh_op_bnr_6')
// (17, 2, 'neigh_op_top_6')
// (17, 3, 'local_g1_6')
// (17, 3, 'lutff_5/in_0')
// (17, 3, 'lutff_6/out')
// (17, 4, 'neigh_op_bot_6')
// (18, 2, 'neigh_op_tnl_6')
// (18, 3, 'neigh_op_lft_6')
// (18, 4, 'neigh_op_bnl_6')

reg n2323 = 0;
// (16, 2, 'neigh_op_tnr_7')
// (16, 3, 'neigh_op_rgt_7')
// (16, 4, 'neigh_op_bnr_7')
// (17, 2, 'neigh_op_top_7')
// (17, 3, 'local_g0_7')
// (17, 3, 'lutff_1/in_2')
// (17, 3, 'lutff_7/out')
// (17, 4, 'neigh_op_bot_7')
// (18, 2, 'neigh_op_tnl_7')
// (18, 3, 'neigh_op_lft_7')
// (18, 4, 'neigh_op_bnl_7')

wire n2324;
// (16, 2, 'sp4_h_r_7')
// (16, 3, 'sp4_r_v_b_39')
// (16, 4, 'local_g0_2')
// (16, 4, 'lutff_global/cen')
// (16, 4, 'sp4_r_v_b_26')
// (16, 5, 'sp4_r_v_b_15')
// (16, 6, 'sp4_r_v_b_2')
// (17, 2, 'local_g0_2')
// (17, 2, 'lutff_global/cen')
// (17, 2, 'sp4_h_r_18')
// (17, 2, 'sp4_h_r_2')
// (17, 2, 'sp4_v_t_39')
// (17, 3, 'local_g1_3')
// (17, 3, 'lutff_global/cen')
// (17, 3, 'sp4_h_r_11')
// (17, 3, 'sp4_v_b_39')
// (17, 4, 'sp4_v_b_26')
// (17, 5, 'sp4_v_b_15')
// (17, 6, 'sp4_v_b_2')
// (18, 2, 'sp4_h_r_15')
// (18, 2, 'sp4_h_r_31')
// (18, 3, 'sp4_h_r_22')
// (19, 2, 'sp4_h_r_26')
// (19, 2, 'sp4_h_r_42')
// (19, 3, 'sp4_h_r_35')
// (20, 1, 'neigh_op_tnr_3')
// (20, 1, 'sp4_r_v_b_35')
// (20, 2, 'local_g3_3')
// (20, 2, 'lutff_global/cen')
// (20, 2, 'neigh_op_rgt_3')
// (20, 2, 'sp4_h_l_42')
// (20, 2, 'sp4_h_r_11')
// (20, 2, 'sp4_h_r_39')
// (20, 2, 'sp4_r_v_b_22')
// (20, 3, 'neigh_op_bnr_3')
// (20, 3, 'sp4_h_r_46')
// (20, 3, 'sp4_r_v_b_11')
// (21, 0, 'span4_vert_35')
// (21, 1, 'neigh_op_top_3')
// (21, 1, 'sp4_v_b_35')
// (21, 2, 'lutff_3/out')
// (21, 2, 'sp4_h_l_39')
// (21, 2, 'sp4_h_r_22')
// (21, 2, 'sp4_h_r_6')
// (21, 2, 'sp4_v_b_22')
// (21, 3, 'neigh_op_bot_3')
// (21, 3, 'sp4_h_l_46')
// (21, 3, 'sp4_v_b_11')
// (22, 1, 'neigh_op_tnl_3')
// (22, 2, 'local_g1_3')
// (22, 2, 'lutff_0/in_2')
// (22, 2, 'neigh_op_lft_3')
// (22, 2, 'sp4_h_r_19')
// (22, 2, 'sp4_h_r_35')
// (22, 3, 'neigh_op_bnl_3')
// (23, 2, 'sp4_h_r_30')
// (23, 2, 'sp4_h_r_46')
// (24, 2, 'sp4_h_l_46')
// (24, 2, 'sp4_h_r_43')
// (25, 2, 'sp4_h_l_43')

reg n2325 = 0;
// (16, 3, 'neigh_op_tnr_0')
// (16, 4, 'neigh_op_rgt_0')
// (16, 5, 'neigh_op_bnr_0')
// (17, 3, 'neigh_op_top_0')
// (17, 4, 'lutff_0/out')
// (17, 5, 'local_g0_0')
// (17, 5, 'lutff_4/in_0')
// (17, 5, 'neigh_op_bot_0')
// (18, 3, 'neigh_op_tnl_0')
// (18, 4, 'neigh_op_lft_0')
// (18, 5, 'neigh_op_bnl_0')

reg n2326 = 0;
// (16, 3, 'neigh_op_tnr_1')
// (16, 4, 'neigh_op_rgt_1')
// (16, 5, 'neigh_op_bnr_1')
// (17, 3, 'neigh_op_top_1')
// (17, 4, 'lutff_1/out')
// (17, 5, 'local_g1_1')
// (17, 5, 'lutff_3/in_1')
// (17, 5, 'neigh_op_bot_1')
// (18, 3, 'neigh_op_tnl_1')
// (18, 4, 'neigh_op_lft_1')
// (18, 5, 'neigh_op_bnl_1')

reg n2327 = 0;
// (16, 3, 'neigh_op_tnr_2')
// (16, 4, 'neigh_op_rgt_2')
// (16, 5, 'neigh_op_bnr_2')
// (17, 2, 'sp4_r_v_b_45')
// (17, 3, 'neigh_op_top_2')
// (17, 3, 'sp4_r_v_b_32')
// (17, 4, 'lutff_2/out')
// (17, 4, 'sp4_r_v_b_21')
// (17, 5, 'neigh_op_bot_2')
// (17, 5, 'sp4_r_v_b_8')
// (18, 1, 'sp4_v_t_45')
// (18, 2, 'local_g3_5')
// (18, 2, 'lutff_0/in_2')
// (18, 2, 'sp4_v_b_45')
// (18, 3, 'neigh_op_tnl_2')
// (18, 3, 'sp4_v_b_32')
// (18, 4, 'neigh_op_lft_2')
// (18, 4, 'sp4_v_b_21')
// (18, 5, 'neigh_op_bnl_2')
// (18, 5, 'sp4_v_b_8')

reg n2328 = 0;
// (16, 3, 'neigh_op_tnr_3')
// (16, 4, 'neigh_op_rgt_3')
// (16, 5, 'neigh_op_bnr_3')
// (17, 3, 'neigh_op_top_3')
// (17, 4, 'lutff_3/out')
// (17, 5, 'local_g0_3')
// (17, 5, 'lutff_7/in_0')
// (17, 5, 'neigh_op_bot_3')
// (18, 3, 'neigh_op_tnl_3')
// (18, 4, 'neigh_op_lft_3')
// (18, 5, 'neigh_op_bnl_3')

reg n2329 = 0;
// (16, 3, 'neigh_op_tnr_4')
// (16, 4, 'neigh_op_rgt_4')
// (16, 5, 'neigh_op_bnr_4')
// (17, 3, 'neigh_op_top_4')
// (17, 4, 'lutff_4/out')
// (17, 5, 'local_g1_4')
// (17, 5, 'lutff_1/in_2')
// (17, 5, 'neigh_op_bot_4')
// (18, 3, 'neigh_op_tnl_4')
// (18, 4, 'neigh_op_lft_4')
// (18, 5, 'neigh_op_bnl_4')

reg n2330 = 0;
// (16, 3, 'neigh_op_tnr_5')
// (16, 4, 'neigh_op_rgt_5')
// (16, 5, 'neigh_op_bnr_5')
// (17, 3, 'neigh_op_top_5')
// (17, 4, 'lutff_5/out')
// (17, 5, 'local_g0_5')
// (17, 5, 'lutff_2/in_3')
// (17, 5, 'neigh_op_bot_5')
// (18, 3, 'neigh_op_tnl_5')
// (18, 4, 'neigh_op_lft_5')
// (18, 5, 'neigh_op_bnl_5')

reg n2331 = 0;
// (16, 3, 'neigh_op_tnr_6')
// (16, 4, 'neigh_op_rgt_6')
// (16, 5, 'neigh_op_bnr_6')
// (17, 3, 'neigh_op_top_6')
// (17, 4, 'lutff_6/out')
// (17, 5, 'local_g1_6')
// (17, 5, 'lutff_0/in_3')
// (17, 5, 'neigh_op_bot_6')
// (18, 3, 'neigh_op_tnl_6')
// (18, 4, 'neigh_op_lft_6')
// (18, 5, 'neigh_op_bnl_6')

reg n2332 = 0;
// (16, 3, 'neigh_op_tnr_7')
// (16, 4, 'neigh_op_rgt_7')
// (16, 5, 'neigh_op_bnr_7')
// (17, 3, 'neigh_op_top_7')
// (17, 4, 'lutff_7/out')
// (17, 5, 'neigh_op_bot_7')
// (18, 3, 'neigh_op_tnl_7')
// (18, 4, 'neigh_op_lft_7')
// (18, 5, 'local_g3_7')
// (18, 5, 'lutff_1/in_1')
// (18, 5, 'neigh_op_bnl_7')

wire n2333;
// (16, 3, 'sp4_r_v_b_38')
// (16, 4, 'local_g1_3')
// (16, 4, 'lutff_2/in_0')
// (16, 4, 'lutff_5/in_3')
// (16, 4, 'sp4_r_v_b_27')
// (16, 5, 'sp4_r_v_b_14')
// (16, 6, 'sp4_r_v_b_3')
// (17, 1, 'neigh_op_tnr_2')
// (17, 2, 'local_g3_2')
// (17, 2, 'lutff_2/in_1')
// (17, 2, 'neigh_op_rgt_2')
// (17, 2, 'sp4_h_r_9')
// (17, 2, 'sp4_v_t_38')
// (17, 3, 'local_g0_2')
// (17, 3, 'lutff_3/in_1')
// (17, 3, 'lutff_4/in_2')
// (17, 3, 'lutff_7/in_1')
// (17, 3, 'neigh_op_bnr_2')
// (17, 3, 'sp4_v_b_38')
// (17, 4, 'sp4_v_b_27')
// (17, 5, 'sp4_v_b_14')
// (17, 6, 'sp4_v_b_3')
// (18, 1, 'neigh_op_top_2')
// (18, 2, 'lutff_2/out')
// (18, 2, 'sp4_h_r_20')
// (18, 2, 'sp4_h_r_4')
// (18, 3, 'neigh_op_bot_2')
// (19, 1, 'neigh_op_tnl_2')
// (19, 2, 'neigh_op_lft_2')
// (19, 2, 'sp4_h_r_17')
// (19, 2, 'sp4_h_r_33')
// (19, 3, 'neigh_op_bnl_2')
// (20, 2, 'local_g2_4')
// (20, 2, 'lutff_0/in_2')
// (20, 2, 'lutff_6/in_2')
// (20, 2, 'sp4_h_r_28')
// (20, 2, 'sp4_h_r_44')
// (21, 2, 'sp4_h_l_44')
// (21, 2, 'sp4_h_r_41')
// (22, 2, 'sp4_h_l_41')

reg n2334 = 0;
// (16, 4, 'neigh_op_tnr_0')
// (16, 5, 'neigh_op_rgt_0')
// (16, 5, 'sp4_h_r_5')
// (16, 6, 'neigh_op_bnr_0')
// (17, 4, 'neigh_op_top_0')
// (17, 5, 'lutff_0/out')
// (17, 5, 'sp4_h_r_16')
// (17, 6, 'neigh_op_bot_0')
// (18, 4, 'neigh_op_tnl_0')
// (18, 5, 'neigh_op_lft_0')
// (18, 5, 'sp4_h_r_29')
// (18, 6, 'neigh_op_bnl_0')
// (19, 5, 'local_g2_0')
// (19, 5, 'ram/WDATA_10')
// (19, 5, 'sp4_h_r_40')
// (20, 5, 'sp4_h_l_40')

reg n2335 = 0;
// (16, 4, 'neigh_op_tnr_1')
// (16, 5, 'neigh_op_rgt_1')
// (16, 6, 'neigh_op_bnr_1')
// (17, 4, 'neigh_op_top_1')
// (17, 5, 'lutff_1/out')
// (17, 5, 'sp4_h_r_2')
// (17, 6, 'neigh_op_bot_1')
// (18, 4, 'neigh_op_tnl_1')
// (18, 5, 'neigh_op_lft_1')
// (18, 5, 'sp4_h_r_15')
// (18, 6, 'neigh_op_bnl_1')
// (19, 5, 'local_g2_2')
// (19, 5, 'ram/WDATA_14')
// (19, 5, 'sp4_h_r_26')
// (20, 5, 'sp4_h_r_39')
// (21, 5, 'sp4_h_l_39')

reg n2336 = 0;
// (16, 4, 'neigh_op_tnr_2')
// (16, 5, 'neigh_op_rgt_2')
// (16, 5, 'sp4_h_r_9')
// (16, 6, 'neigh_op_bnr_2')
// (17, 4, 'neigh_op_top_2')
// (17, 5, 'lutff_2/out')
// (17, 5, 'sp4_h_r_20')
// (17, 6, 'neigh_op_bot_2')
// (18, 4, 'neigh_op_tnl_2')
// (18, 5, 'neigh_op_lft_2')
// (18, 5, 'sp4_h_r_33')
// (18, 6, 'neigh_op_bnl_2')
// (19, 5, 'local_g2_4')
// (19, 5, 'ram/WDATA_12')
// (19, 5, 'sp4_h_r_44')
// (20, 5, 'sp4_h_l_44')

reg n2337 = 0;
// (16, 4, 'neigh_op_tnr_3')
// (16, 5, 'neigh_op_rgt_3')
// (16, 6, 'neigh_op_bnr_3')
// (17, 2, 'sp4_r_v_b_42')
// (17, 3, 'sp4_r_v_b_31')
// (17, 4, 'neigh_op_top_3')
// (17, 4, 'sp4_r_v_b_18')
// (17, 5, 'lutff_3/out')
// (17, 5, 'sp4_r_v_b_7')
// (17, 6, 'neigh_op_bot_3')
// (18, 1, 'sp4_v_t_42')
// (18, 2, 'sp4_v_b_42')
// (18, 3, 'sp4_v_b_31')
// (18, 4, 'neigh_op_tnl_3')
// (18, 4, 'sp4_v_b_18')
// (18, 5, 'neigh_op_lft_3')
// (18, 5, 'sp4_h_r_1')
// (18, 5, 'sp4_v_b_7')
// (18, 6, 'neigh_op_bnl_3')
// (19, 5, 'local_g1_4')
// (19, 5, 'ram/WDATA_13')
// (19, 5, 'sp4_h_r_12')
// (20, 5, 'sp4_h_r_25')
// (21, 5, 'sp4_h_r_36')
// (22, 5, 'sp4_h_l_36')

reg n2338 = 0;
// (16, 4, 'neigh_op_tnr_4')
// (16, 5, 'neigh_op_rgt_4')
// (16, 6, 'neigh_op_bnr_4')
// (17, 4, 'neigh_op_top_4')
// (17, 5, 'lutff_4/out')
// (17, 5, 'sp4_h_r_8')
// (17, 6, 'neigh_op_bot_4')
// (18, 4, 'neigh_op_tnl_4')
// (18, 5, 'neigh_op_lft_4')
// (18, 5, 'sp4_h_r_21')
// (18, 6, 'neigh_op_bnl_4')
// (19, 5, 'local_g3_0')
// (19, 5, 'ram/WDATA_11')
// (19, 5, 'sp4_h_r_32')
// (20, 5, 'sp4_h_r_45')
// (21, 5, 'sp4_h_l_45')

reg n2339 = 0;
// (16, 4, 'neigh_op_tnr_6')
// (16, 5, 'neigh_op_rgt_6')
// (16, 6, 'neigh_op_bnr_6')
// (17, 3, 'sp4_r_v_b_37')
// (17, 4, 'neigh_op_top_6')
// (17, 4, 'sp4_r_v_b_24')
// (17, 5, 'lutff_6/out')
// (17, 5, 'sp4_r_v_b_13')
// (17, 6, 'neigh_op_bot_6')
// (17, 6, 'sp4_r_v_b_0')
// (18, 2, 'sp4_v_t_37')
// (18, 3, 'sp4_v_b_37')
// (18, 4, 'neigh_op_tnl_6')
// (18, 4, 'sp4_v_b_24')
// (18, 5, 'neigh_op_lft_6')
// (18, 5, 'sp4_v_b_13')
// (18, 6, 'neigh_op_bnl_6')
// (18, 6, 'sp4_h_r_0')
// (18, 6, 'sp4_v_b_0')
// (19, 6, 'local_g0_5')
// (19, 6, 'ram/WDATA_7')
// (19, 6, 'sp4_h_r_13')
// (20, 6, 'sp4_h_r_24')
// (21, 6, 'sp4_h_r_37')
// (22, 6, 'sp4_h_l_37')

wire n2340;
// (16, 5, 'neigh_op_tnr_7')
// (16, 6, 'neigh_op_rgt_7')
// (16, 7, 'neigh_op_bnr_7')
// (17, 1, 'sp4_r_v_b_34')
// (17, 2, 'sp4_r_v_b_23')
// (17, 3, 'sp4_r_v_b_10')
// (17, 4, 'sp4_r_v_b_39')
// (17, 5, 'neigh_op_top_7')
// (17, 5, 'sp4_r_v_b_26')
// (17, 6, 'lutff_7/out')
// (17, 6, 'sp4_r_v_b_15')
// (17, 7, 'neigh_op_bot_7')
// (17, 7, 'sp4_r_v_b_2')
// (18, 0, 'span4_vert_34')
// (18, 1, 'sp4_v_b_34')
// (18, 2, 'sp4_v_b_23')
// (18, 3, 'local_g1_2')
// (18, 3, 'lutff_2/in_1')
// (18, 3, 'sp4_v_b_10')
// (18, 3, 'sp4_v_t_39')
// (18, 4, 'sp4_v_b_39')
// (18, 5, 'neigh_op_tnl_7')
// (18, 5, 'sp4_v_b_26')
// (18, 6, 'neigh_op_lft_7')
// (18, 6, 'sp4_v_b_15')
// (18, 7, 'neigh_op_bnl_7')
// (18, 7, 'sp4_v_b_2')

reg n2341 = 0;
// (16, 5, 'sp4_r_v_b_37')
// (16, 6, 'sp4_r_v_b_24')
// (16, 7, 'sp4_r_v_b_13')
// (16, 8, 'sp4_r_v_b_0')
// (16, 9, 'sp4_r_v_b_44')
// (16, 10, 'neigh_op_tnr_2')
// (16, 10, 'sp4_r_v_b_33')
// (16, 11, 'neigh_op_rgt_2')
// (16, 11, 'sp4_r_v_b_20')
// (16, 12, 'neigh_op_bnr_2')
// (16, 12, 'sp4_r_v_b_9')
// (17, 4, 'sp4_v_t_37')
// (17, 5, 'sp4_v_b_37')
// (17, 6, 'sp4_v_b_24')
// (17, 7, 'local_g1_5')
// (17, 7, 'lutff_6/in_0')
// (17, 7, 'lutff_7/in_3')
// (17, 7, 'sp4_v_b_13')
// (17, 8, 'sp4_v_b_0')
// (17, 8, 'sp4_v_t_44')
// (17, 9, 'sp4_r_v_b_45')
// (17, 9, 'sp4_v_b_44')
// (17, 10, 'neigh_op_top_2')
// (17, 10, 'sp4_r_v_b_32')
// (17, 10, 'sp4_v_b_33')
// (17, 11, 'local_g0_2')
// (17, 11, 'lutff_2/in_2')
// (17, 11, 'lutff_2/out')
// (17, 11, 'sp4_h_r_4')
// (17, 11, 'sp4_r_v_b_21')
// (17, 11, 'sp4_v_b_20')
// (17, 12, 'neigh_op_bot_2')
// (17, 12, 'sp4_r_v_b_8')
// (17, 12, 'sp4_v_b_9')
// (18, 8, 'local_g1_1')
// (18, 8, 'lutff_2/in_2')
// (18, 8, 'lutff_3/in_3')
// (18, 8, 'lutff_4/in_2')
// (18, 8, 'sp4_h_r_1')
// (18, 8, 'sp4_v_t_45')
// (18, 9, 'sp4_v_b_45')
// (18, 10, 'neigh_op_tnl_2')
// (18, 10, 'sp4_v_b_32')
// (18, 11, 'neigh_op_lft_2')
// (18, 11, 'sp4_h_r_17')
// (18, 11, 'sp4_v_b_21')
// (18, 12, 'neigh_op_bnl_2')
// (18, 12, 'sp4_v_b_8')
// (19, 8, 'sp4_h_r_12')
// (19, 11, 'sp4_h_r_28')
// (20, 8, 'sp4_h_r_25')
// (20, 8, 'sp4_r_v_b_47')
// (20, 9, 'local_g0_1')
// (20, 9, 'lutff_0/in_1')
// (20, 9, 'sp4_r_v_b_34')
// (20, 10, 'local_g3_7')
// (20, 10, 'lutff_0/in_0')
// (20, 10, 'lutff_1/in_3')
// (20, 10, 'sp4_r_v_b_23')
// (20, 11, 'sp4_h_r_41')
// (20, 11, 'sp4_r_v_b_10')
// (21, 7, 'sp4_v_t_47')
// (21, 8, 'sp4_h_r_36')
// (21, 8, 'sp4_v_b_47')
// (21, 9, 'sp4_v_b_34')
// (21, 10, 'sp4_v_b_23')
// (21, 11, 'sp4_h_l_41')
// (21, 11, 'sp4_v_b_10')
// (22, 8, 'sp4_h_l_36')

wire n2342;
// (16, 6, 'neigh_op_tnr_1')
// (16, 7, 'neigh_op_rgt_1')
// (16, 8, 'neigh_op_bnr_1')
// (17, 4, 'sp4_r_v_b_38')
// (17, 5, 'sp4_r_v_b_27')
// (17, 6, 'neigh_op_top_1')
// (17, 6, 'sp4_r_v_b_14')
// (17, 7, 'lutff_1/out')
// (17, 7, 'sp4_r_v_b_3')
// (17, 8, 'neigh_op_bot_1')
// (18, 3, 'local_g1_0')
// (18, 3, 'lutff_1/in_2')
// (18, 3, 'sp4_h_r_8')
// (18, 3, 'sp4_v_t_38')
// (18, 4, 'sp4_v_b_38')
// (18, 5, 'sp4_v_b_27')
// (18, 6, 'neigh_op_tnl_1')
// (18, 6, 'sp4_v_b_14')
// (18, 7, 'neigh_op_lft_1')
// (18, 7, 'sp4_v_b_3')
// (18, 8, 'neigh_op_bnl_1')
// (19, 3, 'sp4_h_r_21')
// (20, 3, 'sp4_h_r_32')
// (21, 3, 'sp4_h_r_45')
// (22, 3, 'sp4_h_l_45')

wire n2343;
// (16, 6, 'neigh_op_tnr_3')
// (16, 7, 'neigh_op_rgt_3')
// (16, 8, 'neigh_op_bnr_3')
// (17, 4, 'sp4_r_v_b_42')
// (17, 5, 'sp4_r_v_b_31')
// (17, 6, 'neigh_op_top_3')
// (17, 6, 'sp4_r_v_b_18')
// (17, 7, 'lutff_3/out')
// (17, 7, 'sp4_r_v_b_7')
// (17, 8, 'neigh_op_bot_3')
// (18, 3, 'local_g0_0')
// (18, 3, 'lutff_7/in_1')
// (18, 3, 'sp4_h_r_0')
// (18, 3, 'sp4_v_t_42')
// (18, 4, 'sp4_v_b_42')
// (18, 5, 'sp4_v_b_31')
// (18, 6, 'neigh_op_tnl_3')
// (18, 6, 'sp4_v_b_18')
// (18, 7, 'neigh_op_lft_3')
// (18, 7, 'sp4_v_b_7')
// (18, 8, 'neigh_op_bnl_3')
// (19, 3, 'sp4_h_r_13')
// (20, 3, 'sp4_h_r_24')
// (21, 3, 'sp4_h_r_37')
// (22, 3, 'sp4_h_l_37')

wire n2344;
// (16, 6, 'neigh_op_tnr_7')
// (16, 6, 'sp4_r_v_b_43')
// (16, 7, 'neigh_op_rgt_7')
// (16, 7, 'sp4_r_v_b_30')
// (16, 7, 'sp4_r_v_b_46')
// (16, 8, 'local_g3_3')
// (16, 8, 'lutff_global/cen')
// (16, 8, 'neigh_op_bnr_7')
// (16, 8, 'sp4_r_v_b_19')
// (16, 8, 'sp4_r_v_b_35')
// (16, 9, 'sp4_r_v_b_22')
// (16, 9, 'sp4_r_v_b_6')
// (16, 10, 'sp4_r_v_b_11')
// (17, 5, 'sp4_v_t_43')
// (17, 6, 'neigh_op_top_7')
// (17, 6, 'sp4_v_b_43')
// (17, 6, 'sp4_v_t_46')
// (17, 7, 'lutff_7/out')
// (17, 7, 'sp4_v_b_30')
// (17, 7, 'sp4_v_b_46')
// (17, 8, 'local_g3_3')
// (17, 8, 'lutff_global/cen')
// (17, 8, 'neigh_op_bot_7')
// (17, 8, 'sp4_v_b_19')
// (17, 8, 'sp4_v_b_35')
// (17, 9, 'sp4_v_b_22')
// (17, 9, 'sp4_v_b_6')
// (17, 10, 'sp4_v_b_11')
// (18, 6, 'neigh_op_tnl_7')
// (18, 7, 'neigh_op_lft_7')
// (18, 8, 'neigh_op_bnl_7')

wire n2345;
// (16, 6, 'sp4_r_v_b_37')
// (16, 7, 'sp4_r_v_b_24')
// (16, 8, 'sp4_r_v_b_13')
// (16, 9, 'sp4_r_v_b_0')
// (16, 11, 'sp4_h_r_2')
// (17, 5, 'sp4_v_t_37')
// (17, 6, 'sp4_r_v_b_42')
// (17, 6, 'sp4_v_b_37')
// (17, 7, 'local_g3_0')
// (17, 7, 'lutff_6/in_3')
// (17, 7, 'lutff_7/in_0')
// (17, 7, 'sp4_r_v_b_31')
// (17, 7, 'sp4_v_b_24')
// (17, 8, 'sp4_r_v_b_18')
// (17, 8, 'sp4_v_b_13')
// (17, 9, 'sp4_h_r_7')
// (17, 9, 'sp4_r_v_b_7')
// (17, 9, 'sp4_v_b_0')
// (17, 11, 'local_g0_7')
// (17, 11, 'lutff_5/in_2')
// (17, 11, 'sp4_h_r_15')
// (18, 5, 'sp4_v_t_42')
// (18, 6, 'sp4_v_b_42')
// (18, 7, 'sp4_v_b_31')
// (18, 8, 'local_g1_2')
// (18, 8, 'lutff_3/in_2')
// (18, 8, 'sp4_v_b_18')
// (18, 9, 'sp4_h_r_18')
// (18, 9, 'sp4_h_r_2')
// (18, 9, 'sp4_v_b_7')
// (18, 11, 'sp4_h_r_26')
// (19, 8, 'neigh_op_tnr_5')
// (19, 8, 'sp4_r_v_b_39')
// (19, 9, 'neigh_op_rgt_5')
// (19, 9, 'sp4_h_r_15')
// (19, 9, 'sp4_h_r_31')
// (19, 9, 'sp4_r_v_b_26')
// (19, 10, 'neigh_op_bnr_5')
// (19, 10, 'sp4_r_v_b_15')
// (19, 11, 'sp4_h_r_39')
// (19, 11, 'sp4_r_v_b_2')
// (20, 7, 'sp4_v_t_39')
// (20, 8, 'neigh_op_top_5')
// (20, 8, 'sp4_v_b_39')
// (20, 9, 'lutff_5/out')
// (20, 9, 'sp4_h_r_26')
// (20, 9, 'sp4_h_r_42')
// (20, 9, 'sp4_v_b_26')
// (20, 10, 'local_g1_5')
// (20, 10, 'lutff_1/in_1')
// (20, 10, 'neigh_op_bot_5')
// (20, 10, 'sp4_v_b_15')
// (20, 11, 'sp4_h_l_39')
// (20, 11, 'sp4_v_b_2')
// (21, 8, 'neigh_op_tnl_5')
// (21, 9, 'neigh_op_lft_5')
// (21, 9, 'sp4_h_l_42')
// (21, 9, 'sp4_h_r_39')
// (21, 10, 'neigh_op_bnl_5')
// (22, 9, 'sp4_h_l_39')

reg n2346 = 0;
// (16, 7, 'local_g2_4')
// (16, 7, 'lutff_4/in_2')
// (16, 7, 'sp4_r_v_b_36')
// (16, 8, 'neigh_op_tnr_6')
// (16, 8, 'sp4_r_v_b_25')
// (16, 9, 'local_g2_6')
// (16, 9, 'lutff_5/in_3')
// (16, 9, 'neigh_op_rgt_6')
// (16, 9, 'sp4_r_v_b_12')
// (16, 10, 'neigh_op_bnr_6')
// (16, 10, 'sp4_r_v_b_1')
// (17, 6, 'sp4_v_t_36')
// (17, 7, 'sp4_v_b_36')
// (17, 8, 'neigh_op_top_6')
// (17, 8, 'sp4_v_b_25')
// (17, 9, 'lutff_6/out')
// (17, 9, 'sp4_v_b_12')
// (17, 10, 'neigh_op_bot_6')
// (17, 10, 'sp4_v_b_1')
// (18, 8, 'neigh_op_tnl_6')
// (18, 9, 'neigh_op_lft_6')
// (18, 10, 'neigh_op_bnl_6')

reg n2347 = 0;
// (16, 7, 'neigh_op_tnr_0')
// (16, 8, 'neigh_op_rgt_0')
// (16, 9, 'neigh_op_bnr_0')
// (17, 7, 'neigh_op_top_0')
// (17, 8, 'lutff_0/out')
// (17, 9, 'local_g1_0')
// (17, 9, 'lutff_4/in_1')
// (17, 9, 'neigh_op_bot_0')
// (18, 7, 'neigh_op_tnl_0')
// (18, 8, 'neigh_op_lft_0')
// (18, 9, 'neigh_op_bnl_0')

reg n2348 = 0;
// (16, 7, 'neigh_op_tnr_1')
// (16, 8, 'neigh_op_rgt_1')
// (16, 9, 'neigh_op_bnr_1')
// (17, 7, 'neigh_op_top_1')
// (17, 8, 'lutff_1/out')
// (17, 9, 'neigh_op_bot_1')
// (18, 7, 'neigh_op_tnl_1')
// (18, 8, 'neigh_op_lft_1')
// (18, 9, 'local_g2_1')
// (18, 9, 'lutff_4/in_1')
// (18, 9, 'neigh_op_bnl_1')

wire n2349;
// (16, 7, 'neigh_op_tnr_2')
// (16, 8, 'neigh_op_rgt_2')
// (16, 9, 'neigh_op_bnr_2')
// (17, 6, 'sp4_r_v_b_45')
// (17, 7, 'neigh_op_top_2')
// (17, 7, 'sp4_r_v_b_32')
// (17, 8, 'lutff_2/out')
// (17, 8, 'sp4_r_v_b_21')
// (17, 9, 'local_g2_0')
// (17, 9, 'lutff_2/in_2')
// (17, 9, 'neigh_op_bot_2')
// (17, 9, 'sp4_r_v_b_8')
// (18, 5, 'sp4_v_t_45')
// (18, 6, 'sp4_v_b_45')
// (18, 7, 'neigh_op_tnl_2')
// (18, 7, 'sp4_v_b_32')
// (18, 8, 'neigh_op_lft_2')
// (18, 8, 'sp4_v_b_21')
// (18, 9, 'neigh_op_bnl_2')
// (18, 9, 'sp4_v_b_8')

reg n2350 = 0;
// (16, 7, 'neigh_op_tnr_3')
// (16, 8, 'neigh_op_rgt_3')
// (16, 9, 'neigh_op_bnr_3')
// (17, 7, 'neigh_op_top_3')
// (17, 8, 'local_g1_3')
// (17, 8, 'lutff_3/out')
// (17, 8, 'lutff_4/in_2')
// (17, 9, 'neigh_op_bot_3')
// (18, 7, 'neigh_op_tnl_3')
// (18, 8, 'neigh_op_lft_3')
// (18, 9, 'neigh_op_bnl_3')

wire n2351;
// (16, 7, 'neigh_op_tnr_4')
// (16, 8, 'neigh_op_rgt_4')
// (16, 9, 'local_g1_4')
// (16, 9, 'lutff_7/in_2')
// (16, 9, 'neigh_op_bnr_4')
// (17, 7, 'neigh_op_top_4')
// (17, 8, 'lutff_4/out')
// (17, 9, 'neigh_op_bot_4')
// (18, 7, 'neigh_op_tnl_4')
// (18, 8, 'neigh_op_lft_4')
// (18, 9, 'neigh_op_bnl_4')

reg n2352 = 0;
// (16, 7, 'neigh_op_tnr_5')
// (16, 8, 'neigh_op_rgt_5')
// (16, 9, 'neigh_op_bnr_5')
// (17, 7, 'neigh_op_top_5')
// (17, 8, 'lutff_5/out')
// (17, 9, 'local_g0_5')
// (17, 9, 'lutff_3/in_0')
// (17, 9, 'neigh_op_bot_5')
// (18, 7, 'neigh_op_tnl_5')
// (18, 8, 'neigh_op_lft_5')
// (18, 9, 'neigh_op_bnl_5')

reg n2353 = 0;
// (16, 7, 'neigh_op_tnr_6')
// (16, 8, 'neigh_op_rgt_6')
// (16, 9, 'neigh_op_bnr_6')
// (17, 7, 'neigh_op_top_6')
// (17, 8, 'lutff_6/out')
// (17, 8, 'sp4_r_v_b_45')
// (17, 9, 'neigh_op_bot_6')
// (17, 9, 'sp4_r_v_b_32')
// (17, 10, 'sp4_r_v_b_21')
// (17, 11, 'sp4_r_v_b_8')
// (18, 7, 'neigh_op_tnl_6')
// (18, 7, 'sp4_v_t_45')
// (18, 8, 'neigh_op_lft_6')
// (18, 8, 'sp4_v_b_45')
// (18, 9, 'neigh_op_bnl_6')
// (18, 9, 'sp4_v_b_32')
// (18, 10, 'sp4_v_b_21')
// (18, 11, 'local_g0_0')
// (18, 11, 'lutff_2/in_0')
// (18, 11, 'sp4_v_b_8')

reg n2354 = 0;
// (16, 7, 'neigh_op_tnr_7')
// (16, 8, 'neigh_op_rgt_7')
// (16, 9, 'neigh_op_bnr_7')
// (17, 7, 'neigh_op_top_7')
// (17, 8, 'lutff_7/out')
// (17, 9, 'local_g0_7')
// (17, 9, 'lutff_5/in_2')
// (17, 9, 'neigh_op_bot_7')
// (18, 7, 'neigh_op_tnl_7')
// (18, 8, 'neigh_op_lft_7')
// (18, 9, 'neigh_op_bnl_7')

wire n2355;
// (16, 7, 'sp4_r_v_b_39')
// (16, 8, 'sp4_r_v_b_26')
// (16, 9, 'local_g2_1')
// (16, 9, 'local_g3_1')
// (16, 9, 'lutff_0/in_0')
// (16, 9, 'lutff_1/in_3')
// (16, 9, 'lutff_3/in_3')
// (16, 9, 'lutff_6/in_1')
// (16, 9, 'lutff_7/in_0')
// (16, 9, 'neigh_op_tnr_1')
// (16, 9, 'sp4_r_v_b_15')
// (16, 10, 'local_g2_1')
// (16, 10, 'lutff_1/in_2')
// (16, 10, 'lutff_2/in_1')
// (16, 10, 'lutff_4/in_3')
// (16, 10, 'neigh_op_rgt_1')
// (16, 10, 'sp4_r_v_b_2')
// (16, 11, 'local_g0_1')
// (16, 11, 'lutff_5/in_2')
// (16, 11, 'lutff_6/in_1')
// (16, 11, 'neigh_op_bnr_1')
// (17, 6, 'sp4_v_t_39')
// (17, 7, 'sp4_v_b_39')
// (17, 8, 'local_g2_2')
// (17, 8, 'lutff_2/in_0')
// (17, 8, 'sp4_v_b_26')
// (17, 9, 'local_g1_1')
// (17, 9, 'lutff_3/in_3')
// (17, 9, 'lutff_4/in_2')
// (17, 9, 'lutff_5/in_1')
// (17, 9, 'lutff_7/in_1')
// (17, 9, 'neigh_op_top_1')
// (17, 9, 'sp4_v_b_15')
// (17, 10, 'local_g1_1')
// (17, 10, 'lutff_1/out')
// (17, 10, 'lutff_4/in_2')
// (17, 10, 'lutff_5/in_1')
// (17, 10, 'sp4_v_b_2')
// (17, 11, 'local_g1_1')
// (17, 11, 'lutff_3/in_3')
// (17, 11, 'lutff_6/in_2')
// (17, 11, 'neigh_op_bot_1')
// (18, 9, 'local_g3_1')
// (18, 9, 'lutff_1/in_3')
// (18, 9, 'lutff_2/in_2')
// (18, 9, 'lutff_3/in_3')
// (18, 9, 'lutff_4/in_2')
// (18, 9, 'lutff_6/in_2')
// (18, 9, 'lutff_7/in_1')
// (18, 9, 'neigh_op_tnl_1')
// (18, 10, 'local_g1_1')
// (18, 10, 'lutff_1/in_1')
// (18, 10, 'lutff_3/in_1')
// (18, 10, 'lutff_5/in_3')
// (18, 10, 'neigh_op_lft_1')
// (18, 11, 'local_g2_1')
// (18, 11, 'lutff_2/in_1')
// (18, 11, 'lutff_3/in_2')
// (18, 11, 'neigh_op_bnl_1')

reg n2356 = 0;
// (16, 8, 'local_g3_0')
// (16, 8, 'lutff_3/in_0')
// (16, 8, 'neigh_op_tnr_0')
// (16, 9, 'local_g3_0')
// (16, 9, 'lutff_3/in_0')
// (16, 9, 'neigh_op_rgt_0')
// (16, 10, 'neigh_op_bnr_0')
// (17, 8, 'neigh_op_top_0')
// (17, 9, 'lutff_0/out')
// (17, 10, 'neigh_op_bot_0')
// (18, 8, 'neigh_op_tnl_0')
// (18, 9, 'neigh_op_lft_0')
// (18, 10, 'neigh_op_bnl_0')

reg n2357 = 0;
// (16, 8, 'local_g3_1')
// (16, 8, 'lutff_0/in_0')
// (16, 8, 'neigh_op_tnr_1')
// (16, 9, 'neigh_op_rgt_1')
// (16, 10, 'neigh_op_bnr_1')
// (17, 8, 'neigh_op_top_1')
// (17, 9, 'local_g2_1')
// (17, 9, 'lutff_1/out')
// (17, 9, 'lutff_7/in_2')
// (17, 10, 'neigh_op_bot_1')
// (18, 8, 'neigh_op_tnl_1')
// (18, 9, 'neigh_op_lft_1')
// (18, 10, 'neigh_op_bnl_1')

wire n2358;
// (16, 8, 'neigh_op_tnr_2')
// (16, 9, 'neigh_op_rgt_2')
// (16, 9, 'sp4_r_v_b_36')
// (16, 10, 'neigh_op_bnr_2')
// (16, 10, 'sp4_r_v_b_25')
// (16, 11, 'sp4_r_v_b_12')
// (16, 12, 'local_g1_1')
// (16, 12, 'lutff_3/in_1')
// (16, 12, 'sp4_r_v_b_1')
// (17, 8, 'neigh_op_top_2')
// (17, 8, 'sp4_v_t_36')
// (17, 9, 'lutff_2/out')
// (17, 9, 'sp4_v_b_36')
// (17, 10, 'neigh_op_bot_2')
// (17, 10, 'sp4_v_b_25')
// (17, 11, 'sp4_v_b_12')
// (17, 12, 'sp4_v_b_1')
// (18, 8, 'neigh_op_tnl_2')
// (18, 9, 'neigh_op_lft_2')
// (18, 10, 'neigh_op_bnl_2')

wire n2359;
// (16, 8, 'neigh_op_tnr_3')
// (16, 9, 'local_g2_3')
// (16, 9, 'lutff_3/in_2')
// (16, 9, 'neigh_op_rgt_3')
// (16, 10, 'neigh_op_bnr_3')
// (17, 8, 'neigh_op_top_3')
// (17, 9, 'lutff_3/out')
// (17, 10, 'neigh_op_bot_3')
// (18, 8, 'neigh_op_tnl_3')
// (18, 9, 'neigh_op_lft_3')
// (18, 10, 'neigh_op_bnl_3')

wire n2360;
// (16, 8, 'neigh_op_tnr_4')
// (16, 9, 'neigh_op_rgt_4')
// (16, 10, 'neigh_op_bnr_4')
// (17, 8, 'local_g0_4')
// (17, 8, 'lutff_2/in_2')
// (17, 8, 'neigh_op_top_4')
// (17, 9, 'lutff_4/out')
// (17, 10, 'neigh_op_bot_4')
// (18, 8, 'neigh_op_tnl_4')
// (18, 9, 'neigh_op_lft_4')
// (18, 10, 'neigh_op_bnl_4')

wire n2361;
// (16, 8, 'neigh_op_tnr_5')
// (16, 9, 'neigh_op_rgt_5')
// (16, 10, 'local_g0_5')
// (16, 10, 'lutff_6/in_3')
// (16, 10, 'neigh_op_bnr_5')
// (17, 8, 'neigh_op_top_5')
// (17, 9, 'lutff_5/out')
// (17, 10, 'neigh_op_bot_5')
// (18, 8, 'neigh_op_tnl_5')
// (18, 9, 'neigh_op_lft_5')
// (18, 10, 'neigh_op_bnl_5')

wire n2362;
// (16, 8, 'neigh_op_tnr_7')
// (16, 9, 'neigh_op_rgt_7')
// (16, 10, 'neigh_op_bnr_7')
// (17, 8, 'neigh_op_top_7')
// (17, 9, 'lutff_7/out')
// (17, 10, 'neigh_op_bot_7')
// (18, 8, 'neigh_op_tnl_7')
// (18, 9, 'neigh_op_lft_7')
// (18, 10, 'local_g3_7')
// (18, 10, 'lutff_2/in_0')
// (18, 10, 'neigh_op_bnl_7')

wire n2363;
// (16, 8, 'sp4_h_r_9')
// (17, 5, 'sp4_h_r_9')
// (17, 8, 'sp4_h_r_20')
// (18, 5, 'sp4_h_r_20')
// (18, 8, 'sp4_h_r_33')
// (19, 4, 'neigh_op_tnr_6')
// (19, 5, 'local_g2_1')
// (19, 5, 'local_g2_6')
// (19, 5, 'neigh_op_rgt_6')
// (19, 5, 'ram/MASK_10')
// (19, 5, 'ram/MASK_11')
// (19, 5, 'ram/MASK_12')
// (19, 5, 'ram/MASK_13')
// (19, 5, 'ram/MASK_14')
// (19, 5, 'ram/MASK_15')
// (19, 5, 'ram/MASK_8')
// (19, 5, 'ram/MASK_9')
// (19, 5, 'sp4_h_r_33')
// (19, 5, 'sp4_r_v_b_44')
// (19, 6, 'local_g0_6')
// (19, 6, 'local_g1_6')
// (19, 6, 'neigh_op_bnr_6')
// (19, 6, 'ram/MASK_0')
// (19, 6, 'ram/MASK_1')
// (19, 6, 'ram/MASK_2')
// (19, 6, 'ram/MASK_3')
// (19, 6, 'ram/MASK_4')
// (19, 6, 'ram/MASK_5')
// (19, 6, 'ram/MASK_6')
// (19, 6, 'ram/MASK_7')
// (19, 6, 'sp4_r_v_b_33')
// (19, 7, 'sp4_r_v_b_20')
// (19, 8, 'local_g2_1')
// (19, 8, 'local_g2_4')
// (19, 8, 'ram/MASK_0')
// (19, 8, 'ram/MASK_1')
// (19, 8, 'ram/MASK_2')
// (19, 8, 'ram/MASK_3')
// (19, 8, 'sp4_h_r_44')
// (19, 8, 'sp4_r_v_b_9')
// (20, 4, 'neigh_op_top_6')
// (20, 4, 'sp4_v_t_44')
// (20, 5, 'lutff_6/out')
// (20, 5, 'sp4_h_r_44')
// (20, 5, 'sp4_v_b_44')
// (20, 6, 'neigh_op_bot_6')
// (20, 6, 'sp4_v_b_33')
// (20, 7, 'sp4_v_b_20')
// (20, 8, 'sp4_h_l_44')
// (20, 8, 'sp4_v_b_9')
// (21, 4, 'neigh_op_tnl_6')
// (21, 5, 'neigh_op_lft_6')
// (21, 5, 'sp4_h_l_44')
// (21, 6, 'neigh_op_bnl_6')

wire n2364;
// (16, 8, 'sp4_r_v_b_36')
// (16, 9, 'local_g3_6')
// (16, 9, 'lutff_0/in_3')
// (16, 9, 'lutff_1/in_2')
// (16, 9, 'lutff_2/in_1')
// (16, 9, 'lutff_5/in_2')
// (16, 9, 'lutff_6/in_3')
// (16, 9, 'neigh_op_tnr_6')
// (16, 9, 'sp4_r_v_b_25')
// (16, 10, 'local_g2_6')
// (16, 10, 'lutff_2/in_2')
// (16, 10, 'lutff_4/in_0')
// (16, 10, 'lutff_7/in_1')
// (16, 10, 'neigh_op_rgt_6')
// (16, 10, 'sp4_r_v_b_12')
// (16, 11, 'local_g1_6')
// (16, 11, 'lutff_5/in_0')
// (16, 11, 'lutff_6/in_3')
// (16, 11, 'neigh_op_bnr_6')
// (16, 11, 'sp4_r_v_b_1')
// (17, 7, 'sp4_v_t_36')
// (17, 8, 'local_g2_4')
// (17, 8, 'lutff_4/in_0')
// (17, 8, 'sp4_v_b_36')
// (17, 9, 'local_g0_6')
// (17, 9, 'local_g1_6')
// (17, 9, 'lutff_3/in_2')
// (17, 9, 'lutff_4/in_3')
// (17, 9, 'lutff_5/in_3')
// (17, 9, 'neigh_op_top_6')
// (17, 9, 'sp4_v_b_25')
// (17, 10, 'local_g2_6')
// (17, 10, 'lutff_5/in_3')
// (17, 10, 'lutff_6/out')
// (17, 10, 'sp4_v_b_12')
// (17, 11, 'local_g0_6')
// (17, 11, 'lutff_3/in_1')
// (17, 11, 'lutff_6/in_0')
// (17, 11, 'neigh_op_bot_6')
// (17, 11, 'sp4_v_b_1')
// (18, 9, 'local_g2_6')
// (18, 9, 'local_g3_6')
// (18, 9, 'lutff_1/in_1')
// (18, 9, 'lutff_2/in_3')
// (18, 9, 'lutff_3/in_0')
// (18, 9, 'lutff_4/in_0')
// (18, 9, 'lutff_7/in_2')
// (18, 9, 'neigh_op_tnl_6')
// (18, 10, 'local_g1_6')
// (18, 10, 'lutff_1/in_2')
// (18, 10, 'lutff_3/in_0')
// (18, 10, 'lutff_5/in_0')
// (18, 10, 'neigh_op_lft_6')
// (18, 11, 'local_g3_6')
// (18, 11, 'lutff_2/in_3')
// (18, 11, 'neigh_op_bnl_6')

reg n2365 = 0;
// (16, 8, 'sp4_r_v_b_38')
// (16, 9, 'sp4_r_v_b_27')
// (16, 10, 'sp4_r_v_b_14')
// (16, 11, 'sp4_r_v_b_3')
// (17, 7, 'sp4_v_t_38')
// (17, 8, 'sp4_v_b_38')
// (17, 9, 'sp4_v_b_27')
// (17, 10, 'local_g1_6')
// (17, 10, 'lutff_4/in_1')
// (17, 10, 'sp4_v_b_14')
// (17, 11, 'sp4_h_r_3')
// (17, 11, 'sp4_v_b_3')
// (18, 11, 'sp4_h_r_14')
// (19, 11, 'sp4_h_r_27')
// (20, 10, 'neigh_op_tnr_0')
// (20, 11, 'neigh_op_rgt_0')
// (20, 11, 'sp4_h_r_38')
// (20, 12, 'neigh_op_bnr_0')
// (21, 10, 'neigh_op_top_0')
// (21, 11, 'lutff_0/out')
// (21, 11, 'sp4_h_l_38')
// (21, 11, 'sp4_h_r_0')
// (21, 12, 'neigh_op_bot_0')
// (22, 10, 'neigh_op_tnl_0')
// (22, 11, 'neigh_op_lft_0')
// (22, 11, 'sp4_h_r_13')
// (22, 12, 'neigh_op_bnl_0')
// (23, 11, 'sp4_h_r_24')
// (24, 11, 'sp4_h_r_37')
// (25, 11, 'sp4_h_l_37')

wire n2366;
// (16, 9, 'local_g2_2')
// (16, 9, 'lutff_7/in_3')
// (16, 9, 'neigh_op_tnr_2')
// (16, 10, 'local_g2_2')
// (16, 10, 'lutff_1/in_1')
// (16, 10, 'lutff_3/in_1')
// (16, 10, 'lutff_6/in_0')
// (16, 10, 'neigh_op_rgt_2')
// (16, 11, 'local_g0_2')
// (16, 11, 'lutff_3/in_3')
// (16, 11, 'lutff_4/in_2')
// (16, 11, 'neigh_op_bnr_2')
// (17, 9, 'local_g1_2')
// (17, 9, 'lutff_2/in_3')
// (17, 9, 'neigh_op_top_2')
// (17, 10, 'lutff_2/out')
// (17, 11, 'local_g1_2')
// (17, 11, 'lutff_7/in_2')
// (17, 11, 'neigh_op_bot_2')
// (18, 9, 'local_g3_2')
// (18, 9, 'lutff_0/in_3')
// (18, 9, 'neigh_op_tnl_2')
// (18, 10, 'local_g1_2')
// (18, 10, 'lutff_2/in_1')
// (18, 10, 'neigh_op_lft_2')
// (18, 11, 'neigh_op_bnl_2')

reg n2367 = 0;
// (16, 9, 'neigh_op_tnr_3')
// (16, 10, 'neigh_op_rgt_3')
// (16, 11, 'neigh_op_bnr_3')
// (17, 9, 'neigh_op_top_3')
// (17, 10, 'lutff_3/out')
// (17, 11, 'local_g0_3')
// (17, 11, 'lutff_6/in_3')
// (17, 11, 'neigh_op_bot_3')
// (18, 9, 'neigh_op_tnl_3')
// (18, 10, 'neigh_op_lft_3')
// (18, 11, 'neigh_op_bnl_3')

wire n2368;
// (16, 9, 'neigh_op_tnr_4')
// (16, 10, 'local_g2_4')
// (16, 10, 'lutff_6/in_2')
// (16, 10, 'neigh_op_rgt_4')
// (16, 11, 'neigh_op_bnr_4')
// (17, 9, 'neigh_op_top_4')
// (17, 10, 'lutff_4/out')
// (17, 11, 'neigh_op_bot_4')
// (18, 9, 'neigh_op_tnl_4')
// (18, 10, 'neigh_op_lft_4')
// (18, 11, 'neigh_op_bnl_4')

wire n2369;
// (16, 9, 'neigh_op_tnr_5')
// (16, 10, 'neigh_op_rgt_5')
// (16, 11, 'neigh_op_bnr_5')
// (17, 9, 'neigh_op_top_5')
// (17, 10, 'lutff_5/out')
// (17, 11, 'neigh_op_bot_5')
// (18, 9, 'neigh_op_tnl_5')
// (18, 10, 'neigh_op_lft_5')
// (18, 11, 'local_g2_5')
// (18, 11, 'lutff_3/in_0')
// (18, 11, 'neigh_op_bnl_5')

reg n2370 = 0;
// (16, 9, 'neigh_op_tnr_7')
// (16, 10, 'neigh_op_rgt_7')
// (16, 11, 'neigh_op_bnr_7')
// (17, 9, 'neigh_op_top_7')
// (17, 10, 'lutff_7/out')
// (17, 11, 'neigh_op_bot_7')
// (18, 9, 'local_g3_7')
// (18, 9, 'lutff_3/in_1')
// (18, 9, 'neigh_op_tnl_7')
// (18, 10, 'neigh_op_lft_7')
// (18, 11, 'neigh_op_bnl_7')

reg n2371 = 0;
// (16, 9, 'sp4_h_r_3')
// (17, 9, 'sp4_h_r_14')
// (18, 9, 'local_g2_3')
// (18, 9, 'lutff_1/in_0')
// (18, 9, 'sp4_h_r_27')
// (19, 9, 'neigh_op_tnr_3')
// (19, 9, 'sp4_h_r_38')
// (19, 10, 'neigh_op_rgt_3')
// (19, 10, 'sp4_r_v_b_38')
// (19, 11, 'neigh_op_bnr_3')
// (19, 11, 'sp4_r_v_b_27')
// (19, 12, 'sp4_r_v_b_14')
// (19, 13, 'sp4_r_v_b_3')
// (20, 9, 'neigh_op_top_3')
// (20, 9, 'sp4_h_l_38')
// (20, 9, 'sp4_v_t_38')
// (20, 10, 'lutff_3/out')
// (20, 10, 'sp4_v_b_38')
// (20, 11, 'neigh_op_bot_3')
// (20, 11, 'sp4_v_b_27')
// (20, 12, 'sp4_v_b_14')
// (20, 13, 'sp4_v_b_3')
// (21, 9, 'neigh_op_tnl_3')
// (21, 10, 'neigh_op_lft_3')
// (21, 11, 'neigh_op_bnl_3')

reg n2372 = 0;
// (16, 9, 'sp4_h_r_9')
// (17, 9, 'local_g1_4')
// (17, 9, 'lutff_5/in_0')
// (17, 9, 'sp4_h_r_20')
// (18, 9, 'sp4_h_r_33')
// (19, 6, 'sp4_r_v_b_41')
// (19, 7, 'sp4_r_v_b_28')
// (19, 8, 'neigh_op_tnr_2')
// (19, 8, 'sp4_r_v_b_17')
// (19, 9, 'neigh_op_rgt_2')
// (19, 9, 'sp4_h_r_44')
// (19, 9, 'sp4_r_v_b_4')
// (19, 10, 'neigh_op_bnr_2')
// (20, 5, 'sp4_v_t_41')
// (20, 6, 'sp4_v_b_41')
// (20, 7, 'sp4_v_b_28')
// (20, 8, 'neigh_op_top_2')
// (20, 8, 'sp4_v_b_17')
// (20, 9, 'lutff_2/out')
// (20, 9, 'sp4_h_l_44')
// (20, 9, 'sp4_v_b_4')
// (20, 10, 'neigh_op_bot_2')
// (21, 8, 'neigh_op_tnl_2')
// (21, 9, 'neigh_op_lft_2')
// (21, 10, 'neigh_op_bnl_2')

reg n2373 = 0;
// (16, 9, 'sp4_r_v_b_41')
// (16, 10, 'sp4_r_v_b_28')
// (16, 11, 'sp4_r_v_b_17')
// (16, 12, 'sp4_r_v_b_4')
// (17, 8, 'sp4_v_t_41')
// (17, 9, 'sp4_v_b_41')
// (17, 10, 'local_g3_4')
// (17, 10, 'lutff_5/in_0')
// (17, 10, 'sp4_v_b_28')
// (17, 11, 'sp4_v_b_17')
// (17, 12, 'sp4_h_r_11')
// (17, 12, 'sp4_v_b_4')
// (18, 12, 'sp4_h_r_22')
// (19, 11, 'neigh_op_tnr_7')
// (19, 12, 'neigh_op_rgt_7')
// (19, 12, 'sp4_h_r_35')
// (19, 13, 'neigh_op_bnr_7')
// (20, 11, 'neigh_op_top_7')
// (20, 12, 'lutff_7/out')
// (20, 12, 'sp4_h_r_46')
// (20, 13, 'neigh_op_bot_7')
// (21, 11, 'neigh_op_tnl_7')
// (21, 12, 'neigh_op_lft_7')
// (21, 12, 'sp4_h_l_46')
// (21, 13, 'neigh_op_bnl_7')

reg n2374 = 0;
// (16, 10, 'local_g0_0')
// (16, 10, 'lutff_4/in_2')
// (16, 10, 'sp4_h_r_0')
// (17, 9, 'neigh_op_tnr_4')
// (17, 10, 'neigh_op_rgt_4')
// (17, 10, 'sp4_h_r_13')
// (17, 11, 'neigh_op_bnr_4')
// (18, 9, 'neigh_op_top_4')
// (18, 10, 'lutff_4/out')
// (18, 10, 'sp4_h_r_24')
// (18, 11, 'neigh_op_bot_4')
// (19, 9, 'neigh_op_tnl_4')
// (19, 10, 'neigh_op_lft_4')
// (19, 10, 'sp4_h_r_37')
// (19, 11, 'neigh_op_bnl_4')
// (20, 10, 'sp4_h_l_37')

reg n2375 = 0;
// (16, 10, 'neigh_op_tnr_1')
// (16, 11, 'neigh_op_rgt_1')
// (16, 12, 'neigh_op_bnr_1')
// (17, 4, 'sp4_r_v_b_43')
// (17, 5, 'sp4_r_v_b_30')
// (17, 6, 'sp4_r_v_b_19')
// (17, 7, 'local_g1_6')
// (17, 7, 'lutff_6/in_1')
// (17, 7, 'lutff_7/in_2')
// (17, 7, 'sp4_r_v_b_6')
// (17, 8, 'sp4_r_v_b_38')
// (17, 9, 'sp4_r_v_b_27')
// (17, 10, 'neigh_op_top_1')
// (17, 10, 'sp4_r_v_b_14')
// (17, 10, 'sp4_r_v_b_46')
// (17, 11, 'local_g3_1')
// (17, 11, 'lutff_1/in_1')
// (17, 11, 'lutff_1/out')
// (17, 11, 'sp4_h_r_2')
// (17, 11, 'sp4_r_v_b_3')
// (17, 11, 'sp4_r_v_b_35')
// (17, 12, 'neigh_op_bot_1')
// (17, 12, 'sp4_r_v_b_22')
// (17, 13, 'sp4_r_v_b_11')
// (18, 3, 'sp4_v_t_43')
// (18, 4, 'sp4_v_b_43')
// (18, 5, 'sp4_v_b_30')
// (18, 6, 'sp4_v_b_19')
// (18, 7, 'sp4_v_b_6')
// (18, 7, 'sp4_v_t_38')
// (18, 8, 'local_g3_6')
// (18, 8, 'lutff_2/in_3')
// (18, 8, 'lutff_3/in_0')
// (18, 8, 'lutff_4/in_3')
// (18, 8, 'sp4_v_b_38')
// (18, 9, 'sp4_h_r_11')
// (18, 9, 'sp4_v_b_27')
// (18, 9, 'sp4_v_t_46')
// (18, 10, 'neigh_op_tnl_1')
// (18, 10, 'sp4_v_b_14')
// (18, 10, 'sp4_v_b_46')
// (18, 11, 'neigh_op_lft_1')
// (18, 11, 'sp4_h_r_15')
// (18, 11, 'sp4_v_b_3')
// (18, 11, 'sp4_v_b_35')
// (18, 12, 'neigh_op_bnl_1')
// (18, 12, 'sp4_v_b_22')
// (18, 13, 'sp4_v_b_11')
// (19, 9, 'sp4_h_r_22')
// (19, 11, 'sp4_h_r_26')
// (20, 8, 'sp4_r_v_b_39')
// (20, 9, 'local_g2_3')
// (20, 9, 'lutff_0/in_3')
// (20, 9, 'sp4_h_r_35')
// (20, 9, 'sp4_r_v_b_26')
// (20, 10, 'local_g2_7')
// (20, 10, 'lutff_0/in_3')
// (20, 10, 'lutff_1/in_0')
// (20, 10, 'sp4_r_v_b_15')
// (20, 11, 'sp4_h_r_39')
// (20, 11, 'sp4_r_v_b_2')
// (21, 7, 'sp4_v_t_39')
// (21, 8, 'sp4_v_b_39')
// (21, 9, 'sp4_h_r_46')
// (21, 9, 'sp4_v_b_26')
// (21, 10, 'sp4_v_b_15')
// (21, 11, 'sp4_h_l_39')
// (21, 11, 'sp4_v_b_2')
// (22, 9, 'sp4_h_l_46')

wire n2376;
// (16, 10, 'neigh_op_tnr_3')
// (16, 11, 'local_g2_3')
// (16, 11, 'lutff_4/in_3')
// (16, 11, 'neigh_op_rgt_3')
// (16, 12, 'neigh_op_bnr_3')
// (17, 10, 'neigh_op_top_3')
// (17, 11, 'lutff_3/out')
// (17, 12, 'neigh_op_bot_3')
// (18, 10, 'neigh_op_tnl_3')
// (18, 11, 'neigh_op_lft_3')
// (18, 12, 'neigh_op_bnl_3')

reg n2377 = 0;
// (16, 10, 'neigh_op_tnr_5')
// (16, 11, 'neigh_op_rgt_5')
// (16, 11, 'sp4_r_v_b_42')
// (16, 12, 'neigh_op_bnr_5')
// (16, 12, 'sp4_r_v_b_31')
// (16, 13, 'sp4_r_v_b_18')
// (16, 14, 'sp4_r_v_b_7')
// (17, 8, 'sp4_r_v_b_46')
// (17, 9, 'sp4_r_v_b_35')
// (17, 10, 'neigh_op_top_5')
// (17, 10, 'sp4_h_r_7')
// (17, 10, 'sp4_r_v_b_22')
// (17, 10, 'sp4_r_v_b_38')
// (17, 10, 'sp4_v_t_42')
// (17, 11, 'local_g3_5')
// (17, 11, 'lutff_0/in_2')
// (17, 11, 'lutff_1/in_3')
// (17, 11, 'lutff_5/out')
// (17, 11, 'sp4_r_v_b_11')
// (17, 11, 'sp4_r_v_b_27')
// (17, 11, 'sp4_v_b_42')
// (17, 12, 'neigh_op_bot_5')
// (17, 12, 'sp4_r_v_b_14')
// (17, 12, 'sp4_v_b_31')
// (17, 13, 'sp4_r_v_b_3')
// (17, 13, 'sp4_v_b_18')
// (17, 14, 'sp4_v_b_7')
// (18, 7, 'sp4_v_t_46')
// (18, 8, 'local_g2_6')
// (18, 8, 'lutff_2/in_0')
// (18, 8, 'lutff_4/in_0')
// (18, 8, 'sp4_v_b_46')
// (18, 9, 'sp4_h_r_3')
// (18, 9, 'sp4_v_b_35')
// (18, 9, 'sp4_v_t_38')
// (18, 10, 'neigh_op_tnl_5')
// (18, 10, 'sp4_h_r_18')
// (18, 10, 'sp4_v_b_22')
// (18, 10, 'sp4_v_b_38')
// (18, 11, 'neigh_op_lft_5')
// (18, 11, 'sp4_v_b_11')
// (18, 11, 'sp4_v_b_27')
// (18, 12, 'neigh_op_bnl_5')
// (18, 12, 'sp4_v_b_14')
// (18, 13, 'sp4_v_b_3')
// (19, 9, 'sp4_h_r_14')
// (19, 10, 'sp4_h_r_31')
// (20, 9, 'local_g3_3')
// (20, 9, 'lutff_0/in_0')
// (20, 9, 'lutff_5/in_3')
// (20, 9, 'sp4_h_r_27')
// (20, 10, 'local_g3_2')
// (20, 10, 'lutff_0/in_1')
// (20, 10, 'sp4_h_r_42')
// (21, 9, 'sp4_h_r_38')
// (21, 10, 'sp4_h_l_42')
// (22, 9, 'sp4_h_l_38')

wire n2378;
// (16, 10, 'neigh_op_tnr_7')
// (16, 11, 'neigh_op_rgt_7')
// (16, 12, 'neigh_op_bnr_7')
// (17, 10, 'neigh_op_top_7')
// (17, 11, 'lutff_7/out')
// (17, 12, 'local_g0_7')
// (17, 12, 'lutff_5/in_2')
// (17, 12, 'neigh_op_bot_7')
// (18, 10, 'neigh_op_tnl_7')
// (18, 11, 'neigh_op_lft_7')
// (18, 12, 'neigh_op_bnl_7')

wire n2379;
// (16, 10, 'sp4_r_v_b_40')
// (16, 11, 'sp4_r_v_b_29')
// (16, 12, 'sp4_r_v_b_16')
// (16, 13, 'sp4_r_v_b_5')
// (17, 8, 'neigh_op_tnr_0')
// (17, 9, 'neigh_op_rgt_0')
// (17, 9, 'sp4_h_r_5')
// (17, 9, 'sp4_v_t_40')
// (17, 10, 'neigh_op_bnr_0')
// (17, 10, 'sp4_v_b_40')
// (17, 11, 'sp4_v_b_29')
// (17, 12, 'local_g0_0')
// (17, 12, 'lutff_4/in_2')
// (17, 12, 'sp4_v_b_16')
// (17, 13, 'sp4_v_b_5')
// (18, 8, 'neigh_op_top_0')
// (18, 9, 'lutff_0/out')
// (18, 9, 'sp4_h_r_16')
// (18, 10, 'neigh_op_bot_0')
// (19, 8, 'neigh_op_tnl_0')
// (19, 9, 'neigh_op_lft_0')
// (19, 9, 'sp4_h_r_29')
// (19, 10, 'neigh_op_bnl_0')
// (20, 9, 'sp4_h_r_40')
// (21, 9, 'sp4_h_l_40')

reg n2380 = 0;
// (16, 11, 'neigh_op_tnr_0')
// (16, 12, 'neigh_op_rgt_0')
// (16, 13, 'neigh_op_bnr_0')
// (17, 11, 'neigh_op_top_0')
// (17, 12, 'lutff_0/out')
// (17, 12, 'sp4_h_r_0')
// (17, 13, 'neigh_op_bot_0')
// (18, 11, 'neigh_op_tnl_0')
// (18, 12, 'neigh_op_lft_0')
// (18, 12, 'sp4_h_r_13')
// (18, 13, 'neigh_op_bnl_0')
// (19, 12, 'sp4_h_r_24')
// (20, 12, 'local_g3_5')
// (20, 12, 'lutff_0/in_2')
// (20, 12, 'sp4_h_r_37')
// (21, 12, 'sp4_h_l_37')

reg n2381 = 0;
// (16, 11, 'neigh_op_tnr_3')
// (16, 12, 'neigh_op_rgt_3')
// (16, 13, 'neigh_op_bnr_3')
// (17, 11, 'neigh_op_top_3')
// (17, 12, 'lutff_3/out')
// (17, 13, 'neigh_op_bot_3')
// (18, 11, 'neigh_op_tnl_3')
// (18, 12, 'local_g1_3')
// (18, 12, 'lutff_7/in_1')
// (18, 12, 'neigh_op_lft_3')
// (18, 13, 'neigh_op_bnl_3')

wire n2382;
// (16, 11, 'neigh_op_tnr_4')
// (16, 12, 'local_g2_4')
// (16, 12, 'lutff_5/in_1')
// (16, 12, 'neigh_op_rgt_4')
// (16, 13, 'neigh_op_bnr_4')
// (17, 11, 'neigh_op_top_4')
// (17, 12, 'lutff_4/out')
// (17, 13, 'neigh_op_bot_4')
// (18, 11, 'neigh_op_tnl_4')
// (18, 12, 'neigh_op_lft_4')
// (18, 13, 'neigh_op_bnl_4')

wire n2383;
// (16, 11, 'neigh_op_tnr_5')
// (16, 12, 'neigh_op_rgt_5')
// (16, 13, 'local_g1_5')
// (16, 13, 'lutff_0/in_0')
// (16, 13, 'neigh_op_bnr_5')
// (17, 11, 'neigh_op_top_5')
// (17, 12, 'lutff_5/out')
// (17, 13, 'neigh_op_bot_5')
// (18, 11, 'neigh_op_tnl_5')
// (18, 12, 'neigh_op_lft_5')
// (18, 13, 'neigh_op_bnl_5')

wire n2384;
// (16, 11, 'sp4_r_v_b_38')
// (16, 12, 'local_g0_3')
// (16, 12, 'lutff_4/in_3')
// (16, 12, 'sp4_r_v_b_27')
// (16, 13, 'sp4_r_v_b_14')
// (16, 14, 'sp4_r_v_b_3')
// (17, 9, 'neigh_op_tnr_2')
// (17, 10, 'neigh_op_rgt_2')
// (17, 10, 'sp4_h_r_9')
// (17, 10, 'sp4_v_t_38')
// (17, 11, 'neigh_op_bnr_2')
// (17, 11, 'sp4_v_b_38')
// (17, 12, 'sp4_v_b_27')
// (17, 13, 'sp4_v_b_14')
// (17, 14, 'sp4_v_b_3')
// (18, 9, 'neigh_op_top_2')
// (18, 10, 'lutff_2/out')
// (18, 10, 'sp4_h_r_20')
// (18, 11, 'neigh_op_bot_2')
// (19, 9, 'neigh_op_tnl_2')
// (19, 10, 'neigh_op_lft_2')
// (19, 10, 'sp4_h_r_33')
// (19, 11, 'neigh_op_bnl_2')
// (20, 10, 'sp4_h_r_44')
// (21, 10, 'sp4_h_l_44')

reg n2385 = 0;
// (16, 11, 'sp4_r_v_b_44')
// (16, 12, 'neigh_op_tnr_2')
// (16, 12, 'sp4_r_v_b_33')
// (16, 13, 'neigh_op_rgt_2')
// (16, 13, 'sp4_h_r_9')
// (16, 13, 'sp4_r_v_b_20')
// (16, 14, 'neigh_op_bnr_2')
// (16, 14, 'sp4_r_v_b_9')
// (17, 10, 'sp4_v_t_44')
// (17, 11, 'sp4_r_v_b_45')
// (17, 11, 'sp4_v_b_44')
// (17, 12, 'neigh_op_top_2')
// (17, 12, 'sp4_r_v_b_32')
// (17, 12, 'sp4_v_b_33')
// (17, 13, 'local_g0_2')
// (17, 13, 'lutff_2/in_2')
// (17, 13, 'lutff_2/out')
// (17, 13, 'sp4_h_r_20')
// (17, 13, 'sp4_r_v_b_21')
// (17, 13, 'sp4_v_b_20')
// (17, 14, 'neigh_op_bot_2')
// (17, 14, 'sp4_h_r_3')
// (17, 14, 'sp4_r_v_b_8')
// (17, 14, 'sp4_v_b_9')
// (18, 10, 'sp4_h_r_1')
// (18, 10, 'sp4_v_t_45')
// (18, 11, 'sp4_v_b_45')
// (18, 12, 'neigh_op_tnl_2')
// (18, 12, 'sp4_v_b_32')
// (18, 13, 'neigh_op_lft_2')
// (18, 13, 'sp4_h_r_33')
// (18, 13, 'sp4_v_b_21')
// (18, 14, 'neigh_op_bnl_2')
// (18, 14, 'sp4_h_r_14')
// (18, 14, 'sp4_v_b_8')
// (19, 10, 'local_g1_4')
// (19, 10, 'ram/WADDR_2')
// (19, 10, 'sp4_h_r_12')
// (19, 10, 'sp4_r_v_b_44')
// (19, 11, 'sp4_r_v_b_33')
// (19, 12, 'local_g3_4')
// (19, 12, 'ram/WADDR_2')
// (19, 12, 'sp4_r_v_b_20')
// (19, 13, 'sp4_h_r_44')
// (19, 13, 'sp4_r_v_b_9')
// (19, 14, 'local_g2_3')
// (19, 14, 'ram/WADDR_2')
// (19, 14, 'sp4_h_r_27')
// (20, 9, 'sp4_v_t_44')
// (20, 10, 'sp4_h_r_25')
// (20, 10, 'sp4_v_b_44')
// (20, 11, 'sp4_v_b_33')
// (20, 12, 'sp4_v_b_20')
// (20, 13, 'sp4_h_l_44')
// (20, 13, 'sp4_v_b_9')
// (20, 14, 'sp4_h_r_38')
// (21, 10, 'sp4_h_r_36')
// (21, 14, 'sp4_h_l_38')
// (22, 10, 'sp4_h_l_36')

reg n2386 = 0;
// (16, 12, 'neigh_op_tnr_1')
// (16, 13, 'neigh_op_rgt_1')
// (16, 13, 'sp4_h_r_7')
// (16, 14, 'neigh_op_bnr_1')
// (17, 11, 'sp4_r_v_b_43')
// (17, 12, 'neigh_op_top_1')
// (17, 12, 'sp4_r_v_b_30')
// (17, 13, 'local_g1_1')
// (17, 13, 'lutff_1/in_1')
// (17, 13, 'lutff_1/out')
// (17, 13, 'sp4_h_r_18')
// (17, 13, 'sp4_r_v_b_19')
// (17, 14, 'neigh_op_bot_1')
// (17, 14, 'sp4_r_v_b_6')
// (18, 10, 'sp4_v_t_43')
// (18, 11, 'sp4_v_b_43')
// (18, 12, 'neigh_op_tnl_1')
// (18, 12, 'sp4_v_b_30')
// (18, 13, 'neigh_op_lft_1')
// (18, 13, 'sp4_h_r_31')
// (18, 13, 'sp4_v_b_19')
// (18, 14, 'neigh_op_bnl_1')
// (18, 14, 'sp4_h_r_0')
// (18, 14, 'sp4_v_b_6')
// (19, 10, 'local_g2_4')
// (19, 10, 'ram/WADDR_1')
// (19, 10, 'sp4_r_v_b_36')
// (19, 11, 'sp4_r_v_b_25')
// (19, 12, 'local_g2_4')
// (19, 12, 'ram/WADDR_1')
// (19, 12, 'sp4_r_v_b_12')
// (19, 13, 'sp4_h_r_42')
// (19, 13, 'sp4_r_v_b_1')
// (19, 14, 'local_g1_5')
// (19, 14, 'ram/WADDR_1')
// (19, 14, 'sp4_h_r_13')
// (20, 9, 'sp4_v_t_36')
// (20, 10, 'sp4_v_b_36')
// (20, 11, 'sp4_v_b_25')
// (20, 12, 'sp4_v_b_12')
// (20, 13, 'sp4_h_l_42')
// (20, 13, 'sp4_v_b_1')
// (20, 14, 'sp4_h_r_24')
// (21, 14, 'sp4_h_r_37')
// (22, 14, 'sp4_h_l_37')

reg n2387 = 0;
// (16, 12, 'neigh_op_tnr_3')
// (16, 13, 'neigh_op_rgt_3')
// (16, 13, 'sp4_r_v_b_38')
// (16, 14, 'neigh_op_bnr_3')
// (16, 14, 'sp4_r_v_b_27')
// (16, 15, 'sp4_r_v_b_14')
// (16, 16, 'sp4_r_v_b_3')
// (17, 11, 'sp4_r_v_b_47')
// (17, 12, 'neigh_op_top_3')
// (17, 12, 'sp4_h_r_8')
// (17, 12, 'sp4_r_v_b_34')
// (17, 12, 'sp4_v_t_38')
// (17, 13, 'local_g1_3')
// (17, 13, 'lutff_3/in_1')
// (17, 13, 'lutff_3/out')
// (17, 13, 'sp4_r_v_b_23')
// (17, 13, 'sp4_v_b_38')
// (17, 14, 'neigh_op_bot_3')
// (17, 14, 'sp4_r_v_b_10')
// (17, 14, 'sp4_v_b_27')
// (17, 15, 'sp4_v_b_14')
// (17, 16, 'sp4_v_b_3')
// (18, 10, 'sp4_h_r_10')
// (18, 10, 'sp4_v_t_47')
// (18, 11, 'sp4_v_b_47')
// (18, 12, 'neigh_op_tnl_3')
// (18, 12, 'sp4_h_r_21')
// (18, 12, 'sp4_v_b_34')
// (18, 13, 'neigh_op_lft_3')
// (18, 13, 'sp4_v_b_23')
// (18, 14, 'neigh_op_bnl_3')
// (18, 14, 'sp4_h_r_10')
// (18, 14, 'sp4_v_b_10')
// (19, 10, 'local_g1_7')
// (19, 10, 'ram/WADDR_3')
// (19, 10, 'sp4_h_r_23')
// (19, 12, 'local_g2_0')
// (19, 12, 'ram/WADDR_3')
// (19, 12, 'sp4_h_r_32')
// (19, 14, 'local_g1_7')
// (19, 14, 'ram/WADDR_3')
// (19, 14, 'sp4_h_r_23')
// (20, 10, 'sp4_h_r_34')
// (20, 12, 'sp4_h_r_45')
// (20, 14, 'sp4_h_r_34')
// (21, 10, 'sp4_h_r_47')
// (21, 12, 'sp4_h_l_45')
// (21, 14, 'sp4_h_r_47')
// (22, 10, 'sp4_h_l_47')
// (22, 14, 'sp4_h_l_47')

reg n2388 = 0;
// (16, 12, 'neigh_op_tnr_6')
// (16, 13, 'neigh_op_rgt_6')
// (16, 13, 'sp4_h_r_1')
// (16, 14, 'neigh_op_bnr_6')
// (17, 11, 'sp4_r_v_b_37')
// (17, 12, 'neigh_op_top_6')
// (17, 12, 'sp4_r_v_b_24')
// (17, 13, 'local_g2_6')
// (17, 13, 'lutff_6/in_0')
// (17, 13, 'lutff_6/out')
// (17, 13, 'sp4_h_r_12')
// (17, 13, 'sp4_r_v_b_13')
// (17, 14, 'neigh_op_bot_6')
// (17, 14, 'sp4_r_v_b_0')
// (18, 10, 'sp4_v_t_37')
// (18, 11, 'sp4_v_b_37')
// (18, 12, 'neigh_op_tnl_6')
// (18, 12, 'sp4_v_b_24')
// (18, 13, 'neigh_op_lft_6')
// (18, 13, 'sp4_h_r_25')
// (18, 13, 'sp4_v_b_13')
// (18, 14, 'neigh_op_bnl_6')
// (18, 14, 'sp4_h_r_6')
// (18, 14, 'sp4_v_b_0')
// (19, 10, 'local_g3_2')
// (19, 10, 'ram/WADDR_6')
// (19, 10, 'sp4_r_v_b_42')
// (19, 11, 'sp4_r_v_b_31')
// (19, 12, 'local_g3_2')
// (19, 12, 'ram/WADDR_6')
// (19, 12, 'sp4_r_v_b_18')
// (19, 13, 'sp4_h_r_36')
// (19, 13, 'sp4_r_v_b_7')
// (19, 14, 'local_g0_3')
// (19, 14, 'ram/WADDR_6')
// (19, 14, 'sp4_h_r_19')
// (20, 9, 'sp4_v_t_42')
// (20, 10, 'sp4_v_b_42')
// (20, 11, 'sp4_v_b_31')
// (20, 12, 'sp4_v_b_18')
// (20, 13, 'sp4_h_l_36')
// (20, 13, 'sp4_v_b_7')
// (20, 14, 'sp4_h_r_30')
// (21, 14, 'sp4_h_r_43')
// (22, 14, 'sp4_h_l_43')

wire n2389;
// (16, 12, 'sp4_h_r_1')
// (17, 12, 'local_g1_4')
// (17, 12, 'lutff_3/in_0')
// (17, 12, 'sp4_h_r_12')
// (18, 11, 'neigh_op_tnr_2')
// (18, 12, 'neigh_op_rgt_2')
// (18, 12, 'sp4_h_r_25')
// (18, 13, 'neigh_op_bnr_2')
// (19, 11, 'neigh_op_top_2')
// (19, 12, 'ram/RDATA_5')
// (19, 12, 'sp4_h_r_36')
// (19, 13, 'neigh_op_bot_2')
// (20, 11, 'neigh_op_tnl_2')
// (20, 12, 'neigh_op_lft_2')
// (20, 12, 'sp4_h_l_36')
// (20, 13, 'neigh_op_bnl_2')

wire n2390;
// (16, 12, 'sp4_h_r_6')
// (17, 11, 'neigh_op_tnr_7')
// (17, 12, 'neigh_op_rgt_7')
// (17, 12, 'sp4_h_r_19')
// (17, 13, 'neigh_op_bnr_7')
// (18, 11, 'neigh_op_top_7')
// (18, 12, 'lutff_7/out')
// (18, 12, 'sp4_h_r_30')
// (18, 13, 'neigh_op_bot_7')
// (19, 11, 'neigh_op_tnl_7')
// (19, 12, 'neigh_op_lft_7')
// (19, 12, 'sp4_h_r_43')
// (19, 13, 'neigh_op_bnl_7')
// (20, 12, 'sp4_h_l_43')
// (20, 12, 'sp4_h_r_6')
// (21, 12, 'local_g0_3')
// (21, 12, 'lutff_1/in_2')
// (21, 12, 'sp4_h_r_19')
// (22, 12, 'sp4_h_r_30')
// (23, 12, 'sp4_h_r_43')
// (24, 12, 'sp4_h_l_43')

reg n2391 = 0;
// (16, 13, 'neigh_op_tnr_2')
// (16, 14, 'neigh_op_rgt_2')
// (16, 14, 'sp4_h_r_9')
// (16, 15, 'neigh_op_bnr_2')
// (17, 12, 'sp4_r_v_b_45')
// (17, 13, 'neigh_op_top_2')
// (17, 13, 'sp4_r_v_b_32')
// (17, 14, 'local_g3_2')
// (17, 14, 'lutff_2/in_1')
// (17, 14, 'lutff_2/out')
// (17, 14, 'sp4_h_r_20')
// (17, 14, 'sp4_r_v_b_21')
// (17, 14, 'sp4_r_v_b_37')
// (17, 15, 'neigh_op_bot_2')
// (17, 15, 'sp4_r_v_b_24')
// (17, 15, 'sp4_r_v_b_8')
// (17, 16, 'sp4_r_v_b_13')
// (17, 17, 'sp4_r_v_b_0')
// (18, 11, 'sp4_h_r_8')
// (18, 11, 'sp4_v_t_45')
// (18, 12, 'sp4_v_b_45')
// (18, 13, 'neigh_op_tnl_2')
// (18, 13, 'sp4_h_r_5')
// (18, 13, 'sp4_v_b_32')
// (18, 13, 'sp4_v_t_37')
// (18, 14, 'neigh_op_lft_2')
// (18, 14, 'sp4_h_r_33')
// (18, 14, 'sp4_v_b_21')
// (18, 14, 'sp4_v_b_37')
// (18, 15, 'neigh_op_bnl_2')
// (18, 15, 'sp4_v_b_24')
// (18, 15, 'sp4_v_b_8')
// (18, 16, 'sp4_v_b_13')
// (18, 17, 'sp4_v_b_0')
// (19, 7, 'sp4_r_v_b_46')
// (19, 8, 'sp4_r_v_b_35')
// (19, 9, 'local_g3_6')
// (19, 9, 'ram/RADDR_2')
// (19, 9, 'sp4_r_v_b_22')
// (19, 10, 'sp4_r_v_b_11')
// (19, 11, 'local_g0_5')
// (19, 11, 'ram/RADDR_2')
// (19, 11, 'sp4_h_r_21')
// (19, 11, 'sp4_r_v_b_38')
// (19, 12, 'sp4_r_v_b_27')
// (19, 13, 'local_g1_0')
// (19, 13, 'ram/RADDR_2')
// (19, 13, 'sp4_h_r_16')
// (19, 13, 'sp4_r_v_b_14')
// (19, 14, 'sp4_h_r_44')
// (19, 14, 'sp4_r_v_b_3')
// (20, 6, 'sp4_v_t_46')
// (20, 7, 'sp4_v_b_46')
// (20, 8, 'sp4_v_b_35')
// (20, 9, 'sp4_v_b_22')
// (20, 10, 'sp4_v_b_11')
// (20, 10, 'sp4_v_t_38')
// (20, 11, 'sp4_h_r_32')
// (20, 11, 'sp4_v_b_38')
// (20, 12, 'sp4_v_b_27')
// (20, 13, 'sp4_h_r_29')
// (20, 13, 'sp4_v_b_14')
// (20, 14, 'sp4_h_l_44')
// (20, 14, 'sp4_v_b_3')
// (21, 11, 'sp4_h_r_45')
// (21, 13, 'sp4_h_r_40')
// (22, 11, 'sp4_h_l_45')
// (22, 13, 'sp4_h_l_40')

reg n2392 = 0;
// (16, 13, 'neigh_op_tnr_3')
// (16, 14, 'neigh_op_rgt_3')
// (16, 15, 'neigh_op_bnr_3')
// (17, 10, 'sp4_r_v_b_47')
// (17, 11, 'sp4_r_v_b_34')
// (17, 12, 'sp4_r_v_b_23')
// (17, 12, 'sp4_r_v_b_47')
// (17, 13, 'neigh_op_top_3')
// (17, 13, 'sp4_r_v_b_10')
// (17, 13, 'sp4_r_v_b_34')
// (17, 14, 'local_g0_3')
// (17, 14, 'lutff_3/in_2')
// (17, 14, 'lutff_3/out')
// (17, 14, 'sp4_r_v_b_23')
// (17, 14, 'sp4_r_v_b_39')
// (17, 15, 'neigh_op_bot_3')
// (17, 15, 'sp4_r_v_b_10')
// (17, 15, 'sp4_r_v_b_26')
// (17, 16, 'sp4_r_v_b_15')
// (17, 17, 'sp4_r_v_b_2')
// (18, 9, 'sp4_h_r_10')
// (18, 9, 'sp4_v_t_47')
// (18, 10, 'sp4_v_b_47')
// (18, 11, 'sp4_h_r_3')
// (18, 11, 'sp4_v_b_34')
// (18, 11, 'sp4_v_t_47')
// (18, 12, 'sp4_v_b_23')
// (18, 12, 'sp4_v_b_47')
// (18, 13, 'neigh_op_tnl_3')
// (18, 13, 'sp4_h_r_2')
// (18, 13, 'sp4_v_b_10')
// (18, 13, 'sp4_v_b_34')
// (18, 13, 'sp4_v_t_39')
// (18, 14, 'neigh_op_lft_3')
// (18, 14, 'sp4_v_b_23')
// (18, 14, 'sp4_v_b_39')
// (18, 15, 'neigh_op_bnl_3')
// (18, 15, 'sp4_v_b_10')
// (18, 15, 'sp4_v_b_26')
// (18, 16, 'sp4_v_b_15')
// (18, 17, 'sp4_v_b_2')
// (19, 9, 'local_g1_7')
// (19, 9, 'ram/RADDR_3')
// (19, 9, 'sp4_h_r_23')
// (19, 11, 'local_g0_6')
// (19, 11, 'ram/RADDR_3')
// (19, 11, 'sp4_h_r_14')
// (19, 13, 'local_g1_7')
// (19, 13, 'ram/RADDR_3')
// (19, 13, 'sp4_h_r_15')
// (20, 9, 'sp4_h_r_34')
// (20, 11, 'sp4_h_r_27')
// (20, 13, 'sp4_h_r_26')
// (21, 9, 'sp4_h_r_47')
// (21, 11, 'sp4_h_r_38')
// (21, 13, 'sp4_h_r_39')
// (22, 9, 'sp4_h_l_47')
// (22, 11, 'sp4_h_l_38')
// (22, 13, 'sp4_h_l_39')

reg n2393 = 0;
// (16, 13, 'neigh_op_tnr_6')
// (16, 14, 'neigh_op_rgt_6')
// (16, 14, 'sp4_h_r_1')
// (16, 15, 'neigh_op_bnr_6')
// (17, 13, 'neigh_op_top_6')
// (17, 14, 'local_g2_6')
// (17, 14, 'lutff_6/in_0')
// (17, 14, 'lutff_6/out')
// (17, 14, 'sp4_h_r_12')
// (17, 15, 'neigh_op_bot_6')
// (18, 13, 'neigh_op_tnl_6')
// (18, 14, 'neigh_op_lft_6')
// (18, 14, 'sp4_h_r_25')
// (18, 15, 'neigh_op_bnl_6')
// (19, 7, 'sp4_r_v_b_42')
// (19, 8, 'sp4_r_v_b_31')
// (19, 9, 'local_g3_2')
// (19, 9, 'ram/RADDR_6')
// (19, 9, 'sp4_r_v_b_18')
// (19, 10, 'sp4_r_v_b_7')
// (19, 11, 'local_g3_2')
// (19, 11, 'ram/RADDR_6')
// (19, 11, 'sp4_r_v_b_42')
// (19, 12, 'sp4_r_v_b_31')
// (19, 13, 'local_g3_2')
// (19, 13, 'ram/RADDR_6')
// (19, 13, 'sp4_r_v_b_18')
// (19, 14, 'sp4_h_r_36')
// (19, 14, 'sp4_r_v_b_7')
// (20, 6, 'sp4_v_t_42')
// (20, 7, 'sp4_v_b_42')
// (20, 8, 'sp4_v_b_31')
// (20, 9, 'sp4_v_b_18')
// (20, 10, 'sp4_v_b_7')
// (20, 10, 'sp4_v_t_42')
// (20, 11, 'sp4_v_b_42')
// (20, 12, 'sp4_v_b_31')
// (20, 13, 'sp4_v_b_18')
// (20, 14, 'sp4_h_l_36')
// (20, 14, 'sp4_v_b_7')

reg n2394 = 0;
// (16, 13, 'neigh_op_tnr_7')
// (16, 14, 'neigh_op_rgt_7')
// (16, 14, 'sp4_h_r_3')
// (16, 15, 'neigh_op_bnr_7')
// (17, 13, 'neigh_op_top_7')
// (17, 14, 'local_g0_7')
// (17, 14, 'local_g3_7')
// (17, 14, 'lutff_0/in_1')
// (17, 14, 'lutff_1/in_3')
// (17, 14, 'lutff_7/in_2')
// (17, 14, 'lutff_7/out')
// (17, 14, 'sp4_h_r_14')
// (17, 15, 'neigh_op_bot_7')
// (18, 13, 'neigh_op_tnl_7')
// (18, 14, 'neigh_op_lft_7')
// (18, 14, 'sp4_h_r_27')
// (18, 15, 'neigh_op_bnl_7')
// (19, 7, 'sp4_r_v_b_40')
// (19, 8, 'sp4_r_v_b_29')
// (19, 9, 'local_g3_0')
// (19, 9, 'ram/RADDR_0')
// (19, 9, 'sp4_r_v_b_16')
// (19, 10, 'sp4_r_v_b_5')
// (19, 11, 'local_g3_4')
// (19, 11, 'ram/RADDR_0')
// (19, 11, 'sp4_r_v_b_44')
// (19, 12, 'sp4_r_v_b_33')
// (19, 13, 'local_g3_4')
// (19, 13, 'ram/RADDR_0')
// (19, 13, 'sp4_r_v_b_20')
// (19, 14, 'sp4_h_r_38')
// (19, 14, 'sp4_r_v_b_9')
// (20, 6, 'sp4_v_t_40')
// (20, 7, 'sp4_v_b_40')
// (20, 8, 'sp4_v_b_29')
// (20, 9, 'sp4_v_b_16')
// (20, 10, 'sp4_v_b_5')
// (20, 10, 'sp4_v_t_44')
// (20, 11, 'sp4_v_b_44')
// (20, 12, 'sp4_v_b_33')
// (20, 13, 'sp4_v_b_20')
// (20, 14, 'sp4_h_l_38')
// (20, 14, 'sp4_v_b_9')

wire n2395;
// (16, 13, 'sp4_r_v_b_44')
// (16, 14, 'sp4_r_v_b_33')
// (16, 15, 'sp4_r_v_b_20')
// (16, 16, 'sp4_r_v_b_9')
// (17, 12, 'sp4_h_r_3')
// (17, 12, 'sp4_v_t_44')
// (17, 13, 'sp4_v_b_44')
// (17, 14, 'sp4_v_b_33')
// (17, 15, 'local_g0_4')
// (17, 15, 'lutff_3/in_1')
// (17, 15, 'sp4_v_b_20')
// (17, 16, 'local_g1_1')
// (17, 16, 'lutff_4/in_0')
// (17, 16, 'sp4_v_b_9')
// (18, 12, 'sp4_h_r_14')
// (19, 11, 'sp4_h_r_4')
// (19, 12, 'sp4_h_r_27')
// (20, 11, 'sp4_h_r_17')
// (20, 12, 'sp4_h_r_38')
// (21, 11, 'neigh_op_tnr_7')
// (21, 11, 'sp4_h_r_28')
// (21, 12, 'neigh_op_rgt_7')
// (21, 12, 'sp4_h_l_38')
// (21, 12, 'sp4_h_r_3')
// (21, 13, 'neigh_op_bnr_7')
// (22, 10, 'sp4_r_v_b_39')
// (22, 11, 'neigh_op_top_7')
// (22, 11, 'sp4_h_r_41')
// (22, 11, 'sp4_r_v_b_26')
// (22, 12, 'local_g3_7')
// (22, 12, 'lutff_2/in_0')
// (22, 12, 'lutff_7/out')
// (22, 12, 'sp4_h_r_14')
// (22, 12, 'sp4_r_v_b_15')
// (22, 12, 'sp4_r_v_b_47')
// (22, 13, 'local_g0_7')
// (22, 13, 'lutff_4/in_1')
// (22, 13, 'neigh_op_bot_7')
// (22, 13, 'sp4_r_v_b_2')
// (22, 13, 'sp4_r_v_b_34')
// (22, 14, 'sp4_r_v_b_23')
// (22, 15, 'sp4_r_v_b_10')
// (23, 9, 'sp4_v_t_39')
// (23, 10, 'sp4_v_b_39')
// (23, 11, 'local_g0_4')
// (23, 11, 'lutff_global/s_r')
// (23, 11, 'neigh_op_tnl_7')
// (23, 11, 'sp4_h_l_41')
// (23, 11, 'sp4_h_r_4')
// (23, 11, 'sp4_v_b_26')
// (23, 11, 'sp4_v_t_47')
// (23, 12, 'neigh_op_lft_7')
// (23, 12, 'sp4_h_r_27')
// (23, 12, 'sp4_v_b_15')
// (23, 12, 'sp4_v_b_47')
// (23, 13, 'neigh_op_bnl_7')
// (23, 13, 'sp4_h_r_8')
// (23, 13, 'sp4_v_b_2')
// (23, 13, 'sp4_v_b_34')
// (23, 14, 'sp4_v_b_23')
// (23, 15, 'sp4_v_b_10')
// (24, 11, 'sp4_h_r_17')
// (24, 12, 'sp4_h_r_38')
// (24, 13, 'local_g1_5')
// (24, 13, 'lutff_global/s_r')
// (24, 13, 'sp4_h_r_21')
// (25, 11, 'sp4_h_r_28')
// (25, 12, 'sp4_h_l_38')
// (25, 13, 'sp4_h_r_32')

wire n2396;
// (16, 14, 'neigh_op_tnr_2')
// (16, 15, 'neigh_op_rgt_2')
// (16, 16, 'neigh_op_bnr_2')
// (17, 14, 'local_g0_2')
// (17, 14, 'lutff_global/cen')
// (17, 14, 'neigh_op_top_2')
// (17, 15, 'lutff_2/out')
// (17, 16, 'neigh_op_bot_2')
// (18, 14, 'neigh_op_tnl_2')
// (18, 15, 'neigh_op_lft_2')
// (18, 16, 'neigh_op_bnl_2')

reg n2397 = 0;
// (16, 14, 'neigh_op_tnr_4')
// (16, 15, 'neigh_op_rgt_4')
// (16, 16, 'neigh_op_bnr_4')
// (17, 12, 'sp4_r_v_b_44')
// (17, 13, 'sp4_r_v_b_33')
// (17, 14, 'neigh_op_top_4')
// (17, 14, 'sp4_r_v_b_20')
// (17, 15, 'local_g2_4')
// (17, 15, 'lutff_3/in_3')
// (17, 15, 'lutff_4/out')
// (17, 15, 'sp4_r_v_b_9')
// (17, 16, 'local_g1_4')
// (17, 16, 'lutff_4/in_3')
// (17, 16, 'neigh_op_bot_4')
// (17, 16, 'sp4_r_v_b_44')
// (17, 17, 'sp4_r_v_b_33')
// (17, 18, 'sp4_r_v_b_20')
// (17, 19, 'sp4_r_v_b_9')
// (18, 11, 'sp4_v_t_44')
// (18, 12, 'sp4_v_b_44')
// (18, 13, 'sp4_v_b_33')
// (18, 14, 'neigh_op_tnl_4')
// (18, 14, 'sp4_v_b_20')
// (18, 15, 'neigh_op_lft_4')
// (18, 15, 'sp4_v_b_9')
// (18, 15, 'sp4_v_t_44')
// (18, 16, 'neigh_op_bnl_4')
// (18, 16, 'sp4_v_b_44')
// (18, 17, 'sp4_v_b_33')
// (18, 18, 'sp4_v_b_20')
// (18, 19, 'local_g0_1')
// (18, 19, 'lutff_3/in_0')
// (18, 19, 'sp4_v_b_9')

reg n2398 = 0;
// (16, 15, 'neigh_op_tnr_2')
// (16, 16, 'neigh_op_rgt_2')
// (16, 16, 'sp4_h_r_9')
// (16, 17, 'neigh_op_bnr_2')
// (17, 15, 'neigh_op_top_2')
// (17, 16, 'lutff_2/out')
// (17, 16, 'sp4_h_r_20')
// (17, 17, 'neigh_op_bot_2')
// (18, 15, 'neigh_op_tnl_2')
// (18, 16, 'neigh_op_lft_2')
// (18, 16, 'sp4_h_r_33')
// (18, 17, 'neigh_op_bnl_2')
// (19, 9, 'sp4_r_v_b_40')
// (19, 10, 'local_g0_5')
// (19, 10, 'ram/WDATA_1')
// (19, 10, 'sp4_r_v_b_29')
// (19, 11, 'sp4_r_v_b_16')
// (19, 12, 'sp4_r_v_b_5')
// (19, 13, 'sp4_r_v_b_44')
// (19, 14, 'sp4_r_v_b_33')
// (19, 15, 'sp4_r_v_b_20')
// (19, 16, 'sp4_h_r_44')
// (19, 16, 'sp4_r_v_b_9')
// (20, 8, 'sp4_v_t_40')
// (20, 9, 'sp4_v_b_40')
// (20, 10, 'sp4_v_b_29')
// (20, 11, 'sp4_v_b_16')
// (20, 12, 'sp4_v_b_5')
// (20, 12, 'sp4_v_t_44')
// (20, 13, 'sp4_v_b_44')
// (20, 14, 'sp4_v_b_33')
// (20, 15, 'sp4_v_b_20')
// (20, 16, 'sp4_h_l_44')
// (20, 16, 'sp4_v_b_9')

reg n2399 = 0;
// (16, 15, 'neigh_op_tnr_3')
// (16, 16, 'neigh_op_rgt_3')
// (16, 16, 'sp4_h_r_11')
// (16, 17, 'neigh_op_bnr_3')
// (17, 15, 'neigh_op_top_3')
// (17, 16, 'lutff_3/out')
// (17, 16, 'sp4_h_r_22')
// (17, 17, 'neigh_op_bot_3')
// (18, 15, 'neigh_op_tnl_3')
// (18, 16, 'neigh_op_lft_3')
// (18, 16, 'sp4_h_r_35')
// (18, 17, 'neigh_op_bnl_3')
// (19, 13, 'sp4_r_v_b_40')
// (19, 14, 'local_g0_5')
// (19, 14, 'ram/WDATA_5')
// (19, 14, 'sp4_r_v_b_29')
// (19, 15, 'sp4_r_v_b_16')
// (19, 16, 'sp4_h_r_46')
// (19, 16, 'sp4_r_v_b_5')
// (20, 12, 'sp4_v_t_40')
// (20, 13, 'sp4_v_b_40')
// (20, 14, 'sp4_v_b_29')
// (20, 15, 'sp4_v_b_16')
// (20, 16, 'sp4_h_l_46')
// (20, 16, 'sp4_v_b_5')

wire n2400;
// (16, 15, 'neigh_op_tnr_4')
// (16, 16, 'local_g3_4')
// (16, 16, 'lutff_0/in_3')
// (16, 16, 'lutff_2/in_3')
// (16, 16, 'neigh_op_rgt_4')
// (16, 17, 'neigh_op_bnr_4')
// (17, 15, 'neigh_op_top_4')
// (17, 16, 'lutff_4/out')
// (17, 17, 'neigh_op_bot_4')
// (18, 15, 'neigh_op_tnl_4')
// (18, 16, 'neigh_op_lft_4')
// (18, 17, 'neigh_op_bnl_4')

reg n2401 = 0;
// (16, 15, 'neigh_op_tnr_6')
// (16, 15, 'sp4_r_v_b_41')
// (16, 16, 'neigh_op_rgt_6')
// (16, 16, 'sp4_r_v_b_28')
// (16, 17, 'neigh_op_bnr_6')
// (16, 17, 'sp4_r_v_b_17')
// (16, 18, 'sp4_r_v_b_4')
// (17, 14, 'sp4_h_r_4')
// (17, 14, 'sp4_v_t_41')
// (17, 15, 'neigh_op_top_6')
// (17, 15, 'sp4_v_b_41')
// (17, 16, 'lutff_6/out')
// (17, 16, 'sp4_v_b_28')
// (17, 17, 'neigh_op_bot_6')
// (17, 17, 'sp4_v_b_17')
// (17, 18, 'sp4_v_b_4')
// (18, 14, 'sp4_h_r_17')
// (18, 15, 'neigh_op_tnl_6')
// (18, 16, 'neigh_op_lft_6')
// (18, 17, 'neigh_op_bnl_6')
// (19, 14, 'local_g3_4')
// (19, 14, 'ram/WDATA_7')
// (19, 14, 'sp4_h_r_28')
// (20, 14, 'sp4_h_r_41')
// (21, 14, 'sp4_h_l_41')

wire n2402;
// (16, 15, 'sp4_h_r_2')
// (17, 14, 'neigh_op_tnr_5')
// (17, 15, 'neigh_op_rgt_5')
// (17, 15, 'sp4_h_r_15')
// (17, 16, 'neigh_op_bnr_5')
// (18, 14, 'neigh_op_top_5')
// (18, 15, 'local_g2_2')
// (18, 15, 'lutff_5/out')
// (18, 15, 'lutff_global/cen')
// (18, 15, 'sp4_h_r_26')
// (18, 16, 'neigh_op_bot_5')
// (19, 14, 'neigh_op_tnl_5')
// (19, 15, 'neigh_op_lft_5')
// (19, 15, 'sp4_h_r_39')
// (19, 16, 'neigh_op_bnl_5')
// (20, 15, 'sp4_h_l_39')

reg n2403 = 0;
// (16, 15, 'sp4_r_v_b_44')
// (16, 16, 'neigh_op_tnr_2')
// (16, 16, 'sp4_r_v_b_33')
// (16, 17, 'neigh_op_rgt_2')
// (16, 17, 'sp4_r_v_b_20')
// (16, 18, 'neigh_op_bnr_2')
// (16, 18, 'sp4_r_v_b_9')
// (16, 19, 'sp4_r_v_b_37')
// (16, 20, 'sp4_r_v_b_24')
// (16, 21, 'sp4_r_v_b_13')
// (16, 22, 'sp4_r_v_b_0')
// (17, 14, 'sp4_v_t_44')
// (17, 15, 'sp4_r_v_b_45')
// (17, 15, 'sp4_v_b_44')
// (17, 16, 'neigh_op_top_2')
// (17, 16, 'sp4_r_v_b_32')
// (17, 16, 'sp4_v_b_33')
// (17, 17, 'lutff_2/out')
// (17, 17, 'sp4_h_r_4')
// (17, 17, 'sp4_r_v_b_21')
// (17, 17, 'sp4_r_v_b_37')
// (17, 17, 'sp4_v_b_20')
// (17, 18, 'local_g0_2')
// (17, 18, 'lutff_6/in_2')
// (17, 18, 'neigh_op_bot_2')
// (17, 18, 'sp4_r_v_b_24')
// (17, 18, 'sp4_r_v_b_8')
// (17, 18, 'sp4_v_b_9')
// (17, 18, 'sp4_v_t_37')
// (17, 19, 'sp4_r_v_b_13')
// (17, 19, 'sp4_r_v_b_46')
// (17, 19, 'sp4_v_b_37')
// (17, 20, 'sp4_r_v_b_0')
// (17, 20, 'sp4_r_v_b_35')
// (17, 20, 'sp4_v_b_24')
// (17, 21, 'local_g1_5')
// (17, 21, 'lutff_6/in_0')
// (17, 21, 'sp4_r_v_b_22')
// (17, 21, 'sp4_v_b_13')
// (17, 22, 'local_g1_0')
// (17, 22, 'lutff_5/in_2')
// (17, 22, 'sp4_r_v_b_11')
// (17, 22, 'sp4_v_b_0')
// (18, 14, 'sp4_v_t_45')
// (18, 15, 'sp4_v_b_45')
// (18, 16, 'neigh_op_tnl_2')
// (18, 16, 'sp4_v_b_32')
// (18, 16, 'sp4_v_t_37')
// (18, 17, 'local_g0_2')
// (18, 17, 'lutff_6/in_2')
// (18, 17, 'neigh_op_lft_2')
// (18, 17, 'sp4_h_r_17')
// (18, 17, 'sp4_v_b_21')
// (18, 17, 'sp4_v_b_37')
// (18, 18, 'local_g2_2')
// (18, 18, 'lutff_1/in_1')
// (18, 18, 'neigh_op_bnl_2')
// (18, 18, 'sp4_h_r_2')
// (18, 18, 'sp4_v_b_24')
// (18, 18, 'sp4_v_b_8')
// (18, 18, 'sp4_v_t_46')
// (18, 19, 'local_g0_5')
// (18, 19, 'lutff_5/in_0')
// (18, 19, 'sp4_v_b_13')
// (18, 19, 'sp4_v_b_46')
// (18, 20, 'sp4_v_b_0')
// (18, 20, 'sp4_v_b_35')
// (18, 21, 'sp4_v_b_22')
// (18, 22, 'local_g0_3')
// (18, 22, 'lutff_1/in_2')
// (18, 22, 'lutff_2/in_3')
// (18, 22, 'sp4_v_b_11')
// (19, 17, 'sp4_h_r_28')
// (19, 18, 'sp4_h_r_15')
// (20, 14, 'sp4_r_v_b_47')
// (20, 15, 'sp4_r_v_b_34')
// (20, 16, 'sp4_r_v_b_23')
// (20, 17, 'local_g2_1')
// (20, 17, 'lutff_5/in_0')
// (20, 17, 'sp4_h_r_41')
// (20, 17, 'sp4_r_v_b_10')
// (20, 18, 'local_g3_2')
// (20, 18, 'lutff_3/in_0')
// (20, 18, 'lutff_4/in_3')
// (20, 18, 'sp4_h_r_26')
// (20, 18, 'sp4_r_v_b_41')
// (20, 18, 'sp4_r_v_b_44')
// (20, 19, 'sp4_r_v_b_28')
// (20, 19, 'sp4_r_v_b_33')
// (20, 20, 'local_g3_4')
// (20, 20, 'lutff_5/in_0')
// (20, 20, 'sp4_r_v_b_17')
// (20, 20, 'sp4_r_v_b_20')
// (20, 21, 'local_g2_1')
// (20, 21, 'lutff_7/in_0')
// (20, 21, 'sp4_r_v_b_4')
// (20, 21, 'sp4_r_v_b_9')
// (21, 13, 'sp4_v_t_47')
// (21, 14, 'sp4_v_b_47')
// (21, 15, 'sp4_v_b_34')
// (21, 16, 'local_g1_7')
// (21, 16, 'lutff_0/in_0')
// (21, 16, 'sp4_v_b_23')
// (21, 17, 'local_g0_0')
// (21, 17, 'lutff_4/in_2')
// (21, 17, 'lutff_5/in_1')
// (21, 17, 'sp4_h_l_41')
// (21, 17, 'sp4_h_r_0')
// (21, 17, 'sp4_v_b_10')
// (21, 17, 'sp4_v_t_41')
// (21, 17, 'sp4_v_t_44')
// (21, 18, 'sp4_h_r_39')
// (21, 18, 'sp4_v_b_41')
// (21, 18, 'sp4_v_b_44')
// (21, 19, 'sp4_v_b_28')
// (21, 19, 'sp4_v_b_33')
// (21, 20, 'local_g0_1')
// (21, 20, 'lutff_7/in_0')
// (21, 20, 'sp4_v_b_17')
// (21, 20, 'sp4_v_b_20')
// (21, 21, 'local_g1_1')
// (21, 21, 'lutff_1/in_3')
// (21, 21, 'lutff_4/in_0')
// (21, 21, 'lutff_7/in_3')
// (21, 21, 'sp4_h_r_3')
// (21, 21, 'sp4_v_b_4')
// (21, 21, 'sp4_v_b_9')
// (22, 17, 'sp4_h_r_13')
// (22, 18, 'local_g0_5')
// (22, 18, 'lutff_2/in_3')
// (22, 18, 'lutff_7/in_2')
// (22, 18, 'sp4_h_l_39')
// (22, 18, 'sp4_h_r_5')
// (22, 21, 'local_g0_6')
// (22, 21, 'lutff_4/in_2')
// (22, 21, 'sp4_h_r_14')
// (23, 17, 'sp4_h_r_24')
// (23, 18, 'sp4_h_r_16')
// (23, 21, 'sp4_h_r_27')
// (24, 17, 'sp4_h_r_37')
// (24, 18, 'sp4_h_r_29')
// (24, 21, 'sp4_h_r_38')
// (25, 17, 'sp4_h_l_37')
// (25, 18, 'sp4_h_r_40')
// (25, 21, 'sp4_h_l_38')

reg n2404 = 0;
// (16, 15, 'sp4_r_v_b_46')
// (16, 16, 'neigh_op_tnr_3')
// (16, 16, 'sp4_r_v_b_35')
// (16, 17, 'neigh_op_rgt_3')
// (16, 17, 'sp4_h_r_11')
// (16, 17, 'sp4_r_v_b_22')
// (16, 18, 'neigh_op_bnr_3')
// (16, 18, 'sp4_r_v_b_11')
// (16, 19, 'sp4_r_v_b_42')
// (16, 20, 'sp4_r_v_b_31')
// (16, 21, 'sp4_r_v_b_18')
// (16, 22, 'sp4_r_v_b_7')
// (17, 14, 'sp4_v_t_46')
// (17, 15, 'sp4_r_v_b_47')
// (17, 15, 'sp4_v_b_46')
// (17, 16, 'neigh_op_top_3')
// (17, 16, 'sp4_r_v_b_34')
// (17, 16, 'sp4_v_b_35')
// (17, 17, 'lutff_3/out')
// (17, 17, 'sp4_h_r_22')
// (17, 17, 'sp4_h_r_6')
// (17, 17, 'sp4_r_v_b_23')
// (17, 17, 'sp4_r_v_b_39')
// (17, 17, 'sp4_v_b_22')
// (17, 18, 'local_g0_3')
// (17, 18, 'lutff_6/in_3')
// (17, 18, 'neigh_op_bot_3')
// (17, 18, 'sp4_r_v_b_10')
// (17, 18, 'sp4_r_v_b_26')
// (17, 18, 'sp4_v_b_11')
// (17, 18, 'sp4_v_t_42')
// (17, 19, 'sp4_r_v_b_15')
// (17, 19, 'sp4_r_v_b_36')
// (17, 19, 'sp4_v_b_42')
// (17, 20, 'sp4_r_v_b_2')
// (17, 20, 'sp4_r_v_b_25')
// (17, 20, 'sp4_v_b_31')
// (17, 21, 'sp4_r_v_b_12')
// (17, 21, 'sp4_r_v_b_39')
// (17, 21, 'sp4_v_b_18')
// (17, 22, 'local_g1_7')
// (17, 22, 'lutff_5/in_3')
// (17, 22, 'sp4_r_v_b_1')
// (17, 22, 'sp4_r_v_b_26')
// (17, 22, 'sp4_v_b_7')
// (17, 23, 'sp4_r_v_b_15')
// (17, 24, 'sp4_r_v_b_2')
// (18, 14, 'sp4_v_t_47')
// (18, 15, 'sp4_v_b_47')
// (18, 16, 'neigh_op_tnl_3')
// (18, 16, 'sp4_h_r_7')
// (18, 16, 'sp4_v_b_34')
// (18, 16, 'sp4_v_t_39')
// (18, 17, 'local_g1_3')
// (18, 17, 'lutff_2/in_0')
// (18, 17, 'neigh_op_lft_3')
// (18, 17, 'sp4_h_r_19')
// (18, 17, 'sp4_h_r_35')
// (18, 17, 'sp4_v_b_23')
// (18, 17, 'sp4_v_b_39')
// (18, 18, 'local_g3_3')
// (18, 18, 'lutff_1/in_3')
// (18, 18, 'lutff_6/in_0')
// (18, 18, 'neigh_op_bnl_3')
// (18, 18, 'sp4_h_r_10')
// (18, 18, 'sp4_v_b_10')
// (18, 18, 'sp4_v_b_26')
// (18, 18, 'sp4_v_t_36')
// (18, 19, 'local_g1_7')
// (18, 19, 'lutff_5/in_1')
// (18, 19, 'sp4_v_b_15')
// (18, 19, 'sp4_v_b_36')
// (18, 20, 'sp4_v_b_2')
// (18, 20, 'sp4_v_b_25')
// (18, 20, 'sp4_v_t_39')
// (18, 21, 'local_g0_4')
// (18, 21, 'lutff_1/in_3')
// (18, 21, 'sp4_v_b_12')
// (18, 21, 'sp4_v_b_39')
// (18, 22, 'local_g2_2')
// (18, 22, 'lutff_1/in_3')
// (18, 22, 'lutff_2/in_2')
// (18, 22, 'sp4_h_r_1')
// (18, 22, 'sp4_v_b_1')
// (18, 22, 'sp4_v_b_26')
// (18, 23, 'sp4_v_b_15')
// (18, 24, 'sp4_v_b_2')
// (19, 16, 'sp4_h_r_18')
// (19, 17, 'sp4_h_r_30')
// (19, 17, 'sp4_h_r_46')
// (19, 18, 'sp4_h_r_23')
// (19, 22, 'sp4_h_r_12')
// (20, 14, 'sp4_r_v_b_37')
// (20, 15, 'sp4_r_v_b_24')
// (20, 16, 'sp4_h_r_31')
// (20, 16, 'sp4_r_v_b_13')
// (20, 17, 'sp4_h_l_46')
// (20, 17, 'sp4_h_r_43')
// (20, 17, 'sp4_h_r_7')
// (20, 17, 'sp4_r_v_b_0')
// (20, 18, 'local_g2_2')
// (20, 18, 'lutff_3/in_1')
// (20, 18, 'lutff_4/in_0')
// (20, 18, 'sp4_h_r_34')
// (20, 18, 'sp4_r_v_b_43')
// (20, 18, 'sp4_r_v_b_46')
// (20, 19, 'sp4_r_v_b_30')
// (20, 19, 'sp4_r_v_b_35')
// (20, 20, 'local_g3_3')
// (20, 20, 'lutff_5/in_1')
// (20, 20, 'sp4_r_v_b_19')
// (20, 20, 'sp4_r_v_b_22')
// (20, 21, 'local_g1_6')
// (20, 21, 'lutff_3/in_0')
// (20, 21, 'sp4_r_v_b_11')
// (20, 21, 'sp4_r_v_b_6')
// (20, 22, 'local_g3_1')
// (20, 22, 'lutff_5/in_1')
// (20, 22, 'lutff_7/in_1')
// (20, 22, 'sp4_h_r_25')
// (21, 13, 'sp4_v_t_37')
// (21, 14, 'sp4_v_b_37')
// (21, 15, 'sp4_v_b_24')
// (21, 16, 'local_g0_5')
// (21, 16, 'local_g1_5')
// (21, 16, 'lutff_1/in_2')
// (21, 16, 'lutff_3/in_3')
// (21, 16, 'lutff_4/in_0')
// (21, 16, 'sp4_h_r_42')
// (21, 16, 'sp4_v_b_13')
// (21, 17, 'local_g0_2')
// (21, 17, 'local_g1_6')
// (21, 17, 'lutff_4/in_1')
// (21, 17, 'lutff_5/in_3')
// (21, 17, 'sp4_h_l_43')
// (21, 17, 'sp4_h_r_18')
// (21, 17, 'sp4_h_r_2')
// (21, 17, 'sp4_h_r_6')
// (21, 17, 'sp4_v_b_0')
// (21, 17, 'sp4_v_t_43')
// (21, 17, 'sp4_v_t_46')
// (21, 18, 'sp4_h_r_47')
// (21, 18, 'sp4_v_b_43')
// (21, 18, 'sp4_v_b_46')
// (21, 19, 'sp4_v_b_30')
// (21, 19, 'sp4_v_b_35')
// (21, 20, 'local_g1_6')
// (21, 20, 'lutff_2/in_3')
// (21, 20, 'lutff_4/in_3')
// (21, 20, 'sp4_v_b_19')
// (21, 20, 'sp4_v_b_22')
// (21, 21, 'local_g0_6')
// (21, 21, 'local_g1_6')
// (21, 21, 'lutff_2/in_0')
// (21, 21, 'lutff_4/in_3')
// (21, 21, 'lutff_5/in_3')
// (21, 21, 'sp4_v_b_11')
// (21, 21, 'sp4_v_b_6')
// (21, 22, 'sp4_h_r_36')
// (22, 16, 'local_g1_7')
// (22, 16, 'lutff_2/in_0')
// (22, 16, 'sp4_h_l_42')
// (22, 16, 'sp4_h_r_7')
// (22, 17, 'sp4_h_r_15')
// (22, 17, 'sp4_h_r_19')
// (22, 17, 'sp4_h_r_31')
// (22, 18, 'local_g0_2')
// (22, 18, 'lutff_2/in_0')
// (22, 18, 'lutff_7/in_1')
// (22, 18, 'sp4_h_l_47')
// (22, 18, 'sp4_h_r_10')
// (22, 22, 'sp4_h_l_36')
// (23, 16, 'sp4_h_r_18')
// (23, 17, 'local_g2_6')
// (23, 17, 'lutff_7/in_1')
// (23, 17, 'sp4_h_r_26')
// (23, 17, 'sp4_h_r_30')
// (23, 17, 'sp4_h_r_42')
// (23, 18, 'sp4_h_r_23')
// (23, 18, 'sp4_r_v_b_37')
// (23, 19, 'local_g1_0')
// (23, 19, 'lutff_1/in_0')
// (23, 19, 'sp4_r_v_b_24')
// (23, 20, 'sp4_r_v_b_13')
// (23, 21, 'sp4_r_v_b_0')
// (24, 16, 'sp4_h_r_31')
// (24, 17, 'sp4_h_l_42')
// (24, 17, 'sp4_h_r_39')
// (24, 17, 'sp4_h_r_43')
// (24, 17, 'sp4_v_t_37')
// (24, 18, 'sp4_h_r_34')
// (24, 18, 'sp4_v_b_37')
// (24, 19, 'sp4_v_b_24')
// (24, 20, 'sp4_v_b_13')
// (24, 21, 'sp4_v_b_0')
// (25, 16, 'sp4_h_r_42')
// (25, 17, 'sp4_h_l_39')
// (25, 17, 'sp4_h_l_43')
// (25, 18, 'sp4_h_r_47')

reg n2405 = 0;
// (16, 16, 'neigh_op_tnr_1')
// (16, 17, 'neigh_op_rgt_1')
// (16, 18, 'neigh_op_bnr_1')
// (17, 15, 'sp4_r_v_b_43')
// (17, 16, 'neigh_op_top_1')
// (17, 16, 'sp4_r_v_b_30')
// (17, 17, 'lutff_1/out')
// (17, 17, 'sp4_r_v_b_19')
// (17, 18, 'neigh_op_bot_1')
// (17, 18, 'sp4_r_v_b_6')
// (18, 14, 'sp4_v_t_43')
// (18, 15, 'sp4_v_b_43')
// (18, 16, 'neigh_op_tnl_1')
// (18, 16, 'sp4_v_b_30')
// (18, 17, 'neigh_op_lft_1')
// (18, 17, 'sp4_v_b_19')
// (18, 18, 'neigh_op_bnl_1')
// (18, 18, 'sp4_h_r_6')
// (18, 18, 'sp4_v_b_6')
// (19, 18, 'sp4_h_r_19')
// (20, 18, 'local_g2_6')
// (20, 18, 'lutff_0/in_0')
// (20, 18, 'sp4_h_r_30')
// (21, 18, 'sp4_h_r_43')
// (22, 18, 'sp4_h_l_43')

reg n2406 = 0;
// (16, 16, 'neigh_op_tnr_4')
// (16, 17, 'neigh_op_rgt_4')
// (16, 17, 'sp4_r_v_b_40')
// (16, 18, 'neigh_op_bnr_4')
// (16, 18, 'sp4_r_v_b_29')
// (16, 19, 'sp4_r_v_b_16')
// (16, 20, 'sp4_r_v_b_5')
// (17, 9, 'sp12_v_t_23')
// (17, 10, 'sp12_v_b_23')
// (17, 11, 'sp12_v_b_20')
// (17, 12, 'sp12_v_b_19')
// (17, 13, 'sp12_v_b_16')
// (17, 14, 'sp12_v_b_15')
// (17, 15, 'sp12_v_b_12')
// (17, 16, 'neigh_op_top_4')
// (17, 16, 'sp12_v_b_11')
// (17, 16, 'sp4_v_t_40')
// (17, 17, 'lutff_4/out')
// (17, 17, 'sp12_v_b_8')
// (17, 17, 'sp4_h_r_8')
// (17, 17, 'sp4_r_v_b_41')
// (17, 17, 'sp4_v_b_40')
// (17, 18, 'neigh_op_bot_4')
// (17, 18, 'sp12_v_b_7')
// (17, 18, 'sp4_r_v_b_28')
// (17, 18, 'sp4_v_b_29')
// (17, 19, 'sp12_v_b_4')
// (17, 19, 'sp4_r_v_b_17')
// (17, 19, 'sp4_v_b_16')
// (17, 20, 'sp12_v_b_3')
// (17, 20, 'sp4_h_r_5')
// (17, 20, 'sp4_r_v_b_4')
// (17, 20, 'sp4_v_b_5')
// (17, 21, 'local_g3_0')
// (17, 21, 'lutff_6/in_3')
// (17, 21, 'sp12_v_b_0')
// (18, 16, 'neigh_op_tnl_4')
// (18, 16, 'sp4_h_r_9')
// (18, 16, 'sp4_v_t_41')
// (18, 17, 'local_g1_4')
// (18, 17, 'lutff_6/in_1')
// (18, 17, 'neigh_op_lft_4')
// (18, 17, 'sp4_h_r_21')
// (18, 17, 'sp4_v_b_41')
// (18, 18, 'local_g2_4')
// (18, 18, 'lutff_7/in_1')
// (18, 18, 'neigh_op_bnl_4')
// (18, 18, 'sp4_v_b_28')
// (18, 19, 'sp4_v_b_17')
// (18, 20, 'sp4_h_r_16')
// (18, 20, 'sp4_v_b_4')
// (19, 16, 'sp4_h_r_20')
// (19, 17, 'sp4_h_r_32')
// (19, 20, 'sp4_h_r_29')
// (20, 14, 'sp4_r_v_b_39')
// (20, 15, 'sp4_r_v_b_26')
// (20, 16, 'sp4_h_r_33')
// (20, 16, 'sp4_r_v_b_15')
// (20, 17, 'local_g2_5')
// (20, 17, 'lutff_5/in_2')
// (20, 17, 'sp4_h_r_45')
// (20, 17, 'sp4_r_v_b_2')
// (20, 18, 'local_g3_5')
// (20, 18, 'lutff_6/in_2')
// (20, 18, 'lutff_7/in_1')
// (20, 18, 'sp4_r_v_b_45')
// (20, 19, 'sp4_r_v_b_32')
// (20, 20, 'local_g2_0')
// (20, 20, 'lutff_3/in_3')
// (20, 20, 'lutff_7/in_3')
// (20, 20, 'sp4_h_r_40')
// (20, 20, 'sp4_r_v_b_21')
// (20, 21, 'local_g2_0')
// (20, 21, 'lutff_7/in_3')
// (20, 21, 'sp4_r_v_b_8')
// (21, 13, 'sp4_v_t_39')
// (21, 14, 'sp4_v_b_39')
// (21, 15, 'sp4_v_b_26')
// (21, 16, 'local_g0_7')
// (21, 16, 'lutff_1/in_0')
// (21, 16, 'lutff_4/in_3')
// (21, 16, 'sp4_h_r_44')
// (21, 16, 'sp4_v_b_15')
// (21, 17, 'local_g1_3')
// (21, 17, 'lutff_3/in_1')
// (21, 17, 'sp4_h_l_45')
// (21, 17, 'sp4_h_r_11')
// (21, 17, 'sp4_v_b_2')
// (21, 17, 'sp4_v_t_45')
// (21, 18, 'local_g2_5')
// (21, 18, 'lutff_3/in_0')
// (21, 18, 'sp4_v_b_45')
// (21, 19, 'sp4_v_b_32')
// (21, 20, 'local_g1_5')
// (21, 20, 'lutff_7/in_3')
// (21, 20, 'sp4_h_l_40')
// (21, 20, 'sp4_v_b_21')
// (21, 21, 'local_g0_0')
// (21, 21, 'local_g1_0')
// (21, 21, 'lutff_1/in_1')
// (21, 21, 'lutff_7/in_0')
// (21, 21, 'sp4_h_r_2')
// (21, 21, 'sp4_v_b_8')
// (22, 16, 'local_g1_0')
// (22, 16, 'lutff_2/in_3')
// (22, 16, 'sp4_h_l_44')
// (22, 16, 'sp4_h_r_0')
// (22, 17, 'sp4_h_r_22')
// (22, 21, 'local_g0_7')
// (22, 21, 'lutff_4/in_1')
// (22, 21, 'sp4_h_r_15')
// (23, 16, 'sp4_h_r_13')
// (23, 17, 'sp4_h_r_35')
// (23, 21, 'sp4_h_r_26')
// (24, 16, 'sp4_h_r_24')
// (24, 17, 'sp4_h_r_46')
// (24, 21, 'sp4_h_r_39')
// (25, 16, 'sp4_h_r_37')
// (25, 17, 'sp4_h_l_46')
// (25, 21, 'sp4_h_l_39')

reg n2407 = 0;
// (16, 16, 'neigh_op_tnr_5')
// (16, 16, 'sp4_r_v_b_39')
// (16, 17, 'neigh_op_rgt_5')
// (16, 17, 'sp4_r_v_b_26')
// (16, 18, 'neigh_op_bnr_5')
// (16, 18, 'sp4_r_v_b_15')
// (16, 19, 'sp4_r_v_b_2')
// (17, 15, 'sp4_v_t_39')
// (17, 16, 'neigh_op_top_5')
// (17, 16, 'sp4_r_v_b_38')
// (17, 16, 'sp4_v_b_39')
// (17, 17, 'lutff_5/out')
// (17, 17, 'sp4_r_v_b_27')
// (17, 17, 'sp4_v_b_26')
// (17, 18, 'neigh_op_bot_5')
// (17, 18, 'sp4_r_v_b_14')
// (17, 18, 'sp4_v_b_15')
// (17, 19, 'sp4_h_r_2')
// (17, 19, 'sp4_r_v_b_3')
// (17, 19, 'sp4_v_b_2')
// (18, 15, 'sp4_v_t_38')
// (18, 16, 'neigh_op_tnl_5')
// (18, 16, 'sp4_v_b_38')
// (18, 17, 'neigh_op_lft_5')
// (18, 17, 'sp4_v_b_27')
// (18, 18, 'neigh_op_bnl_5')
// (18, 18, 'sp4_v_b_14')
// (18, 19, 'sp4_h_r_15')
// (18, 19, 'sp4_h_r_3')
// (18, 19, 'sp4_v_b_3')
// (19, 19, 'sp4_h_r_14')
// (19, 19, 'sp4_h_r_26')
// (20, 16, 'sp4_r_v_b_39')
// (20, 17, 'sp4_r_v_b_26')
// (20, 18, 'local_g2_7')
// (20, 18, 'lutff_1/in_0')
// (20, 18, 'sp4_r_v_b_15')
// (20, 19, 'local_g3_3')
// (20, 19, 'lutff_1/in_3')
// (20, 19, 'sp4_h_r_27')
// (20, 19, 'sp4_h_r_39')
// (20, 19, 'sp4_r_v_b_2')
// (21, 15, 'sp4_v_t_39')
// (21, 16, 'sp4_v_b_39')
// (21, 17, 'sp4_v_b_26')
// (21, 18, 'sp4_v_b_15')
// (21, 19, 'sp4_h_l_39')
// (21, 19, 'sp4_h_r_38')
// (21, 19, 'sp4_v_b_2')
// (22, 19, 'sp4_h_l_38')

reg n2408 = 0;
// (16, 16, 'neigh_op_tnr_7')
// (16, 17, 'neigh_op_rgt_7')
// (16, 17, 'sp4_h_r_3')
// (16, 18, 'neigh_op_bnr_7')
// (17, 16, 'neigh_op_top_7')
// (17, 17, 'lutff_7/out')
// (17, 17, 'sp4_h_r_14')
// (17, 18, 'neigh_op_bot_7')
// (18, 16, 'neigh_op_tnl_7')
// (18, 17, 'neigh_op_lft_7')
// (18, 17, 'sp4_h_r_27')
// (18, 18, 'local_g2_7')
// (18, 18, 'lutff_7/in_0')
// (18, 18, 'neigh_op_bnl_7')
// (19, 17, 'sp4_h_r_38')
// (19, 18, 'sp4_r_v_b_38')
// (19, 18, 'sp4_r_v_b_45')
// (19, 19, 'sp4_r_v_b_27')
// (19, 19, 'sp4_r_v_b_32')
// (19, 20, 'sp4_r_v_b_14')
// (19, 20, 'sp4_r_v_b_21')
// (19, 21, 'sp4_r_v_b_3')
// (19, 21, 'sp4_r_v_b_8')
// (20, 17, 'local_g0_6')
// (20, 17, 'lutff_0/in_2')
// (20, 17, 'sp4_h_l_38')
// (20, 17, 'sp4_h_r_3')
// (20, 17, 'sp4_h_r_6')
// (20, 17, 'sp4_v_t_38')
// (20, 17, 'sp4_v_t_45')
// (20, 18, 'sp4_v_b_38')
// (20, 18, 'sp4_v_b_45')
// (20, 19, 'sp4_v_b_27')
// (20, 19, 'sp4_v_b_32')
// (20, 20, 'local_g1_5')
// (20, 20, 'local_g1_6')
// (20, 20, 'lutff_1/in_0')
// (20, 20, 'lutff_3/in_0')
// (20, 20, 'lutff_7/in_1')
// (20, 20, 'sp4_v_b_14')
// (20, 20, 'sp4_v_b_21')
// (20, 21, 'sp4_h_r_2')
// (20, 21, 'sp4_v_b_3')
// (20, 21, 'sp4_v_b_8')
// (21, 17, 'local_g0_6')
// (21, 17, 'lutff_3/in_3')
// (21, 17, 'sp4_h_r_14')
// (21, 17, 'sp4_h_r_19')
// (21, 21, 'local_g1_7')
// (21, 21, 'lutff_2/in_2')
// (21, 21, 'sp4_h_r_15')
// (22, 17, 'sp4_h_r_27')
// (22, 17, 'sp4_h_r_30')
// (22, 21, 'sp4_h_r_26')
// (23, 17, 'sp4_h_r_38')
// (23, 17, 'sp4_h_r_43')
// (23, 21, 'sp4_h_r_39')
// (24, 17, 'sp4_h_l_38')
// (24, 17, 'sp4_h_l_43')
// (24, 21, 'sp4_h_l_39')

reg n2409 = 0;
// (16, 17, 'neigh_op_tnr_1')
// (16, 18, 'neigh_op_rgt_1')
// (16, 19, 'neigh_op_bnr_1')
// (17, 15, 'sp4_r_v_b_38')
// (17, 16, 'sp4_r_v_b_27')
// (17, 17, 'local_g1_1')
// (17, 17, 'lutff_4/in_2')
// (17, 17, 'neigh_op_top_1')
// (17, 17, 'sp4_r_v_b_14')
// (17, 17, 'sp4_r_v_b_46')
// (17, 18, 'local_g0_1')
// (17, 18, 'lutff_1/in_2')
// (17, 18, 'lutff_1/out')
// (17, 18, 'sp4_r_v_b_3')
// (17, 18, 'sp4_r_v_b_35')
// (17, 19, 'neigh_op_bot_1')
// (17, 19, 'sp4_r_v_b_22')
// (17, 20, 'local_g2_3')
// (17, 20, 'lutff_1/in_0')
// (17, 20, 'sp4_r_v_b_11')
// (18, 14, 'sp4_v_t_38')
// (18, 15, 'sp4_v_b_38')
// (18, 16, 'local_g2_3')
// (18, 16, 'lutff_3/in_0')
// (18, 16, 'sp4_v_b_27')
// (18, 16, 'sp4_v_t_46')
// (18, 17, 'neigh_op_tnl_1')
// (18, 17, 'sp4_v_b_14')
// (18, 17, 'sp4_v_b_46')
// (18, 18, 'neigh_op_lft_1')
// (18, 18, 'sp4_v_b_3')
// (18, 18, 'sp4_v_b_35')
// (18, 19, 'neigh_op_bnl_1')
// (18, 19, 'sp4_v_b_22')
// (18, 20, 'sp4_v_b_11')

reg n2410 = 0;
// (16, 17, 'neigh_op_tnr_2')
// (16, 18, 'neigh_op_rgt_2')
// (16, 18, 'sp4_r_v_b_36')
// (16, 19, 'neigh_op_bnr_2')
// (16, 19, 'sp4_r_v_b_25')
// (16, 20, 'sp4_r_v_b_12')
// (16, 21, 'sp4_r_v_b_1')
// (17, 15, 'sp4_r_v_b_40')
// (17, 16, 'sp4_r_v_b_29')
// (17, 17, 'local_g1_2')
// (17, 17, 'lutff_3/in_0')
// (17, 17, 'neigh_op_top_2')
// (17, 17, 'sp4_r_v_b_16')
// (17, 17, 'sp4_v_t_36')
// (17, 18, 'local_g2_2')
// (17, 18, 'lutff_2/in_2')
// (17, 18, 'lutff_2/out')
// (17, 18, 'sp4_r_v_b_5')
// (17, 18, 'sp4_v_b_36')
// (17, 19, 'neigh_op_bot_2')
// (17, 19, 'sp4_v_b_25')
// (17, 20, 'local_g0_4')
// (17, 20, 'lutff_3/in_3')
// (17, 20, 'sp4_v_b_12')
// (17, 21, 'sp4_v_b_1')
// (18, 14, 'sp4_v_t_40')
// (18, 15, 'sp4_v_b_40')
// (18, 16, 'local_g2_5')
// (18, 16, 'lutff_6/in_1')
// (18, 16, 'sp4_v_b_29')
// (18, 17, 'neigh_op_tnl_2')
// (18, 17, 'sp4_v_b_16')
// (18, 18, 'neigh_op_lft_2')
// (18, 18, 'sp4_v_b_5')
// (18, 19, 'neigh_op_bnl_2')

reg n2411 = 0;
// (16, 17, 'neigh_op_tnr_3')
// (16, 18, 'neigh_op_rgt_3')
// (16, 18, 'sp4_r_v_b_38')
// (16, 19, 'neigh_op_bnr_3')
// (16, 19, 'sp4_r_v_b_27')
// (16, 20, 'sp4_r_v_b_14')
// (16, 21, 'sp4_r_v_b_3')
// (17, 15, 'sp4_r_v_b_42')
// (17, 16, 'sp4_r_v_b_31')
// (17, 17, 'local_g1_3')
// (17, 17, 'lutff_5/in_1')
// (17, 17, 'neigh_op_top_3')
// (17, 17, 'sp4_r_v_b_18')
// (17, 17, 'sp4_v_t_38')
// (17, 18, 'local_g3_3')
// (17, 18, 'lutff_3/in_1')
// (17, 18, 'lutff_3/out')
// (17, 18, 'sp4_r_v_b_7')
// (17, 18, 'sp4_v_b_38')
// (17, 19, 'neigh_op_bot_3')
// (17, 19, 'sp4_v_b_27')
// (17, 20, 'local_g0_6')
// (17, 20, 'lutff_2/in_2')
// (17, 20, 'sp4_v_b_14')
// (17, 21, 'sp4_v_b_3')
// (18, 14, 'sp4_v_t_42')
// (18, 15, 'sp4_v_b_42')
// (18, 16, 'local_g3_7')
// (18, 16, 'lutff_1/in_1')
// (18, 16, 'sp4_v_b_31')
// (18, 17, 'neigh_op_tnl_3')
// (18, 17, 'sp4_v_b_18')
// (18, 18, 'neigh_op_lft_3')
// (18, 18, 'sp4_v_b_7')
// (18, 19, 'neigh_op_bnl_3')

reg n2412 = 0;
// (16, 17, 'neigh_op_tnr_4')
// (16, 17, 'sp4_r_v_b_37')
// (16, 18, 'neigh_op_rgt_4')
// (16, 18, 'sp4_r_v_b_24')
// (16, 19, 'neigh_op_bnr_4')
// (16, 19, 'sp4_r_v_b_13')
// (16, 20, 'sp4_r_v_b_0')
// (17, 15, 'sp4_r_v_b_44')
// (17, 16, 'sp4_r_v_b_33')
// (17, 16, 'sp4_v_t_37')
// (17, 17, 'local_g0_4')
// (17, 17, 'lutff_1/in_1')
// (17, 17, 'neigh_op_top_4')
// (17, 17, 'sp4_r_v_b_20')
// (17, 17, 'sp4_v_b_37')
// (17, 18, 'local_g0_4')
// (17, 18, 'lutff_4/in_2')
// (17, 18, 'lutff_4/out')
// (17, 18, 'sp4_r_v_b_9')
// (17, 18, 'sp4_v_b_24')
// (17, 19, 'neigh_op_bot_4')
// (17, 19, 'sp4_v_b_13')
// (17, 20, 'local_g0_0')
// (17, 20, 'lutff_7/in_1')
// (17, 20, 'sp4_v_b_0')
// (18, 14, 'sp4_v_t_44')
// (18, 15, 'sp4_v_b_44')
// (18, 16, 'local_g3_1')
// (18, 16, 'lutff_4/in_0')
// (18, 16, 'sp4_v_b_33')
// (18, 17, 'neigh_op_tnl_4')
// (18, 17, 'sp4_v_b_20')
// (18, 18, 'neigh_op_lft_4')
// (18, 18, 'sp4_v_b_9')
// (18, 19, 'neigh_op_bnl_4')

reg n2413 = 0;
// (16, 17, 'neigh_op_tnr_5')
// (16, 18, 'neigh_op_rgt_5')
// (16, 19, 'neigh_op_bnr_5')
// (17, 15, 'sp4_r_v_b_46')
// (17, 16, 'sp4_r_v_b_35')
// (17, 17, 'local_g1_5')
// (17, 17, 'lutff_7/in_1')
// (17, 17, 'neigh_op_top_5')
// (17, 17, 'sp4_r_v_b_22')
// (17, 17, 'sp4_r_v_b_38')
// (17, 18, 'local_g3_5')
// (17, 18, 'lutff_5/in_1')
// (17, 18, 'lutff_5/out')
// (17, 18, 'sp4_r_v_b_11')
// (17, 18, 'sp4_r_v_b_27')
// (17, 19, 'neigh_op_bot_5')
// (17, 19, 'sp4_r_v_b_14')
// (17, 20, 'local_g1_3')
// (17, 20, 'lutff_0/in_0')
// (17, 20, 'sp4_r_v_b_3')
// (18, 14, 'sp4_v_t_46')
// (18, 15, 'sp4_v_b_46')
// (18, 16, 'local_g3_3')
// (18, 16, 'lutff_0/in_0')
// (18, 16, 'sp4_v_b_35')
// (18, 16, 'sp4_v_t_38')
// (18, 17, 'neigh_op_tnl_5')
// (18, 17, 'sp4_v_b_22')
// (18, 17, 'sp4_v_b_38')
// (18, 18, 'neigh_op_lft_5')
// (18, 18, 'sp4_v_b_11')
// (18, 18, 'sp4_v_b_27')
// (18, 19, 'neigh_op_bnl_5')
// (18, 19, 'sp4_v_b_14')
// (18, 20, 'sp4_v_b_3')

wire n2414;
// (16, 17, 'neigh_op_tnr_6')
// (16, 18, 'neigh_op_rgt_6')
// (16, 18, 'sp4_h_r_1')
// (16, 19, 'neigh_op_bnr_6')
// (17, 17, 'neigh_op_top_6')
// (17, 18, 'lutff_6/out')
// (17, 18, 'sp4_h_r_12')
// (17, 19, 'neigh_op_bot_6')
// (18, 17, 'neigh_op_tnl_6')
// (18, 18, 'neigh_op_lft_6')
// (18, 18, 'sp4_h_r_25')
// (18, 19, 'neigh_op_bnl_6')
// (19, 18, 'sp4_h_r_36')
// (20, 18, 'local_g1_4')
// (20, 18, 'lutff_6/in_3')
// (20, 18, 'sp4_h_l_36')
// (20, 18, 'sp4_h_r_4')
// (21, 18, 'sp4_h_r_17')
// (22, 18, 'sp4_h_r_28')
// (23, 18, 'sp4_h_r_41')
// (24, 18, 'sp4_h_l_41')

reg n2415 = 0;
// (16, 17, 'neigh_op_tnr_7')
// (16, 18, 'neigh_op_rgt_7')
// (16, 19, 'neigh_op_bnr_7')
// (17, 16, 'sp4_r_v_b_39')
// (17, 17, 'local_g1_7')
// (17, 17, 'lutff_2/in_0')
// (17, 17, 'neigh_op_top_7')
// (17, 17, 'sp4_r_v_b_26')
// (17, 17, 'sp4_r_v_b_42')
// (17, 18, 'local_g3_7')
// (17, 18, 'lutff_0/in_2')
// (17, 18, 'lutff_1/in_3')
// (17, 18, 'lutff_7/in_1')
// (17, 18, 'lutff_7/out')
// (17, 18, 'sp4_r_v_b_15')
// (17, 18, 'sp4_r_v_b_31')
// (17, 19, 'neigh_op_bot_7')
// (17, 19, 'sp4_r_v_b_18')
// (17, 19, 'sp4_r_v_b_2')
// (17, 20, 'local_g1_7')
// (17, 20, 'lutff_5/in_1')
// (17, 20, 'sp4_r_v_b_7')
// (18, 15, 'sp4_v_t_39')
// (18, 16, 'local_g2_7')
// (18, 16, 'lutff_5/in_0')
// (18, 16, 'sp4_v_b_39')
// (18, 16, 'sp4_v_t_42')
// (18, 17, 'neigh_op_tnl_7')
// (18, 17, 'sp4_v_b_26')
// (18, 17, 'sp4_v_b_42')
// (18, 18, 'neigh_op_lft_7')
// (18, 18, 'sp4_v_b_15')
// (18, 18, 'sp4_v_b_31')
// (18, 19, 'neigh_op_bnl_7')
// (18, 19, 'sp4_v_b_18')
// (18, 19, 'sp4_v_b_2')
// (18, 20, 'sp4_v_b_7')

wire n2416;
// (16, 18, 'lutff_1/cout')
// (16, 18, 'lutff_2/in_3')

wire n2417;
// (16, 18, 'lutff_3/cout')
// (16, 18, 'lutff_4/in_3')

wire n2418;
// (16, 18, 'lutff_5/cout')
// (16, 18, 'lutff_6/in_3')

wire n2419;
// (16, 18, 'lutff_7/cout')
// (16, 19, 'carry_in')
// (16, 19, 'carry_in_mux')
// (16, 19, 'lutff_0/in_3')

wire n2420;
// (16, 18, 'neigh_op_tnr_2')
// (16, 19, 'neigh_op_rgt_2')
// (16, 20, 'neigh_op_bnr_2')
// (17, 18, 'neigh_op_top_2')
// (17, 19, 'lutff_2/out')
// (17, 20, 'local_g1_2')
// (17, 20, 'lutff_3/in_2')
// (17, 20, 'neigh_op_bot_2')
// (18, 18, 'neigh_op_tnl_2')
// (18, 19, 'neigh_op_lft_2')
// (18, 20, 'neigh_op_bnl_2')

wire n2421;
// (16, 18, 'neigh_op_tnr_4')
// (16, 19, 'neigh_op_rgt_4')
// (16, 20, 'neigh_op_bnr_4')
// (17, 18, 'neigh_op_top_4')
// (17, 19, 'lutff_4/out')
// (17, 20, 'local_g1_4')
// (17, 20, 'lutff_2/in_3')
// (17, 20, 'neigh_op_bot_4')
// (18, 18, 'neigh_op_tnl_4')
// (18, 19, 'neigh_op_lft_4')
// (18, 20, 'neigh_op_bnl_4')

wire n2422;
// (16, 18, 'neigh_op_tnr_6')
// (16, 19, 'neigh_op_rgt_6')
// (16, 20, 'neigh_op_bnr_6')
// (17, 18, 'neigh_op_top_6')
// (17, 19, 'lutff_6/out')
// (17, 20, 'local_g1_6')
// (17, 20, 'lutff_7/in_2')
// (17, 20, 'neigh_op_bot_6')
// (18, 18, 'neigh_op_tnl_6')
// (18, 19, 'neigh_op_lft_6')
// (18, 20, 'neigh_op_bnl_6')

wire n2423;
// (16, 18, 'sp4_r_v_b_45')
// (16, 19, 'sp4_r_v_b_32')
// (16, 20, 'neigh_op_tnr_4')
// (16, 20, 'sp4_r_v_b_21')
// (16, 21, 'neigh_op_rgt_4')
// (16, 21, 'sp4_r_v_b_8')
// (16, 22, 'neigh_op_bnr_4')
// (17, 17, 'sp4_v_t_45')
// (17, 18, 'sp4_v_b_45')
// (17, 19, 'sp4_v_b_32')
// (17, 20, 'neigh_op_top_4')
// (17, 20, 'sp4_v_b_21')
// (17, 21, 'local_g0_2')
// (17, 21, 'lutff_4/out')
// (17, 21, 'lutff_global/cen')
// (17, 21, 'sp4_h_r_2')
// (17, 21, 'sp4_v_b_8')
// (17, 22, 'neigh_op_bot_4')
// (18, 20, 'neigh_op_tnl_4')
// (18, 21, 'neigh_op_lft_4')
// (18, 21, 'sp4_h_r_15')
// (18, 22, 'neigh_op_bnl_4')
// (19, 21, 'sp4_h_r_26')
// (20, 21, 'sp4_h_r_39')
// (21, 21, 'sp4_h_l_39')

wire n2424;
// (16, 19, 'lutff_1/cout')
// (16, 19, 'lutff_2/in_3')

wire n2425;
// (16, 19, 'lutff_3/cout')
// (16, 19, 'lutff_4/in_3')

reg n2426 = 0;
// (16, 19, 'neigh_op_tnr_3')
// (16, 20, 'neigh_op_rgt_3')
// (16, 21, 'neigh_op_bnr_3')
// (17, 18, 'sp4_r_v_b_47')
// (17, 19, 'local_g1_3')
// (17, 19, 'lutff_3/in_1')
// (17, 19, 'neigh_op_top_3')
// (17, 19, 'sp4_r_v_b_34')
// (17, 20, 'local_g3_3')
// (17, 20, 'lutff_3/in_1')
// (17, 20, 'lutff_3/out')
// (17, 20, 'lutff_6/in_2')
// (17, 20, 'sp4_h_r_6')
// (17, 20, 'sp4_r_v_b_23')
// (17, 20, 'sp4_r_v_b_39')
// (17, 21, 'local_g1_3')
// (17, 21, 'lutff_0/in_0')
// (17, 21, 'lutff_2/in_0')
// (17, 21, 'lutff_5/in_3')
// (17, 21, 'lutff_7/in_3')
// (17, 21, 'neigh_op_bot_3')
// (17, 21, 'sp4_r_v_b_10')
// (17, 21, 'sp4_r_v_b_26')
// (17, 22, 'sp4_r_v_b_15')
// (17, 23, 'sp4_r_v_b_2')
// (18, 17, 'sp4_v_t_47')
// (18, 18, 'sp4_v_b_47')
// (18, 19, 'neigh_op_tnl_3')
// (18, 19, 'sp4_h_r_7')
// (18, 19, 'sp4_v_b_34')
// (18, 19, 'sp4_v_t_39')
// (18, 20, 'neigh_op_lft_3')
// (18, 20, 'sp4_h_r_19')
// (18, 20, 'sp4_v_b_23')
// (18, 20, 'sp4_v_b_39')
// (18, 21, 'neigh_op_bnl_3')
// (18, 21, 'sp4_h_r_4')
// (18, 21, 'sp4_v_b_10')
// (18, 21, 'sp4_v_b_26')
// (18, 22, 'sp4_v_b_15')
// (18, 23, 'sp4_v_b_2')
// (19, 19, 'sp4_h_r_18')
// (19, 20, 'sp4_h_r_30')
// (19, 21, 'sp4_h_r_17')
// (20, 17, 'sp4_r_v_b_37')
// (20, 18, 'sp4_r_v_b_24')
// (20, 19, 'sp4_h_r_31')
// (20, 19, 'sp4_r_v_b_13')
// (20, 20, 'sp4_h_r_43')
// (20, 20, 'sp4_r_v_b_0')
// (20, 21, 'sp4_h_r_28')
// (21, 16, 'sp4_v_t_37')
// (21, 17, 'sp4_v_b_37')
// (21, 18, 'sp4_v_b_24')
// (21, 19, 'local_g0_5')
// (21, 19, 'lutff_3/in_0')
// (21, 19, 'sp4_h_r_42')
// (21, 19, 'sp4_v_b_13')
// (21, 20, 'sp4_h_l_43')
// (21, 20, 'sp4_v_b_0')
// (21, 21, 'local_g2_1')
// (21, 21, 'lutff_6/in_3')
// (21, 21, 'sp4_h_r_41')
// (22, 19, 'local_g1_7')
// (22, 19, 'lutff_5/in_3')
// (22, 19, 'lutff_7/in_1')
// (22, 19, 'sp4_h_l_42')
// (22, 19, 'sp4_h_r_7')
// (22, 21, 'sp4_h_l_41')
// (23, 19, 'sp4_h_r_18')
// (24, 19, 'sp4_h_r_31')
// (25, 19, 'sp4_h_r_42')

reg n2427 = 0;
// (16, 19, 'neigh_op_tnr_5')
// (16, 20, 'neigh_op_rgt_5')
// (16, 21, 'neigh_op_bnr_5')
// (17, 19, 'local_g1_5')
// (17, 19, 'lutff_0/in_2')
// (17, 19, 'neigh_op_top_5')
// (17, 20, 'local_g1_5')
// (17, 20, 'lutff_1/in_1')
// (17, 20, 'lutff_5/in_3')
// (17, 20, 'lutff_5/out')
// (17, 20, 'lutff_6/in_0')
// (17, 20, 'sp4_h_r_10')
// (17, 20, 'sp4_r_v_b_43')
// (17, 21, 'local_g0_5')
// (17, 21, 'lutff_0/in_1')
// (17, 21, 'lutff_1/in_2')
// (17, 21, 'lutff_5/in_2')
// (17, 21, 'lutff_7/in_0')
// (17, 21, 'neigh_op_bot_5')
// (17, 21, 'sp4_r_v_b_30')
// (17, 22, 'sp4_r_v_b_19')
// (17, 23, 'sp4_r_v_b_6')
// (18, 19, 'neigh_op_tnl_5')
// (18, 19, 'sp4_h_r_6')
// (18, 19, 'sp4_v_t_43')
// (18, 20, 'neigh_op_lft_5')
// (18, 20, 'sp4_h_r_23')
// (18, 20, 'sp4_v_b_43')
// (18, 21, 'neigh_op_bnl_5')
// (18, 21, 'sp4_v_b_30')
// (18, 22, 'sp4_v_b_19')
// (18, 23, 'sp4_v_b_6')
// (19, 19, 'sp4_h_r_19')
// (19, 20, 'sp4_h_r_34')
// (20, 17, 'sp4_r_v_b_41')
// (20, 18, 'sp4_r_v_b_28')
// (20, 19, 'sp4_h_r_30')
// (20, 19, 'sp4_r_v_b_17')
// (20, 20, 'sp4_h_r_47')
// (20, 20, 'sp4_r_v_b_4')
// (20, 21, 'sp4_r_v_b_38')
// (20, 22, 'sp4_r_v_b_27')
// (20, 23, 'sp4_r_v_b_14')
// (20, 24, 'sp4_r_v_b_3')
// (21, 16, 'sp4_v_t_41')
// (21, 17, 'sp4_v_b_41')
// (21, 18, 'sp4_v_b_28')
// (21, 19, 'local_g1_1')
// (21, 19, 'lutff_3/in_3')
// (21, 19, 'sp4_h_r_43')
// (21, 19, 'sp4_v_b_17')
// (21, 20, 'sp4_h_l_47')
// (21, 20, 'sp4_v_b_4')
// (21, 20, 'sp4_v_t_38')
// (21, 21, 'local_g2_6')
// (21, 21, 'lutff_6/in_0')
// (21, 21, 'sp4_v_b_38')
// (21, 22, 'sp4_v_b_27')
// (21, 23, 'sp4_v_b_14')
// (21, 24, 'sp4_v_b_3')
// (22, 19, 'local_g1_2')
// (22, 19, 'lutff_5/in_2')
// (22, 19, 'lutff_7/in_2')
// (22, 19, 'sp4_h_l_43')
// (22, 19, 'sp4_h_r_2')
// (23, 19, 'sp4_h_r_15')
// (24, 19, 'sp4_h_r_26')
// (25, 19, 'sp4_h_r_39')

wire n2428;
// (16, 20, 'local_g2_0')
// (16, 20, 'lutff_2/in_0')
// (16, 20, 'neigh_op_tnr_0')
// (16, 21, 'neigh_op_rgt_0')
// (16, 22, 'local_g1_0')
// (16, 22, 'lutff_2/in_1')
// (16, 22, 'neigh_op_bnr_0')
// (17, 18, 'sp4_r_v_b_36')
// (17, 19, 'sp4_r_v_b_25')
// (17, 19, 'sp4_r_v_b_41')
// (17, 20, 'neigh_op_top_0')
// (17, 20, 'sp4_r_v_b_12')
// (17, 20, 'sp4_r_v_b_28')
// (17, 21, 'local_g1_0')
// (17, 21, 'lutff_0/out')
// (17, 21, 'lutff_4/in_3')
// (17, 21, 'sp4_h_r_0')
// (17, 21, 'sp4_r_v_b_1')
// (17, 21, 'sp4_r_v_b_17')
// (17, 22, 'neigh_op_bot_0')
// (17, 22, 'sp4_r_v_b_4')
// (18, 17, 'sp4_h_r_6')
// (18, 17, 'sp4_v_t_36')
// (18, 18, 'sp4_h_r_4')
// (18, 18, 'sp4_v_b_36')
// (18, 18, 'sp4_v_t_41')
// (18, 19, 'sp4_v_b_25')
// (18, 19, 'sp4_v_b_41')
// (18, 20, 'neigh_op_tnl_0')
// (18, 20, 'sp4_v_b_12')
// (18, 20, 'sp4_v_b_28')
// (18, 21, 'local_g0_0')
// (18, 21, 'lutff_2/in_2')
// (18, 21, 'neigh_op_lft_0')
// (18, 21, 'sp4_h_r_13')
// (18, 21, 'sp4_v_b_1')
// (18, 21, 'sp4_v_b_17')
// (18, 22, 'neigh_op_bnl_0')
// (18, 22, 'sp4_h_r_10')
// (18, 22, 'sp4_v_b_4')
// (19, 17, 'sp4_h_r_19')
// (19, 18, 'sp4_h_r_17')
// (19, 21, 'sp4_h_r_24')
// (19, 22, 'sp4_h_r_23')
// (20, 17, 'sp4_h_r_30')
// (20, 18, 'local_g3_4')
// (20, 18, 'lutff_5/in_2')
// (20, 18, 'sp4_h_r_28')
// (20, 21, 'local_g3_5')
// (20, 21, 'lutff_6/in_2')
// (20, 21, 'sp4_h_r_37')
// (20, 22, 'sp4_h_r_34')
// (21, 14, 'sp4_r_v_b_37')
// (21, 15, 'sp4_r_v_b_24')
// (21, 16, 'local_g2_5')
// (21, 16, 'lutff_5/in_0')
// (21, 16, 'sp4_r_v_b_13')
// (21, 17, 'sp4_h_r_43')
// (21, 17, 'sp4_r_v_b_0')
// (21, 18, 'sp4_h_r_41')
// (21, 21, 'sp4_h_l_37')
// (21, 22, 'local_g3_7')
// (21, 22, 'lutff_5/in_3')
// (21, 22, 'sp4_h_r_47')
// (22, 13, 'sp4_v_t_37')
// (22, 14, 'sp4_v_b_37')
// (22, 15, 'sp4_v_b_24')
// (22, 16, 'sp4_v_b_13')
// (22, 17, 'sp4_h_l_43')
// (22, 17, 'sp4_v_b_0')
// (22, 18, 'sp4_h_l_41')
// (22, 22, 'sp4_h_l_47')

wire n2429;
// (16, 20, 'neigh_op_tnr_1')
// (16, 21, 'neigh_op_rgt_1')
// (16, 22, 'neigh_op_bnr_1')
// (17, 20, 'neigh_op_top_1')
// (17, 21, 'local_g2_1')
// (17, 21, 'lutff_1/out')
// (17, 21, 'lutff_2/in_3')
// (17, 22, 'neigh_op_bot_1')
// (18, 20, 'neigh_op_tnl_1')
// (18, 21, 'neigh_op_lft_1')
// (18, 22, 'neigh_op_bnl_1')

reg n2430 = 0;
// (16, 20, 'neigh_op_tnr_3')
// (16, 21, 'neigh_op_rgt_3')
// (16, 22, 'neigh_op_bnr_3')
// (17, 18, 'sp4_r_v_b_42')
// (17, 19, 'sp4_r_v_b_31')
// (17, 20, 'neigh_op_top_3')
// (17, 20, 'sp4_r_v_b_18')
// (17, 21, 'lutff_3/out')
// (17, 21, 'sp4_r_v_b_7')
// (17, 22, 'neigh_op_bot_3')
// (18, 17, 'sp4_v_t_42')
// (18, 18, 'sp4_v_b_42')
// (18, 19, 'local_g2_7')
// (18, 19, 'lutff_5/in_2')
// (18, 19, 'sp4_v_b_31')
// (18, 20, 'neigh_op_tnl_3')
// (18, 20, 'sp4_v_b_18')
// (18, 21, 'neigh_op_lft_3')
// (18, 21, 'sp4_v_b_7')
// (18, 22, 'neigh_op_bnl_3')

wire n2431;
// (16, 20, 'neigh_op_tnr_6')
// (16, 21, 'neigh_op_rgt_6')
// (16, 21, 'sp4_h_r_1')
// (16, 22, 'neigh_op_bnr_6')
// (17, 20, 'neigh_op_top_6')
// (17, 21, 'lutff_6/out')
// (17, 21, 'sp4_h_r_12')
// (17, 22, 'neigh_op_bot_6')
// (18, 20, 'neigh_op_tnl_6')
// (18, 21, 'neigh_op_lft_6')
// (18, 21, 'sp4_h_r_25')
// (18, 22, 'neigh_op_bnl_6')
// (19, 21, 'sp4_h_r_36')
// (20, 21, 'sp4_h_l_36')
// (20, 21, 'sp4_h_r_9')
// (21, 21, 'local_g1_4')
// (21, 21, 'lutff_2/in_1')
// (21, 21, 'sp4_h_r_20')
// (22, 21, 'sp4_h_r_33')
// (23, 21, 'sp4_h_r_44')
// (24, 21, 'sp4_h_l_44')

wire n2432;
// (16, 20, 'neigh_op_tnr_7')
// (16, 21, 'neigh_op_rgt_7')
// (16, 21, 'sp4_h_r_3')
// (16, 22, 'neigh_op_bnr_7')
// (17, 15, 'sp4_r_v_b_39')
// (17, 16, 'sp4_r_v_b_26')
// (17, 17, 'sp4_r_v_b_15')
// (17, 18, 'sp4_r_v_b_2')
// (17, 19, 'sp4_r_v_b_39')
// (17, 20, 'neigh_op_top_7')
// (17, 20, 'sp4_r_v_b_26')
// (17, 20, 'sp4_r_v_b_42')
// (17, 21, 'lutff_7/out')
// (17, 21, 'sp4_h_r_14')
// (17, 21, 'sp4_r_v_b_15')
// (17, 21, 'sp4_r_v_b_31')
// (17, 22, 'local_g0_7')
// (17, 22, 'lutff_6/in_1')
// (17, 22, 'neigh_op_bot_7')
// (17, 22, 'sp4_r_v_b_18')
// (17, 22, 'sp4_r_v_b_2')
// (17, 23, 'local_g1_7')
// (17, 23, 'lutff_2/in_2')
// (17, 23, 'sp4_r_v_b_7')
// (18, 14, 'sp4_v_t_39')
// (18, 15, 'local_g3_7')
// (18, 15, 'lutff_5/in_3')
// (18, 15, 'sp4_v_b_39')
// (18, 16, 'sp4_v_b_26')
// (18, 17, 'local_g0_7')
// (18, 17, 'lutff_3/in_0')
// (18, 17, 'sp4_v_b_15')
// (18, 18, 'local_g1_2')
// (18, 18, 'lutff_2/in_1')
// (18, 18, 'sp4_v_b_2')
// (18, 18, 'sp4_v_t_39')
// (18, 19, 'sp4_v_b_39')
// (18, 19, 'sp4_v_t_42')
// (18, 20, 'neigh_op_tnl_7')
// (18, 20, 'sp4_v_b_26')
// (18, 20, 'sp4_v_b_42')
// (18, 21, 'neigh_op_lft_7')
// (18, 21, 'sp4_h_r_27')
// (18, 21, 'sp4_v_b_15')
// (18, 21, 'sp4_v_b_31')
// (18, 22, 'neigh_op_bnl_7')
// (18, 22, 'sp4_v_b_18')
// (18, 22, 'sp4_v_b_2')
// (18, 23, 'sp4_v_b_7')
// (19, 14, 'sp4_r_v_b_37')
// (19, 15, 'sp4_r_v_b_24')
// (19, 16, 'sp4_r_v_b_13')
// (19, 17, 'sp4_r_v_b_0')
// (19, 18, 'sp4_r_v_b_44')
// (19, 19, 'sp4_r_v_b_33')
// (19, 20, 'sp4_r_v_b_20')
// (19, 21, 'sp4_h_r_38')
// (19, 21, 'sp4_r_v_b_9')
// (19, 22, 'sp4_r_v_b_45')
// (19, 23, 'sp4_r_v_b_32')
// (19, 24, 'sp4_r_v_b_21')
// (19, 25, 'sp4_r_v_b_8')
// (20, 13, 'sp4_v_t_37')
// (20, 14, 'sp4_v_b_37')
// (20, 15, 'local_g2_0')
// (20, 15, 'lutff_5/in_1')
// (20, 15, 'sp4_v_b_24')
// (20, 16, 'sp4_v_b_13')
// (20, 17, 'sp4_v_b_0')
// (20, 17, 'sp4_v_t_44')
// (20, 18, 'sp4_v_b_44')
// (20, 19, 'sp4_v_b_33')
// (20, 20, 'local_g1_4')
// (20, 20, 'lutff_4/in_3')
// (20, 20, 'sp4_v_b_20')
// (20, 21, 'sp4_h_l_38')
// (20, 21, 'sp4_v_b_9')
// (20, 21, 'sp4_v_t_45')
// (20, 22, 'sp4_v_b_45')
// (20, 23, 'local_g3_0')
// (20, 23, 'lutff_3/in_0')
// (20, 23, 'sp4_v_b_32')
// (20, 24, 'sp4_v_b_21')
// (20, 25, 'sp4_v_b_8')

reg n2433 = 0;
// (16, 21, 'neigh_op_tnr_1')
// (16, 22, 'neigh_op_rgt_1')
// (16, 23, 'neigh_op_bnr_1')
// (17, 21, 'local_g0_1')
// (17, 21, 'lutff_6/in_1')
// (17, 21, 'neigh_op_top_1')
// (17, 22, 'lutff_1/out')
// (17, 23, 'neigh_op_bot_1')
// (18, 21, 'neigh_op_tnl_1')
// (18, 22, 'neigh_op_lft_1')
// (18, 23, 'neigh_op_bnl_1')

wire n2434;
// (16, 21, 'neigh_op_tnr_5')
// (16, 22, 'neigh_op_rgt_5')
// (16, 23, 'neigh_op_bnr_5')
// (17, 21, 'neigh_op_top_5')
// (17, 21, 'sp4_r_v_b_38')
// (17, 22, 'lutff_5/out')
// (17, 22, 'sp4_r_v_b_27')
// (17, 23, 'neigh_op_bot_5')
// (17, 23, 'sp4_r_v_b_14')
// (17, 24, 'sp4_r_v_b_3')
// (18, 20, 'sp4_h_r_8')
// (18, 20, 'sp4_v_t_38')
// (18, 21, 'neigh_op_tnl_5')
// (18, 21, 'sp4_v_b_38')
// (18, 22, 'neigh_op_lft_5')
// (18, 22, 'sp4_v_b_27')
// (18, 23, 'neigh_op_bnl_5')
// (18, 23, 'sp4_v_b_14')
// (18, 24, 'sp4_v_b_3')
// (19, 20, 'sp4_h_r_21')
// (20, 20, 'local_g3_0')
// (20, 20, 'lutff_7/in_0')
// (20, 20, 'sp4_h_r_32')
// (21, 20, 'sp4_h_r_45')
// (22, 20, 'sp4_h_l_45')

reg n2435 = 0;
// (16, 21, 'sp4_r_v_b_41')
// (16, 22, 'sp4_r_v_b_28')
// (16, 23, 'neigh_op_tnr_2')
// (16, 23, 'sp4_r_v_b_17')
// (16, 24, 'neigh_op_rgt_2')
// (16, 24, 'sp4_r_v_b_4')
// (16, 25, 'neigh_op_bnr_2')
// (17, 20, 'sp4_v_t_41')
// (17, 21, 'local_g3_1')
// (17, 21, 'lutff_6/in_2')
// (17, 21, 'sp4_v_b_41')
// (17, 22, 'sp4_v_b_28')
// (17, 23, 'neigh_op_top_2')
// (17, 23, 'sp4_v_b_17')
// (17, 24, 'lutff_2/out')
// (17, 24, 'sp4_v_b_4')
// (17, 25, 'neigh_op_bot_2')
// (18, 23, 'neigh_op_tnl_2')
// (18, 24, 'neigh_op_lft_2')
// (18, 25, 'neigh_op_bnl_2')

reg n2436 = 0;
// (16, 22, 'neigh_op_tnr_1')
// (16, 23, 'neigh_op_rgt_1')
// (16, 23, 'sp4_h_r_7')
// (16, 24, 'neigh_op_bnr_1')
// (17, 22, 'neigh_op_top_1')
// (17, 23, 'lutff_1/out')
// (17, 23, 'sp4_h_r_18')
// (17, 24, 'neigh_op_bot_1')
// (18, 22, 'neigh_op_tnl_1')
// (18, 23, 'neigh_op_lft_1')
// (18, 23, 'sp4_h_r_31')
// (18, 24, 'neigh_op_bnl_1')
// (19, 20, 'sp4_r_v_b_36')
// (19, 21, 'sp4_r_v_b_25')
// (19, 22, 'sp4_r_v_b_12')
// (19, 23, 'sp4_h_r_42')
// (19, 23, 'sp4_r_v_b_1')
// (20, 19, 'sp4_v_t_36')
// (20, 20, 'sp4_v_b_36')
// (20, 21, 'sp4_v_b_25')
// (20, 22, 'local_g1_4')
// (20, 22, 'lutff_5/in_2')
// (20, 22, 'sp4_v_b_12')
// (20, 23, 'sp4_h_l_42')
// (20, 23, 'sp4_v_b_1')

wire n2437;
// (16, 22, 'neigh_op_tnr_2')
// (16, 23, 'neigh_op_rgt_2')
// (16, 24, 'neigh_op_bnr_2')
// (17, 22, 'neigh_op_top_2')
// (17, 23, 'local_g2_2')
// (17, 23, 'lutff_2/out')
// (17, 23, 'lutff_global/cen')
// (17, 24, 'neigh_op_bot_2')
// (18, 22, 'neigh_op_tnl_2')
// (18, 23, 'neigh_op_lft_2')
// (18, 24, 'neigh_op_bnl_2')

wire n2438;
// (16, 23, 'neigh_op_tnr_7')
// (16, 24, 'neigh_op_rgt_7')
// (16, 24, 'sp4_h_r_3')
// (16, 24, 'sp4_h_r_6')
// (16, 25, 'neigh_op_bnr_7')
// (17, 23, 'neigh_op_top_7')
// (17, 24, 'local_g1_3')
// (17, 24, 'lutff_7/out')
// (17, 24, 'lutff_global/cen')
// (17, 24, 'sp4_h_r_14')
// (17, 24, 'sp4_h_r_19')
// (17, 25, 'neigh_op_bot_7')
// (18, 23, 'neigh_op_tnl_7')
// (18, 24, 'neigh_op_lft_7')
// (18, 24, 'sp4_h_r_27')
// (18, 24, 'sp4_h_r_30')
// (18, 25, 'neigh_op_bnl_7')
// (19, 24, 'sp4_h_r_38')
// (19, 24, 'sp4_h_r_43')
// (20, 24, 'sp4_h_l_38')
// (20, 24, 'sp4_h_l_43')
// (20, 24, 'sp4_h_r_6')
// (21, 24, 'sp4_h_r_19')
// (22, 24, 'sp4_h_r_30')
// (23, 24, 'sp4_h_r_43')
// (24, 24, 'sp4_h_l_43')

wire n2439;
// (17, 0, 'logic_op_tnr_1')
// (17, 1, 'local_g2_1')
// (17, 1, 'lutff_1/in_0')
// (17, 1, 'lutff_2/in_3')
// (17, 1, 'lutff_3/in_0')
// (17, 1, 'neigh_op_rgt_1')
// (17, 2, 'neigh_op_bnr_1')
// (18, 0, 'logic_op_top_1')
// (18, 1, 'local_g3_1')
// (18, 1, 'lutff_1/out')
// (18, 1, 'lutff_5/in_1')
// (18, 2, 'neigh_op_bot_1')
// (19, 0, 'logic_op_tnl_1')
// (19, 1, 'neigh_op_lft_1')
// (19, 2, 'neigh_op_bnl_1')

wire n2440;
// (17, 0, 'logic_op_tnr_2')
// (17, 1, 'neigh_op_rgt_2')
// (17, 2, 'neigh_op_bnr_2')
// (18, 0, 'logic_op_top_2')
// (18, 1, 'lutff_2/out')
// (18, 2, 'local_g1_2')
// (18, 2, 'lutff_2/in_3')
// (18, 2, 'lutff_7/in_2')
// (18, 2, 'neigh_op_bot_2')
// (19, 0, 'logic_op_tnl_2')
// (19, 1, 'neigh_op_lft_2')
// (19, 2, 'neigh_op_bnl_2')

wire n2441;
// (17, 0, 'logic_op_tnr_3')
// (17, 1, 'neigh_op_rgt_3')
// (17, 2, 'neigh_op_bnr_3')
// (18, 0, 'logic_op_top_3')
// (18, 1, 'lutff_3/out')
// (18, 2, 'local_g0_3')
// (18, 2, 'lutff_2/in_1')
// (18, 2, 'lutff_7/in_0')
// (18, 2, 'neigh_op_bot_3')
// (19, 0, 'logic_op_tnl_3')
// (19, 1, 'neigh_op_lft_3')
// (19, 2, 'neigh_op_bnl_3')

wire n2442;
// (17, 0, 'logic_op_tnr_4')
// (17, 1, 'local_g2_4')
// (17, 1, 'lutff_1/in_1')
// (17, 1, 'lutff_2/in_0')
// (17, 1, 'lutff_3/in_3')
// (17, 1, 'neigh_op_rgt_4')
// (17, 2, 'neigh_op_bnr_4')
// (18, 0, 'logic_op_top_4')
// (18, 1, 'lutff_4/out')
// (18, 2, 'neigh_op_bot_4')
// (19, 0, 'logic_op_tnl_4')
// (19, 1, 'neigh_op_lft_4')
// (19, 2, 'neigh_op_bnl_4')

reg n2443 = 0;
// (17, 1, 'neigh_op_tnr_0')
// (17, 2, 'neigh_op_rgt_0')
// (17, 3, 'neigh_op_bnr_0')
// (18, 1, 'neigh_op_top_0')
// (18, 1, 'sp4_r_v_b_28')
// (18, 2, 'lutff_0/out')
// (18, 2, 'sp4_r_v_b_17')
// (18, 3, 'neigh_op_bot_0')
// (18, 3, 'sp4_r_v_b_4')
// (18, 4, 'sp4_r_v_b_42')
// (18, 5, 'sp4_r_v_b_31')
// (18, 6, 'sp4_r_v_b_18')
// (18, 7, 'sp4_r_v_b_7')
// (19, 0, 'span4_vert_28')
// (19, 1, 'neigh_op_tnl_0')
// (19, 1, 'sp4_v_b_28')
// (19, 2, 'neigh_op_lft_0')
// (19, 2, 'sp4_v_b_17')
// (19, 3, 'neigh_op_bnl_0')
// (19, 3, 'sp4_v_b_4')
// (19, 3, 'sp4_v_t_42')
// (19, 4, 'sp4_v_b_42')
// (19, 5, 'local_g3_7')
// (19, 5, 'ram/WDATA_8')
// (19, 5, 'sp4_v_b_31')
// (19, 6, 'sp4_v_b_18')
// (19, 7, 'sp4_v_b_7')

reg n2444 = 0;
// (17, 1, 'neigh_op_tnr_1')
// (17, 2, 'neigh_op_rgt_1')
// (17, 3, 'neigh_op_bnr_1')
// (18, 1, 'neigh_op_top_1')
// (18, 1, 'sp4_r_v_b_46')
// (18, 2, 'lutff_1/out')
// (18, 2, 'sp4_r_v_b_35')
// (18, 3, 'neigh_op_bot_1')
// (18, 3, 'sp4_r_v_b_22')
// (18, 4, 'sp4_r_v_b_11')
// (18, 5, 'sp4_r_v_b_42')
// (18, 6, 'sp4_r_v_b_31')
// (18, 7, 'sp4_r_v_b_18')
// (18, 8, 'sp4_r_v_b_7')
// (19, 0, 'span4_vert_46')
// (19, 1, 'neigh_op_tnl_1')
// (19, 1, 'sp4_v_b_46')
// (19, 2, 'neigh_op_lft_1')
// (19, 2, 'sp4_v_b_35')
// (19, 3, 'neigh_op_bnl_1')
// (19, 3, 'sp4_v_b_22')
// (19, 4, 'sp4_v_b_11')
// (19, 4, 'sp4_v_t_42')
// (19, 5, 'sp4_v_b_42')
// (19, 6, 'local_g3_7')
// (19, 6, 'ram/WDATA_6')
// (19, 6, 'sp4_v_b_31')
// (19, 7, 'sp4_v_b_18')
// (19, 8, 'sp4_v_b_7')

reg n2445 = 0;
// (17, 1, 'neigh_op_tnr_3')
// (17, 2, 'neigh_op_rgt_3')
// (17, 3, 'neigh_op_bnr_3')
// (18, 1, 'neigh_op_top_3')
// (18, 1, 'sp4_r_v_b_34')
// (18, 2, 'lutff_3/out')
// (18, 2, 'sp4_r_v_b_23')
// (18, 3, 'neigh_op_bot_3')
// (18, 3, 'sp4_r_v_b_10')
// (18, 4, 'sp4_r_v_b_47')
// (18, 5, 'sp4_r_v_b_34')
// (18, 6, 'sp4_r_v_b_23')
// (18, 7, 'sp4_r_v_b_10')
// (19, 0, 'span4_vert_34')
// (19, 1, 'neigh_op_tnl_3')
// (19, 1, 'sp4_v_b_34')
// (19, 2, 'neigh_op_lft_3')
// (19, 2, 'sp4_v_b_23')
// (19, 3, 'neigh_op_bnl_3')
// (19, 3, 'sp4_v_b_10')
// (19, 3, 'sp4_v_t_47')
// (19, 4, 'sp4_v_b_47')
// (19, 5, 'sp4_v_b_34')
// (19, 6, 'local_g0_7')
// (19, 6, 'ram/WDATA_1')
// (19, 6, 'sp4_v_b_23')
// (19, 7, 'sp4_v_b_10')

reg n2446 = 0;
// (17, 1, 'neigh_op_tnr_5')
// (17, 2, 'neigh_op_rgt_5')
// (17, 3, 'neigh_op_bnr_5')
// (18, 1, 'neigh_op_top_5')
// (18, 1, 'sp4_r_v_b_22')
// (18, 2, 'lutff_5/out')
// (18, 2, 'sp4_r_v_b_11')
// (18, 3, 'neigh_op_bot_5')
// (18, 3, 'sp4_r_v_b_42')
// (18, 4, 'sp4_r_v_b_31')
// (18, 5, 'sp4_r_v_b_18')
// (18, 6, 'sp4_r_v_b_7')
// (19, 0, 'span4_vert_22')
// (19, 1, 'neigh_op_tnl_5')
// (19, 1, 'sp4_v_b_22')
// (19, 2, 'neigh_op_lft_5')
// (19, 2, 'sp4_v_b_11')
// (19, 2, 'sp4_v_t_42')
// (19, 3, 'neigh_op_bnl_5')
// (19, 3, 'sp4_v_b_42')
// (19, 4, 'sp4_v_b_31')
// (19, 5, 'sp4_v_b_18')
// (19, 6, 'local_g1_7')
// (19, 6, 'ram/WDATA_2')
// (19, 6, 'sp4_v_b_7')

reg n2447 = 0;
// (17, 1, 'sp4_h_r_1')
// (18, 1, 'local_g0_4')
// (18, 1, 'lutff_2/in_2')
// (18, 1, 'sp4_h_r_12')
// (19, 0, 'logic_op_tnr_2')
// (19, 1, 'neigh_op_rgt_2')
// (19, 1, 'sp4_h_r_25')
// (19, 2, 'neigh_op_bnr_2')
// (20, 0, 'logic_op_top_2')
// (20, 1, 'local_g1_2')
// (20, 1, 'lutff_2/in_1')
// (20, 1, 'lutff_2/out')
// (20, 1, 'sp4_h_r_36')
// (20, 2, 'neigh_op_bot_2')
// (21, 0, 'logic_op_tnl_2')
// (21, 1, 'local_g1_2')
// (21, 1, 'lutff_0/in_1')
// (21, 1, 'lutff_5/in_0')
// (21, 1, 'neigh_op_lft_2')
// (21, 1, 'sp4_h_l_36')
// (21, 2, 'neigh_op_bnl_2')

reg n2448 = 0;
// (17, 1, 'sp4_h_r_3')
// (18, 1, 'local_g0_6')
// (18, 1, 'lutff_3/in_1')
// (18, 1, 'sp4_h_r_14')
// (19, 0, 'logic_op_tnr_3')
// (19, 1, 'neigh_op_rgt_3')
// (19, 1, 'sp4_h_r_27')
// (19, 2, 'neigh_op_bnr_3')
// (20, 0, 'logic_op_top_3')
// (20, 1, 'local_g2_3')
// (20, 1, 'lutff_3/in_0')
// (20, 1, 'lutff_3/out')
// (20, 1, 'sp4_h_r_38')
// (20, 2, 'neigh_op_bot_3')
// (21, 0, 'logic_op_tnl_3')
// (21, 1, 'local_g1_3')
// (21, 1, 'lutff_0/in_2')
// (21, 1, 'lutff_5/in_3')
// (21, 1, 'neigh_op_lft_3')
// (21, 1, 'sp4_h_l_38')
// (21, 2, 'neigh_op_bnl_3')

wire n2449;
// (17, 2, 'sp4_h_r_5')
// (17, 4, 'local_g0_6')
// (17, 4, 'lutff_4/in_0')
// (17, 4, 'sp4_h_r_6')
// (18, 2, 'local_g0_0')
// (18, 2, 'lutff_1/in_1')
// (18, 2, 'sp4_h_r_16')
// (18, 4, 'sp4_h_r_19')
// (19, 1, 'neigh_op_tnr_4')
// (19, 2, 'neigh_op_rgt_4')
// (19, 2, 'sp4_h_r_29')
// (19, 3, 'neigh_op_bnr_4')
// (19, 4, 'sp4_h_r_30')
// (20, 1, 'neigh_op_top_4')
// (20, 1, 'sp4_r_v_b_36')
// (20, 2, 'local_g1_4')
// (20, 2, 'lutff_0/in_1')
// (20, 2, 'lutff_4/out')
// (20, 2, 'sp4_h_r_40')
// (20, 2, 'sp4_r_v_b_25')
// (20, 3, 'neigh_op_bot_4')
// (20, 3, 'sp4_r_v_b_12')
// (20, 4, 'sp4_h_r_43')
// (20, 4, 'sp4_r_v_b_1')
// (21, 0, 'span4_vert_36')
// (21, 1, 'neigh_op_tnl_4')
// (21, 1, 'sp4_v_b_36')
// (21, 2, 'neigh_op_lft_4')
// (21, 2, 'sp4_h_l_40')
// (21, 2, 'sp4_v_b_25')
// (21, 3, 'neigh_op_bnl_4')
// (21, 3, 'sp4_v_b_12')
// (21, 4, 'sp4_h_l_43')
// (21, 4, 'sp4_v_b_1')

reg n2450 = 0;
// (17, 3, 'neigh_op_tnr_0')
// (17, 4, 'neigh_op_rgt_0')
// (17, 5, 'neigh_op_bnr_0')
// (18, 3, 'neigh_op_top_0')
// (18, 4, 'lutff_0/out')
// (18, 5, 'local_g0_0')
// (18, 5, 'lutff_0/in_0')
// (18, 5, 'lutff_6/in_0')
// (18, 5, 'neigh_op_bot_0')
// (19, 3, 'neigh_op_tnl_0')
// (19, 4, 'neigh_op_lft_0')
// (19, 5, 'neigh_op_bnl_0')

reg n2451 = 0;
// (17, 3, 'neigh_op_tnr_1')
// (17, 4, 'neigh_op_rgt_1')
// (17, 5, 'neigh_op_bnr_1')
// (18, 3, 'neigh_op_top_1')
// (18, 4, 'lutff_1/out')
// (18, 5, 'local_g1_1')
// (18, 5, 'lutff_0/in_2')
// (18, 5, 'lutff_4/in_2')
// (18, 5, 'neigh_op_bot_1')
// (19, 3, 'neigh_op_tnl_1')
// (19, 4, 'neigh_op_lft_1')
// (19, 5, 'neigh_op_bnl_1')

reg n2452 = 0;
// (17, 3, 'neigh_op_tnr_2')
// (17, 4, 'neigh_op_rgt_2')
// (17, 5, 'neigh_op_bnr_2')
// (18, 3, 'neigh_op_top_2')
// (18, 4, 'lutff_2/out')
// (18, 5, 'local_g1_2')
// (18, 5, 'lutff_0/in_3')
// (18, 5, 'lutff_5/in_2')
// (18, 5, 'neigh_op_bot_2')
// (19, 3, 'neigh_op_tnl_2')
// (19, 4, 'neigh_op_lft_2')
// (19, 5, 'neigh_op_bnl_2')

reg n2453 = 0;
// (17, 3, 'neigh_op_tnr_3')
// (17, 4, 'neigh_op_rgt_3')
// (17, 5, 'neigh_op_bnr_3')
// (18, 3, 'neigh_op_top_3')
// (18, 4, 'lutff_3/out')
// (18, 5, 'local_g0_3')
// (18, 5, 'lutff_0/in_1')
// (18, 5, 'lutff_2/in_1')
// (18, 5, 'neigh_op_bot_3')
// (19, 3, 'neigh_op_tnl_3')
// (19, 4, 'neigh_op_lft_3')
// (19, 5, 'neigh_op_bnl_3')

reg n2454 = 0;
// (17, 3, 'sp4_r_v_b_39')
// (17, 4, 'sp4_r_v_b_26')
// (17, 5, 'sp4_r_v_b_15')
// (17, 6, 'sp4_r_v_b_2')
// (18, 2, 'sp4_v_t_39')
// (18, 3, 'local_g2_7')
// (18, 3, 'lutff_7/in_2')
// (18, 3, 'sp4_v_b_39')
// (18, 4, 'sp4_v_b_26')
// (18, 5, 'sp4_v_b_15')
// (18, 6, 'sp4_h_r_9')
// (18, 6, 'sp4_v_b_2')
// (19, 6, 'sp4_h_r_20')
// (20, 1, 'sp4_r_v_b_28')
// (20, 2, 'sp4_r_v_b_17')
// (20, 3, 'local_g1_4')
// (20, 3, 'lutff_1/in_0')
// (20, 3, 'sp4_r_v_b_4')
// (20, 4, 'sp4_r_v_b_36')
// (20, 5, 'neigh_op_tnr_6')
// (20, 5, 'sp4_r_v_b_25')
// (20, 6, 'neigh_op_rgt_6')
// (20, 6, 'sp4_h_r_33')
// (20, 6, 'sp4_r_v_b_12')
// (20, 7, 'neigh_op_bnr_6')
// (20, 7, 'sp4_r_v_b_1')
// (21, 0, 'span4_vert_28')
// (21, 1, 'sp4_v_b_28')
// (21, 2, 'sp4_v_b_17')
// (21, 3, 'sp4_v_b_4')
// (21, 3, 'sp4_v_t_36')
// (21, 4, 'sp4_v_b_36')
// (21, 5, 'neigh_op_top_6')
// (21, 5, 'sp4_v_b_25')
// (21, 6, 'lutff_6/out')
// (21, 6, 'sp4_h_r_44')
// (21, 6, 'sp4_v_b_12')
// (21, 7, 'neigh_op_bot_6')
// (21, 7, 'sp4_v_b_1')
// (22, 5, 'neigh_op_tnl_6')
// (22, 6, 'neigh_op_lft_6')
// (22, 6, 'sp4_h_l_44')
// (22, 7, 'neigh_op_bnl_6')

reg n2455 = 0;
// (17, 3, 'sp4_r_v_b_40')
// (17, 4, 'sp4_r_v_b_29')
// (17, 5, 'sp4_r_v_b_16')
// (17, 6, 'sp4_r_v_b_5')
// (18, 2, 'sp4_v_t_40')
// (18, 3, 'local_g2_0')
// (18, 3, 'lutff_2/in_2')
// (18, 3, 'sp4_v_b_40')
// (18, 4, 'sp4_v_b_29')
// (18, 5, 'sp4_v_b_16')
// (18, 6, 'sp4_h_r_5')
// (18, 6, 'sp4_v_b_5')
// (19, 6, 'sp4_h_r_16')
// (20, 5, 'neigh_op_tnr_4')
// (20, 6, 'neigh_op_rgt_4')
// (20, 6, 'sp4_h_r_29')
// (20, 7, 'neigh_op_bnr_4')
// (21, 5, 'neigh_op_top_4')
// (21, 6, 'lutff_4/out')
// (21, 6, 'sp4_h_r_40')
// (21, 7, 'neigh_op_bot_4')
// (22, 5, 'neigh_op_tnl_4')
// (22, 6, 'local_g1_4')
// (22, 6, 'lutff_1/in_0')
// (22, 6, 'neigh_op_lft_4')
// (22, 6, 'sp4_h_l_40')
// (22, 7, 'neigh_op_bnl_4')

wire n2456;
// (17, 3, 'sp4_r_v_b_43')
// (17, 4, 'sp4_r_v_b_30')
// (17, 5, 'local_g3_3')
// (17, 5, 'lutff_global/cen')
// (17, 5, 'sp4_r_v_b_19')
// (17, 6, 'sp4_r_v_b_6')
// (18, 2, 'local_g0_2')
// (18, 2, 'lutff_global/cen')
// (18, 2, 'sp4_h_r_10')
// (18, 2, 'sp4_v_t_43')
// (18, 3, 'sp4_v_b_43')
// (18, 4, 'sp4_v_b_30')
// (18, 5, 'local_g0_2')
// (18, 5, 'lutff_global/cen')
// (18, 5, 'sp4_h_r_10')
// (18, 5, 'sp4_v_b_19')
// (18, 6, 'sp4_h_r_1')
// (18, 6, 'sp4_v_b_6')
// (19, 2, 'sp4_h_r_23')
// (19, 5, 'sp4_h_r_23')
// (19, 6, 'sp4_h_r_12')
// (20, 2, 'sp4_h_r_34')
// (20, 5, 'sp4_h_r_34')
// (20, 6, 'sp4_h_r_25')
// (21, 2, 'sp4_h_r_47')
// (21, 2, 'sp4_r_v_b_38')
// (21, 3, 'sp4_r_v_b_27')
// (21, 3, 'sp4_r_v_b_47')
// (21, 4, 'sp4_r_v_b_14')
// (21, 4, 'sp4_r_v_b_34')
// (21, 5, 'neigh_op_tnr_5')
// (21, 5, 'sp4_h_r_47')
// (21, 5, 'sp4_r_v_b_23')
// (21, 5, 'sp4_r_v_b_3')
// (21, 6, 'neigh_op_rgt_5')
// (21, 6, 'sp4_h_r_36')
// (21, 6, 'sp4_r_v_b_10')
// (21, 6, 'sp4_r_v_b_42')
// (21, 7, 'neigh_op_bnr_5')
// (21, 7, 'sp4_r_v_b_31')
// (21, 8, 'sp4_r_v_b_18')
// (21, 9, 'sp4_r_v_b_7')
// (22, 1, 'sp4_v_t_38')
// (22, 2, 'sp4_h_l_47')
// (22, 2, 'sp4_v_b_38')
// (22, 2, 'sp4_v_t_47')
// (22, 3, 'sp4_v_b_27')
// (22, 3, 'sp4_v_b_47')
// (22, 4, 'sp4_v_b_14')
// (22, 4, 'sp4_v_b_34')
// (22, 5, 'local_g1_3')
// (22, 5, 'lutff_global/cen')
// (22, 5, 'neigh_op_top_5')
// (22, 5, 'sp4_h_l_47')
// (22, 5, 'sp4_h_r_7')
// (22, 5, 'sp4_v_b_23')
// (22, 5, 'sp4_v_b_3')
// (22, 5, 'sp4_v_t_42')
// (22, 6, 'lutff_5/out')
// (22, 6, 'sp4_h_l_36')
// (22, 6, 'sp4_h_r_10')
// (22, 6, 'sp4_v_b_10')
// (22, 6, 'sp4_v_b_42')
// (22, 7, 'neigh_op_bot_5')
// (22, 7, 'sp4_v_b_31')
// (22, 8, 'sp4_v_b_18')
// (22, 9, 'sp4_v_b_7')
// (23, 5, 'neigh_op_tnl_5')
// (23, 5, 'sp4_h_r_18')
// (23, 6, 'neigh_op_lft_5')
// (23, 6, 'sp4_h_r_23')
// (23, 7, 'neigh_op_bnl_5')
// (24, 5, 'sp4_h_r_31')
// (24, 6, 'sp4_h_r_34')
// (25, 5, 'sp4_h_r_42')
// (25, 6, 'sp4_h_r_47')

wire n2457;
// (17, 4, 'neigh_op_tnr_0')
// (17, 5, 'neigh_op_rgt_0')
// (17, 6, 'neigh_op_bnr_0')
// (18, 4, 'neigh_op_top_0')
// (18, 5, 'lutff_0/out')
// (18, 5, 'sp4_h_r_0')
// (18, 6, 'neigh_op_bot_0')
// (19, 4, 'neigh_op_tnl_0')
// (19, 5, 'neigh_op_lft_0')
// (19, 5, 'sp4_h_r_13')
// (19, 6, 'neigh_op_bnl_0')
// (20, 5, 'sp4_h_r_24')
// (21, 5, 'sp4_h_r_37')
// (22, 5, 'local_g0_0')
// (22, 5, 'lutff_6/in_2')
// (22, 5, 'sp4_h_l_37')
// (22, 5, 'sp4_h_r_0')
// (23, 5, 'local_g0_5')
// (23, 5, 'lutff_6/in_3')
// (23, 5, 'sp4_h_r_13')
// (24, 5, 'sp4_h_r_24')
// (25, 5, 'sp4_h_r_37')

reg n2458 = 0;
// (17, 4, 'neigh_op_tnr_1')
// (17, 5, 'neigh_op_rgt_1')
// (17, 6, 'neigh_op_bnr_1')
// (18, 4, 'neigh_op_top_1')
// (18, 5, 'lutff_1/out')
// (18, 6, 'neigh_op_bot_1')
// (19, 4, 'neigh_op_tnl_1')
// (19, 5, 'local_g0_1')
// (19, 5, 'neigh_op_lft_1')
// (19, 5, 'ram/WDATA_9')
// (19, 6, 'neigh_op_bnl_1')

reg n2459 = 0;
// (17, 4, 'neigh_op_tnr_2')
// (17, 5, 'neigh_op_rgt_2')
// (17, 6, 'neigh_op_bnr_2')
// (18, 4, 'neigh_op_top_2')
// (18, 5, 'lutff_2/out')
// (18, 5, 'sp4_r_v_b_37')
// (18, 6, 'neigh_op_bot_2')
// (18, 6, 'sp4_r_v_b_24')
// (18, 7, 'sp4_r_v_b_13')
// (18, 8, 'sp4_r_v_b_0')
// (19, 4, 'neigh_op_tnl_2')
// (19, 4, 'sp4_v_t_37')
// (19, 5, 'neigh_op_lft_2')
// (19, 5, 'sp4_v_b_37')
// (19, 6, 'neigh_op_bnl_2')
// (19, 6, 'sp4_v_b_24')
// (19, 7, 'sp4_v_b_13')
// (19, 8, 'local_g0_0')
// (19, 8, 'ram/WDATA_0')
// (19, 8, 'sp4_v_b_0')

reg n2460 = 0;
// (17, 4, 'neigh_op_tnr_3')
// (17, 5, 'neigh_op_rgt_3')
// (17, 6, 'neigh_op_bnr_3')
// (18, 4, 'neigh_op_top_3')
// (18, 5, 'lutff_3/out')
// (18, 6, 'neigh_op_bot_3')
// (19, 4, 'neigh_op_tnl_3')
// (19, 5, 'neigh_op_lft_3')
// (19, 6, 'local_g3_3')
// (19, 6, 'neigh_op_bnl_3')
// (19, 6, 'ram/WDATA_4')

reg n2461 = 0;
// (17, 4, 'neigh_op_tnr_4')
// (17, 5, 'neigh_op_rgt_4')
// (17, 6, 'neigh_op_bnr_4')
// (18, 4, 'neigh_op_top_4')
// (18, 5, 'lutff_4/out')
// (18, 5, 'sp4_r_v_b_41')
// (18, 6, 'neigh_op_bot_4')
// (18, 6, 'sp4_r_v_b_28')
// (18, 7, 'sp4_r_v_b_17')
// (18, 8, 'sp4_r_v_b_4')
// (19, 4, 'neigh_op_tnl_4')
// (19, 4, 'sp4_v_t_41')
// (19, 5, 'neigh_op_lft_4')
// (19, 5, 'sp4_v_b_41')
// (19, 6, 'neigh_op_bnl_4')
// (19, 6, 'sp4_v_b_28')
// (19, 7, 'sp4_v_b_17')
// (19, 8, 'local_g1_4')
// (19, 8, 'ram/WDATA_1')
// (19, 8, 'sp4_v_b_4')

reg n2462 = 0;
// (17, 4, 'neigh_op_tnr_5')
// (17, 5, 'neigh_op_rgt_5')
// (17, 6, 'neigh_op_bnr_5')
// (18, 4, 'neigh_op_top_5')
// (18, 5, 'lutff_5/out')
// (18, 5, 'sp4_r_v_b_43')
// (18, 6, 'neigh_op_bot_5')
// (18, 6, 'sp4_r_v_b_30')
// (18, 7, 'sp4_r_v_b_19')
// (18, 8, 'sp4_r_v_b_6')
// (19, 4, 'neigh_op_tnl_5')
// (19, 4, 'sp4_v_t_43')
// (19, 5, 'neigh_op_lft_5')
// (19, 5, 'sp4_v_b_43')
// (19, 6, 'neigh_op_bnl_5')
// (19, 6, 'sp4_v_b_30')
// (19, 7, 'sp4_v_b_19')
// (19, 8, 'local_g0_6')
// (19, 8, 'ram/WDATA_2')
// (19, 8, 'sp4_v_b_6')

reg n2463 = 0;
// (17, 4, 'neigh_op_tnr_6')
// (17, 5, 'neigh_op_rgt_6')
// (17, 6, 'neigh_op_bnr_6')
// (18, 4, 'neigh_op_top_6')
// (18, 5, 'lutff_6/out')
// (18, 5, 'sp4_r_v_b_45')
// (18, 6, 'neigh_op_bot_6')
// (18, 6, 'sp4_r_v_b_32')
// (18, 7, 'sp4_r_v_b_21')
// (18, 8, 'sp4_r_v_b_8')
// (19, 4, 'neigh_op_tnl_6')
// (19, 4, 'sp4_v_t_45')
// (19, 5, 'neigh_op_lft_6')
// (19, 5, 'sp4_v_b_45')
// (19, 6, 'neigh_op_bnl_6')
// (19, 6, 'sp4_v_b_32')
// (19, 7, 'sp4_v_b_21')
// (19, 8, 'local_g1_0')
// (19, 8, 'ram/WDATA_3')
// (19, 8, 'sp4_v_b_8')

reg n2464 = 0;
// (17, 4, 'neigh_op_tnr_7')
// (17, 5, 'neigh_op_rgt_7')
// (17, 6, 'neigh_op_bnr_7')
// (18, 4, 'neigh_op_top_7')
// (18, 5, 'lutff_7/out')
// (18, 6, 'neigh_op_bot_7')
// (19, 4, 'neigh_op_tnl_7')
// (19, 5, 'neigh_op_lft_7')
// (19, 6, 'local_g2_7')
// (19, 6, 'neigh_op_bnl_7')
// (19, 6, 'ram/WDATA_3')

reg n2465 = 0;
// (17, 5, 'neigh_op_tnr_1')
// (17, 5, 'sp4_r_v_b_47')
// (17, 6, 'neigh_op_rgt_1')
// (17, 6, 'sp4_r_v_b_34')
// (17, 7, 'neigh_op_bnr_1')
// (17, 7, 'sp4_r_v_b_23')
// (17, 8, 'sp4_r_v_b_10')
// (18, 4, 'sp4_v_t_47')
// (18, 5, 'neigh_op_top_1')
// (18, 5, 'sp4_v_b_47')
// (18, 6, 'local_g2_1')
// (18, 6, 'lutff_1/in_2')
// (18, 6, 'lutff_1/out')
// (18, 6, 'sp4_v_b_34')
// (18, 7, 'neigh_op_bot_1')
// (18, 7, 'sp4_v_b_23')
// (18, 8, 'sp4_h_r_4')
// (18, 8, 'sp4_v_b_10')
// (19, 5, 'neigh_op_tnl_1')
// (19, 6, 'local_g1_1')
// (19, 6, 'neigh_op_lft_1')
// (19, 6, 'ram/WADDR_1')
// (19, 7, 'neigh_op_bnl_1')
// (19, 8, 'local_g1_1')
// (19, 8, 'ram/WADDR_1')
// (19, 8, 'sp4_h_r_17')
// (20, 8, 'sp4_h_r_28')
// (21, 8, 'sp4_h_r_41')
// (22, 8, 'sp4_h_l_41')

reg n2466 = 0;
// (17, 5, 'neigh_op_tnr_2')
// (17, 6, 'neigh_op_rgt_2')
// (17, 7, 'neigh_op_bnr_2')
// (18, 4, 'sp4_r_v_b_45')
// (18, 5, 'neigh_op_top_2')
// (18, 5, 'sp4_r_v_b_32')
// (18, 6, 'local_g3_2')
// (18, 6, 'lutff_2/in_1')
// (18, 6, 'lutff_2/out')
// (18, 6, 'sp4_r_v_b_21')
// (18, 7, 'neigh_op_bot_2')
// (18, 7, 'sp4_r_v_b_8')
// (18, 8, 'sp4_r_v_b_45')
// (18, 9, 'sp4_r_v_b_32')
// (18, 10, 'sp4_r_v_b_21')
// (18, 11, 'sp4_r_v_b_8')
// (19, 3, 'sp4_v_t_45')
// (19, 4, 'sp4_v_b_45')
// (19, 5, 'neigh_op_tnl_2')
// (19, 5, 'sp4_v_b_32')
// (19, 6, 'local_g1_2')
// (19, 6, 'neigh_op_lft_2')
// (19, 6, 'ram/WADDR_2')
// (19, 6, 'sp4_v_b_21')
// (19, 7, 'neigh_op_bnl_2')
// (19, 7, 'sp4_v_b_8')
// (19, 7, 'sp4_v_t_45')
// (19, 8, 'local_g2_5')
// (19, 8, 'ram/WADDR_2')
// (19, 8, 'sp4_v_b_45')
// (19, 9, 'sp4_v_b_32')
// (19, 10, 'sp4_v_b_21')
// (19, 11, 'sp4_v_b_8')

reg n2467 = 0;
// (17, 5, 'neigh_op_tnr_3')
// (17, 6, 'neigh_op_rgt_3')
// (17, 7, 'neigh_op_bnr_3')
// (18, 5, 'neigh_op_top_3')
// (18, 6, 'local_g2_3')
// (18, 6, 'lutff_3/in_2')
// (18, 6, 'lutff_3/out')
// (18, 6, 'sp4_r_v_b_39')
// (18, 7, 'neigh_op_bot_3')
// (18, 7, 'sp4_r_v_b_26')
// (18, 8, 'sp4_r_v_b_15')
// (18, 9, 'sp4_r_v_b_2')
// (19, 5, 'neigh_op_tnl_3')
// (19, 5, 'sp4_v_t_39')
// (19, 6, 'local_g1_3')
// (19, 6, 'neigh_op_lft_3')
// (19, 6, 'ram/WADDR_3')
// (19, 6, 'sp4_v_b_39')
// (19, 7, 'neigh_op_bnl_3')
// (19, 7, 'sp4_v_b_26')
// (19, 8, 'local_g1_7')
// (19, 8, 'ram/WADDR_3')
// (19, 8, 'sp4_v_b_15')
// (19, 9, 'sp4_v_b_2')

reg n2468 = 0;
// (17, 5, 'neigh_op_tnr_4')
// (17, 6, 'neigh_op_rgt_4')
// (17, 7, 'neigh_op_bnr_4')
// (18, 5, 'neigh_op_top_4')
// (18, 5, 'sp4_r_v_b_36')
// (18, 6, 'local_g3_4')
// (18, 6, 'lutff_4/in_1')
// (18, 6, 'lutff_4/out')
// (18, 6, 'sp4_r_v_b_25')
// (18, 7, 'neigh_op_bot_4')
// (18, 7, 'sp4_r_v_b_12')
// (18, 8, 'sp4_r_v_b_1')
// (19, 4, 'sp4_v_t_36')
// (19, 5, 'neigh_op_tnl_4')
// (19, 5, 'sp4_v_b_36')
// (19, 6, 'local_g1_4')
// (19, 6, 'neigh_op_lft_4')
// (19, 6, 'ram/WADDR_4')
// (19, 6, 'sp4_v_b_25')
// (19, 7, 'neigh_op_bnl_4')
// (19, 7, 'sp4_v_b_12')
// (19, 8, 'local_g0_1')
// (19, 8, 'ram/WADDR_4')
// (19, 8, 'sp4_v_b_1')

reg n2469 = 0;
// (17, 5, 'neigh_op_tnr_5')
// (17, 6, 'neigh_op_rgt_5')
// (17, 7, 'neigh_op_bnr_5')
// (18, 5, 'neigh_op_top_5')
// (18, 5, 'sp4_r_v_b_38')
// (18, 6, 'local_g1_5')
// (18, 6, 'lutff_5/in_1')
// (18, 6, 'lutff_5/out')
// (18, 6, 'sp4_r_v_b_27')
// (18, 7, 'neigh_op_bot_5')
// (18, 7, 'sp4_r_v_b_14')
// (18, 8, 'sp4_r_v_b_3')
// (19, 4, 'sp4_v_t_38')
// (19, 5, 'neigh_op_tnl_5')
// (19, 5, 'sp4_v_b_38')
// (19, 6, 'local_g1_5')
// (19, 6, 'neigh_op_lft_5')
// (19, 6, 'ram/WADDR_5')
// (19, 6, 'sp4_v_b_27')
// (19, 7, 'neigh_op_bnl_5')
// (19, 7, 'sp4_v_b_14')
// (19, 8, 'local_g1_3')
// (19, 8, 'ram/WADDR_5')
// (19, 8, 'sp4_v_b_3')

reg n2470 = 0;
// (17, 5, 'neigh_op_tnr_6')
// (17, 6, 'neigh_op_rgt_6')
// (17, 6, 'sp4_h_r_1')
// (17, 7, 'neigh_op_bnr_6')
// (18, 5, 'neigh_op_top_6')
// (18, 6, 'local_g3_6')
// (18, 6, 'lutff_6/in_1')
// (18, 6, 'lutff_6/out')
// (18, 6, 'sp4_h_r_12')
// (18, 6, 'sp4_r_v_b_45')
// (18, 7, 'neigh_op_bot_6')
// (18, 7, 'sp4_r_v_b_32')
// (18, 8, 'sp4_r_v_b_21')
// (18, 9, 'sp4_r_v_b_8')
// (19, 5, 'neigh_op_tnl_6')
// (19, 5, 'sp4_v_t_45')
// (19, 6, 'local_g2_1')
// (19, 6, 'neigh_op_lft_6')
// (19, 6, 'ram/WADDR_6')
// (19, 6, 'sp4_h_r_25')
// (19, 6, 'sp4_v_b_45')
// (19, 7, 'neigh_op_bnl_6')
// (19, 7, 'sp4_v_b_32')
// (19, 8, 'local_g0_5')
// (19, 8, 'ram/WADDR_6')
// (19, 8, 'sp4_v_b_21')
// (19, 9, 'sp4_v_b_8')
// (20, 6, 'sp4_h_r_36')
// (21, 6, 'sp4_h_l_36')

wire n2471;
// (17, 5, 'sp4_h_r_11')
// (18, 5, 'sp4_h_r_22')
// (19, 4, 'neigh_op_tnr_7')
// (19, 5, 'neigh_op_rgt_7')
// (19, 5, 'sp4_h_r_35')
// (19, 6, 'neigh_op_bnr_7')
// (20, 2, 'sp4_r_v_b_40')
// (20, 3, 'sp4_r_v_b_29')
// (20, 4, 'neigh_op_top_7')
// (20, 4, 'sp4_r_v_b_16')
// (20, 5, 'local_g1_5')
// (20, 5, 'lutff_7/out')
// (20, 5, 'lutff_global/s_r')
// (20, 5, 'sp4_h_r_46')
// (20, 5, 'sp4_r_v_b_5')
// (20, 6, 'neigh_op_bot_7')
// (21, 1, 'sp4_v_t_40')
// (21, 2, 'sp4_v_b_40')
// (21, 3, 'sp4_v_b_29')
// (21, 4, 'neigh_op_tnl_7')
// (21, 4, 'sp4_v_b_16')
// (21, 5, 'neigh_op_lft_7')
// (21, 5, 'sp4_h_l_46')
// (21, 5, 'sp4_v_b_5')
// (21, 6, 'neigh_op_bnl_7')

wire n2472;
// (17, 5, 'sp4_h_r_6')
// (18, 5, 'sp4_h_r_19')
// (19, 5, 'sp4_h_r_30')
// (20, 5, 'local_g3_3')
// (20, 5, 'lutff_global/cen')
// (20, 5, 'sp4_h_r_43')
// (21, 4, 'neigh_op_tnr_7')
// (21, 5, 'neigh_op_rgt_7')
// (21, 5, 'sp4_h_l_43')
// (21, 5, 'sp4_h_r_3')
// (21, 6, 'neigh_op_bnr_7')
// (22, 4, 'neigh_op_top_7')
// (22, 5, 'lutff_7/out')
// (22, 5, 'sp4_h_r_14')
// (22, 6, 'neigh_op_bot_7')
// (23, 4, 'neigh_op_tnl_7')
// (23, 5, 'neigh_op_lft_7')
// (23, 5, 'sp4_h_r_27')
// (23, 6, 'neigh_op_bnl_7')
// (24, 5, 'sp4_h_r_38')
// (25, 5, 'sp4_h_l_38')

wire n2473;
// (17, 6, 'lutff_0/cout')
// (17, 6, 'lutff_1/in_3')

wire n2474;
// (17, 6, 'lutff_2/cout')
// (17, 6, 'lutff_3/in_3')

wire n2475;
// (17, 6, 'lutff_4/cout')
// (17, 6, 'lutff_5/in_3')

wire n2476;
// (17, 6, 'lutff_6/cout')
// (17, 6, 'lutff_7/in_3')

wire n2477;
// (17, 6, 'lutff_7/cout')
// (17, 7, 'carry_in')
// (17, 7, 'carry_in_mux')

reg n2478 = 0;
// (17, 6, 'neigh_op_tnr_2')
// (17, 7, 'neigh_op_rgt_2')
// (17, 7, 'sp4_r_v_b_36')
// (17, 8, 'neigh_op_bnr_2')
// (17, 8, 'sp4_r_v_b_25')
// (17, 9, 'sp4_r_v_b_12')
// (17, 10, 'sp4_r_v_b_1')
// (18, 6, 'neigh_op_top_2')
// (18, 6, 'sp4_v_t_36')
// (18, 7, 'lutff_2/out')
// (18, 7, 'sp4_v_b_36')
// (18, 8, 'neigh_op_bot_2')
// (18, 8, 'sp4_v_b_25')
// (18, 9, 'local_g0_4')
// (18, 9, 'lutff_7/in_3')
// (18, 9, 'sp4_v_b_12')
// (18, 10, 'sp4_v_b_1')
// (19, 6, 'neigh_op_tnl_2')
// (19, 7, 'neigh_op_lft_2')
// (19, 8, 'neigh_op_bnl_2')

reg n2479 = 0;
// (17, 6, 'neigh_op_tnr_3')
// (17, 7, 'neigh_op_rgt_3')
// (17, 7, 'sp4_r_v_b_38')
// (17, 8, 'neigh_op_bnr_3')
// (17, 8, 'sp4_r_v_b_27')
// (17, 9, 'sp4_r_v_b_14')
// (17, 10, 'sp4_r_v_b_3')
// (18, 6, 'neigh_op_top_3')
// (18, 6, 'sp4_v_t_38')
// (18, 7, 'lutff_3/out')
// (18, 7, 'sp4_v_b_38')
// (18, 8, 'neigh_op_bot_3')
// (18, 8, 'sp4_v_b_27')
// (18, 9, 'sp4_v_b_14')
// (18, 10, 'local_g0_3')
// (18, 10, 'lutff_1/in_0')
// (18, 10, 'sp4_v_b_3')
// (19, 6, 'neigh_op_tnl_3')
// (19, 7, 'neigh_op_lft_3')
// (19, 8, 'neigh_op_bnl_3')

reg n2480 = 0;
// (17, 6, 'neigh_op_tnr_5')
// (17, 7, 'neigh_op_rgt_5')
// (17, 7, 'sp4_r_v_b_42')
// (17, 8, 'neigh_op_bnr_5')
// (17, 8, 'sp4_r_v_b_31')
// (17, 9, 'sp4_r_v_b_18')
// (17, 10, 'sp4_r_v_b_7')
// (18, 6, 'neigh_op_top_5')
// (18, 6, 'sp4_v_t_42')
// (18, 7, 'lutff_5/out')
// (18, 7, 'sp4_v_b_42')
// (18, 8, 'neigh_op_bot_5')
// (18, 8, 'sp4_v_b_31')
// (18, 9, 'sp4_v_b_18')
// (18, 10, 'local_g0_7')
// (18, 10, 'lutff_3/in_2')
// (18, 10, 'sp4_v_b_7')
// (19, 6, 'neigh_op_tnl_5')
// (19, 7, 'neigh_op_lft_5')
// (19, 8, 'neigh_op_bnl_5')

reg n2481 = 0;
// (17, 6, 'sp4_h_r_2')
// (18, 6, 'local_g1_7')
// (18, 6, 'lutff_0/in_2')
// (18, 6, 'lutff_1/in_3')
// (18, 6, 'sp4_h_r_15')
// (19, 2, 'sp4_r_v_b_40')
// (19, 3, 'neigh_op_tnr_0')
// (19, 3, 'sp4_r_v_b_29')
// (19, 4, 'neigh_op_rgt_0')
// (19, 4, 'sp4_r_v_b_16')
// (19, 5, 'neigh_op_bnr_0')
// (19, 5, 'sp4_r_v_b_5')
// (19, 6, 'local_g3_0')
// (19, 6, 'ram/WADDR_0')
// (19, 6, 'sp4_h_r_26')
// (19, 6, 'sp4_r_v_b_40')
// (19, 7, 'sp4_r_v_b_29')
// (19, 8, 'local_g3_0')
// (19, 8, 'ram/WADDR_0')
// (19, 8, 'sp4_r_v_b_16')
// (19, 9, 'sp4_r_v_b_5')
// (20, 1, 'sp4_v_t_40')
// (20, 2, 'sp4_v_b_40')
// (20, 3, 'neigh_op_top_0')
// (20, 3, 'sp4_r_v_b_44')
// (20, 3, 'sp4_v_b_29')
// (20, 4, 'local_g0_0')
// (20, 4, 'lutff_0/in_2')
// (20, 4, 'lutff_0/out')
// (20, 4, 'sp4_r_v_b_33')
// (20, 4, 'sp4_v_b_16')
// (20, 5, 'neigh_op_bot_0')
// (20, 5, 'sp4_r_v_b_20')
// (20, 5, 'sp4_v_b_5')
// (20, 5, 'sp4_v_t_40')
// (20, 6, 'sp4_h_r_39')
// (20, 6, 'sp4_r_v_b_9')
// (20, 6, 'sp4_v_b_40')
// (20, 7, 'sp4_v_b_29')
// (20, 8, 'sp4_v_b_16')
// (20, 9, 'sp4_v_b_5')
// (21, 2, 'sp4_v_t_44')
// (21, 3, 'neigh_op_tnl_0')
// (21, 3, 'sp4_v_b_44')
// (21, 4, 'neigh_op_lft_0')
// (21, 4, 'sp4_v_b_33')
// (21, 5, 'neigh_op_bnl_0')
// (21, 5, 'sp4_v_b_20')
// (21, 6, 'sp4_h_l_39')
// (21, 6, 'sp4_v_b_9')

wire n2482;
// (17, 6, 'sp4_h_r_4')
// (18, 5, 'neigh_op_tnr_6')
// (18, 6, 'neigh_op_rgt_6')
// (18, 6, 'sp4_h_r_17')
// (18, 7, 'neigh_op_bnr_6')
// (19, 5, 'neigh_op_top_6')
// (19, 6, 'ram/RDATA_1')
// (19, 6, 'sp4_h_r_28')
// (19, 7, 'neigh_op_bot_6')
// (20, 5, 'neigh_op_tnl_6')
// (20, 6, 'neigh_op_lft_6')
// (20, 6, 'sp4_h_r_41')
// (20, 7, 'neigh_op_bnl_6')
// (21, 6, 'local_g1_0')
// (21, 6, 'lutff_5/in_0')
// (21, 6, 'sp4_h_l_41')
// (21, 6, 'sp4_h_r_0')
// (22, 6, 'sp4_h_r_13')
// (23, 6, 'sp4_h_r_24')
// (24, 6, 'sp4_h_r_37')
// (25, 6, 'sp4_h_l_37')

reg n2483 = 0;
// (17, 6, 'sp4_r_v_b_37')
// (17, 7, 'sp4_r_v_b_24')
// (17, 8, 'local_g2_5')
// (17, 8, 'lutff_4/in_1')
// (17, 8, 'sp4_r_v_b_13')
// (17, 9, 'sp4_r_v_b_0')
// (18, 5, 'sp4_v_t_37')
// (18, 6, 'sp4_v_b_37')
// (18, 7, 'sp4_v_b_24')
// (18, 8, 'sp4_v_b_13')
// (18, 9, 'sp4_h_r_0')
// (18, 9, 'sp4_v_b_0')
// (19, 8, 'neigh_op_tnr_4')
// (19, 9, 'neigh_op_rgt_4')
// (19, 9, 'sp4_h_r_13')
// (19, 10, 'neigh_op_bnr_4')
// (20, 8, 'neigh_op_top_4')
// (20, 9, 'lutff_4/out')
// (20, 9, 'sp4_h_r_24')
// (20, 10, 'neigh_op_bot_4')
// (21, 8, 'neigh_op_tnl_4')
// (21, 9, 'neigh_op_lft_4')
// (21, 9, 'sp4_h_r_37')
// (21, 10, 'neigh_op_bnl_4')
// (22, 9, 'sp4_h_l_37')

reg n2484 = 0;
// (17, 7, 'local_g0_3')
// (17, 7, 'lutff_5/in_0')
// (17, 7, 'sp4_h_r_11')
// (18, 7, 'sp4_h_r_22')
// (19, 7, 'sp4_h_r_35')
// (20, 4, 'sp4_r_v_b_46')
// (20, 5, 'neigh_op_tnr_3')
// (20, 5, 'sp4_r_v_b_35')
// (20, 6, 'neigh_op_rgt_3')
// (20, 6, 'sp4_r_v_b_22')
// (20, 6, 'sp4_r_v_b_38')
// (20, 7, 'neigh_op_bnr_3')
// (20, 7, 'sp4_h_r_46')
// (20, 7, 'sp4_r_v_b_11')
// (20, 7, 'sp4_r_v_b_27')
// (20, 8, 'sp4_r_v_b_14')
// (20, 9, 'sp4_r_v_b_3')
// (21, 3, 'sp4_v_t_46')
// (21, 4, 'sp4_v_b_46')
// (21, 5, 'neigh_op_top_3')
// (21, 5, 'sp4_v_b_35')
// (21, 5, 'sp4_v_t_38')
// (21, 6, 'lutff_3/out')
// (21, 6, 'sp4_v_b_22')
// (21, 6, 'sp4_v_b_38')
// (21, 7, 'neigh_op_bot_3')
// (21, 7, 'sp4_h_l_46')
// (21, 7, 'sp4_v_b_11')
// (21, 7, 'sp4_v_b_27')
// (21, 8, 'sp4_v_b_14')
// (21, 9, 'local_g1_3')
// (21, 9, 'lutff_2/in_0')
// (21, 9, 'sp4_v_b_3')
// (22, 5, 'neigh_op_tnl_3')
// (22, 6, 'neigh_op_lft_3')
// (22, 7, 'neigh_op_bnl_3')

wire n2485;
// (17, 7, 'lutff_0/cout')
// (17, 7, 'lutff_1/in_3')

wire n2486;
// (17, 7, 'lutff_2/cout')
// (17, 7, 'lutff_3/in_3')

wire n2487;
// (17, 7, 'lutff_4/cout')
// (17, 7, 'lutff_5/in_3')

reg n2488 = 0;
// (17, 7, 'neigh_op_tnr_0')
// (17, 7, 'sp4_r_v_b_45')
// (17, 8, 'neigh_op_rgt_0')
// (17, 8, 'sp4_r_v_b_32')
// (17, 9, 'neigh_op_bnr_0')
// (17, 9, 'sp4_r_v_b_21')
// (17, 10, 'sp4_r_v_b_8')
// (18, 6, 'sp4_v_t_45')
// (18, 7, 'neigh_op_top_0')
// (18, 7, 'sp4_v_b_45')
// (18, 8, 'lutff_0/out')
// (18, 8, 'sp4_v_b_32')
// (18, 9, 'neigh_op_bot_0')
// (18, 9, 'sp4_v_b_21')
// (18, 10, 'local_g1_0')
// (18, 10, 'lutff_5/in_2')
// (18, 10, 'sp4_v_b_8')
// (19, 7, 'neigh_op_tnl_0')
// (19, 8, 'neigh_op_lft_0')
// (19, 9, 'neigh_op_bnl_0')

reg n2489 = 0;
// (17, 7, 'neigh_op_tnr_5')
// (17, 8, 'neigh_op_rgt_5')
// (17, 9, 'neigh_op_bnr_5')
// (18, 7, 'neigh_op_top_5')
// (18, 8, 'lutff_5/out')
// (18, 9, 'local_g0_5')
// (18, 9, 'lutff_1/in_2')
// (18, 9, 'neigh_op_bot_5')
// (19, 7, 'neigh_op_tnl_5')
// (19, 8, 'neigh_op_lft_5')
// (19, 9, 'neigh_op_bnl_5')

reg n2490 = 0;
// (17, 7, 'neigh_op_tnr_6')
// (17, 7, 'sp4_r_v_b_41')
// (17, 8, 'neigh_op_rgt_6')
// (17, 8, 'sp4_r_v_b_28')
// (17, 9, 'neigh_op_bnr_6')
// (17, 9, 'sp4_r_v_b_17')
// (17, 10, 'local_g1_4')
// (17, 10, 'lutff_4/in_3')
// (17, 10, 'sp4_r_v_b_4')
// (18, 6, 'sp4_v_t_41')
// (18, 7, 'neigh_op_top_6')
// (18, 7, 'sp4_v_b_41')
// (18, 8, 'lutff_6/out')
// (18, 8, 'sp4_v_b_28')
// (18, 9, 'neigh_op_bot_6')
// (18, 9, 'sp4_v_b_17')
// (18, 10, 'sp4_v_b_4')
// (19, 7, 'neigh_op_tnl_6')
// (19, 8, 'neigh_op_lft_6')
// (19, 9, 'neigh_op_bnl_6')

reg n2491 = 0;
// (17, 7, 'neigh_op_tnr_7')
// (17, 8, 'neigh_op_rgt_7')
// (17, 9, 'neigh_op_bnr_7')
// (18, 7, 'neigh_op_top_7')
// (18, 8, 'lutff_7/out')
// (18, 9, 'local_g0_7')
// (18, 9, 'lutff_3/in_2')
// (18, 9, 'neigh_op_bot_7')
// (19, 7, 'neigh_op_tnl_7')
// (19, 8, 'neigh_op_lft_7')
// (19, 9, 'neigh_op_bnl_7')

wire n2492;
// (17, 8, 'neigh_op_tnr_1')
// (17, 9, 'neigh_op_rgt_1')
// (17, 10, 'neigh_op_bnr_1')
// (18, 8, 'neigh_op_top_1')
// (18, 9, 'local_g1_1')
// (18, 9, 'lutff_0/in_2')
// (18, 9, 'lutff_1/out')
// (18, 10, 'neigh_op_bot_1')
// (19, 8, 'neigh_op_tnl_1')
// (19, 9, 'neigh_op_lft_1')
// (19, 10, 'neigh_op_bnl_1')

wire n2493;
// (17, 8, 'neigh_op_tnr_2')
// (17, 9, 'neigh_op_rgt_2')
// (17, 10, 'neigh_op_bnr_2')
// (18, 8, 'neigh_op_top_2')
// (18, 9, 'local_g0_2')
// (18, 9, 'lutff_0/in_0')
// (18, 9, 'lutff_2/out')
// (18, 10, 'neigh_op_bot_2')
// (19, 8, 'neigh_op_tnl_2')
// (19, 9, 'neigh_op_lft_2')
// (19, 10, 'neigh_op_bnl_2')

wire n2494;
// (17, 8, 'neigh_op_tnr_3')
// (17, 9, 'local_g3_3')
// (17, 9, 'lutff_2/in_0')
// (17, 9, 'neigh_op_rgt_3')
// (17, 10, 'neigh_op_bnr_3')
// (18, 8, 'neigh_op_top_3')
// (18, 9, 'lutff_3/out')
// (18, 10, 'neigh_op_bot_3')
// (19, 8, 'neigh_op_tnl_3')
// (19, 9, 'neigh_op_lft_3')
// (19, 10, 'neigh_op_bnl_3')

wire n2495;
// (17, 8, 'neigh_op_tnr_4')
// (17, 9, 'neigh_op_rgt_4')
// (17, 10, 'neigh_op_bnr_4')
// (18, 8, 'neigh_op_top_4')
// (18, 9, 'local_g3_4')
// (18, 9, 'lutff_4/out')
// (18, 9, 'lutff_6/in_3')
// (18, 10, 'neigh_op_bot_4')
// (19, 8, 'neigh_op_tnl_4')
// (19, 9, 'neigh_op_lft_4')
// (19, 10, 'neigh_op_bnl_4')

reg n2496 = 0;
// (17, 8, 'neigh_op_tnr_5')
// (17, 9, 'neigh_op_rgt_5')
// (17, 10, 'neigh_op_bnr_5')
// (18, 8, 'neigh_op_top_5')
// (18, 9, 'local_g1_5')
// (18, 9, 'lutff_2/in_0')
// (18, 9, 'lutff_5/out')
// (18, 10, 'neigh_op_bot_5')
// (19, 8, 'neigh_op_tnl_5')
// (19, 9, 'neigh_op_lft_5')
// (19, 10, 'neigh_op_bnl_5')

wire n2497;
// (17, 8, 'neigh_op_tnr_6')
// (17, 9, 'neigh_op_rgt_6')
// (17, 10, 'neigh_op_bnr_6')
// (18, 8, 'neigh_op_top_6')
// (18, 9, 'local_g1_6')
// (18, 9, 'lutff_0/in_1')
// (18, 9, 'lutff_6/out')
// (18, 10, 'neigh_op_bot_6')
// (19, 8, 'neigh_op_tnl_6')
// (19, 9, 'neigh_op_lft_6')
// (19, 10, 'neigh_op_bnl_6')

wire n2498;
// (17, 8, 'neigh_op_tnr_7')
// (17, 9, 'local_g2_7')
// (17, 9, 'lutff_2/in_1')
// (17, 9, 'neigh_op_rgt_7')
// (17, 10, 'neigh_op_bnr_7')
// (18, 8, 'neigh_op_top_7')
// (18, 9, 'lutff_7/out')
// (18, 10, 'neigh_op_bot_7')
// (19, 8, 'neigh_op_tnl_7')
// (19, 9, 'neigh_op_lft_7')
// (19, 10, 'neigh_op_bnl_7')

reg n2499 = 0;
// (17, 8, 'sp4_r_v_b_37')
// (17, 9, 'sp4_r_v_b_24')
// (17, 10, 'sp4_r_v_b_13')
// (17, 11, 'local_g1_0')
// (17, 11, 'lutff_3/in_2')
// (17, 11, 'sp4_r_v_b_0')
// (18, 7, 'sp4_v_t_37')
// (18, 8, 'sp4_v_b_37')
// (18, 9, 'sp4_v_b_24')
// (18, 10, 'sp4_v_b_13')
// (18, 11, 'sp4_h_r_7')
// (18, 11, 'sp4_v_b_0')
// (19, 11, 'sp4_h_r_18')
// (20, 10, 'neigh_op_tnr_5')
// (20, 11, 'neigh_op_rgt_5')
// (20, 11, 'sp4_h_r_31')
// (20, 12, 'neigh_op_bnr_5')
// (21, 10, 'neigh_op_top_5')
// (21, 11, 'lutff_5/out')
// (21, 11, 'sp4_h_r_42')
// (21, 12, 'neigh_op_bot_5')
// (22, 10, 'neigh_op_tnl_5')
// (22, 11, 'neigh_op_lft_5')
// (22, 11, 'sp4_h_l_42')
// (22, 12, 'neigh_op_bnl_5')

reg n2500 = 0;
// (17, 8, 'sp4_r_v_b_39')
// (17, 9, 'sp4_r_v_b_26')
// (17, 10, 'sp4_r_v_b_15')
// (17, 11, 'sp4_r_v_b_2')
// (18, 7, 'sp4_v_t_39')
// (18, 8, 'sp4_v_b_39')
// (18, 9, 'sp4_r_v_b_41')
// (18, 9, 'sp4_v_b_26')
// (18, 10, 'local_g1_7')
// (18, 10, 'lutff_0/in_2')
// (18, 10, 'sp4_r_v_b_28')
// (18, 10, 'sp4_v_b_15')
// (18, 11, 'local_g0_2')
// (18, 11, 'lutff_1/in_3')
// (18, 11, 'sp4_h_r_2')
// (18, 11, 'sp4_r_v_b_17')
// (18, 11, 'sp4_v_b_2')
// (18, 12, 'local_g1_4')
// (18, 12, 'lutff_1/in_0')
// (18, 12, 'lutff_7/in_0')
// (18, 12, 'sp4_r_v_b_4')
// (19, 8, 'sp4_v_t_41')
// (19, 9, 'sp4_v_b_41')
// (19, 10, 'sp4_v_b_28')
// (19, 11, 'sp4_h_r_15')
// (19, 11, 'sp4_v_b_17')
// (19, 12, 'sp4_h_r_4')
// (19, 12, 'sp4_r_v_b_44')
// (19, 12, 'sp4_v_b_4')
// (19, 13, 'sp4_r_v_b_33')
// (19, 14, 'sp4_r_v_b_20')
// (19, 15, 'sp4_r_v_b_9')
// (20, 11, 'sp4_h_r_26')
// (20, 11, 'sp4_h_r_3')
// (20, 11, 'sp4_v_t_44')
// (20, 12, 'local_g1_1')
// (20, 12, 'lutff_1/in_3')
// (20, 12, 'lutff_6/in_2')
// (20, 12, 'sp4_h_r_17')
// (20, 12, 'sp4_h_r_3')
// (20, 12, 'sp4_v_b_44')
// (20, 13, 'local_g2_1')
// (20, 13, 'local_g3_1')
// (20, 13, 'lutff_1/in_3')
// (20, 13, 'lutff_2/in_3')
// (20, 13, 'lutff_6/in_3')
// (20, 13, 'lutff_7/in_2')
// (20, 13, 'sp4_v_b_33')
// (20, 14, 'sp4_v_b_20')
// (20, 15, 'sp4_v_b_9')
// (21, 11, 'sp4_h_r_14')
// (21, 11, 'sp4_h_r_39')
// (21, 12, 'local_g1_6')
// (21, 12, 'lutff_3/in_2')
// (21, 12, 'sp4_h_r_14')
// (21, 12, 'sp4_h_r_28')
// (22, 9, 'sp4_r_v_b_46')
// (22, 10, 'neigh_op_tnr_3')
// (22, 10, 'sp4_r_v_b_35')
// (22, 11, 'neigh_op_rgt_3')
// (22, 11, 'sp4_h_l_39')
// (22, 11, 'sp4_h_r_11')
// (22, 11, 'sp4_h_r_27')
// (22, 11, 'sp4_r_v_b_22')
// (22, 12, 'local_g1_3')
// (22, 12, 'lutff_4/in_0')
// (22, 12, 'lutff_7/in_1')
// (22, 12, 'neigh_op_bnr_3')
// (22, 12, 'sp4_h_r_27')
// (22, 12, 'sp4_h_r_41')
// (22, 12, 'sp4_r_v_b_11')
// (23, 8, 'sp4_v_t_46')
// (23, 9, 'sp4_r_v_b_47')
// (23, 9, 'sp4_v_b_46')
// (23, 10, 'neigh_op_top_3')
// (23, 10, 'sp4_r_v_b_34')
// (23, 10, 'sp4_v_b_35')
// (23, 11, 'local_g2_3')
// (23, 11, 'lutff_3/in_2')
// (23, 11, 'lutff_3/out')
// (23, 11, 'sp4_h_r_22')
// (23, 11, 'sp4_h_r_38')
// (23, 11, 'sp4_r_v_b_23')
// (23, 11, 'sp4_v_b_22')
// (23, 12, 'local_g0_3')
// (23, 12, 'local_g1_3')
// (23, 12, 'lutff_0/in_1')
// (23, 12, 'lutff_1/in_3')
// (23, 12, 'neigh_op_bot_3')
// (23, 12, 'sp4_h_l_41')
// (23, 12, 'sp4_h_r_38')
// (23, 12, 'sp4_r_v_b_10')
// (23, 12, 'sp4_v_b_11')
// (24, 8, 'sp4_v_t_47')
// (24, 9, 'sp4_v_b_47')
// (24, 10, 'neigh_op_tnl_3')
// (24, 10, 'sp4_v_b_34')
// (24, 11, 'neigh_op_lft_3')
// (24, 11, 'sp4_h_l_38')
// (24, 11, 'sp4_h_r_35')
// (24, 11, 'sp4_v_b_23')
// (24, 12, 'neigh_op_bnl_3')
// (24, 12, 'sp4_h_l_38')
// (24, 12, 'sp4_v_b_10')
// (25, 11, 'sp4_h_r_46')

reg n2501 = 0;
// (17, 8, 'sp4_r_v_b_40')
// (17, 9, 'sp4_r_v_b_29')
// (17, 10, 'sp4_r_v_b_16')
// (17, 11, 'sp4_r_v_b_5')
// (18, 7, 'sp4_v_t_40')
// (18, 8, 'sp4_v_b_40')
// (18, 9, 'local_g2_5')
// (18, 9, 'lutff_2/in_1')
// (18, 9, 'sp4_v_b_29')
// (18, 10, 'sp4_v_b_16')
// (18, 11, 'sp4_h_r_5')
// (18, 11, 'sp4_v_b_5')
// (19, 11, 'sp4_h_r_16')
// (20, 10, 'neigh_op_tnr_4')
// (20, 11, 'neigh_op_rgt_4')
// (20, 11, 'sp4_h_r_29')
// (20, 12, 'neigh_op_bnr_4')
// (21, 10, 'neigh_op_top_4')
// (21, 11, 'lutff_4/out')
// (21, 11, 'sp4_h_r_40')
// (21, 12, 'neigh_op_bot_4')
// (22, 10, 'neigh_op_tnl_4')
// (22, 11, 'neigh_op_lft_4')
// (22, 11, 'sp4_h_l_40')
// (22, 12, 'neigh_op_bnl_4')

reg n2502 = 0;
// (17, 9, 'local_g1_3')
// (17, 9, 'lutff_3/in_1')
// (17, 9, 'sp4_h_r_11')
// (18, 9, 'sp4_h_r_22')
// (19, 8, 'neigh_op_tnr_7')
// (19, 9, 'neigh_op_rgt_7')
// (19, 9, 'sp4_h_r_35')
// (19, 10, 'neigh_op_bnr_7')
// (20, 8, 'neigh_op_top_7')
// (20, 9, 'lutff_7/out')
// (20, 9, 'sp4_h_r_46')
// (20, 10, 'neigh_op_bot_7')
// (21, 8, 'neigh_op_tnl_7')
// (21, 9, 'neigh_op_lft_7')
// (21, 9, 'sp4_h_l_46')
// (21, 10, 'neigh_op_bnl_7')

wire n2503;
// (17, 9, 'neigh_op_tnr_0')
// (17, 10, 'neigh_op_rgt_0')
// (17, 11, 'neigh_op_bnr_0')
// (18, 9, 'neigh_op_top_0')
// (18, 10, 'lutff_0/out')
// (18, 10, 'sp4_h_r_0')
// (18, 11, 'neigh_op_bot_0')
// (19, 9, 'neigh_op_tnl_0')
// (19, 10, 'neigh_op_lft_0')
// (19, 10, 'sp4_h_r_13')
// (19, 11, 'neigh_op_bnl_0')
// (20, 10, 'sp4_h_r_24')
// (21, 10, 'sp4_h_r_37')
// (21, 11, 'sp4_r_v_b_37')
// (21, 12, 'local_g1_0')
// (21, 12, 'lutff_2/in_1')
// (21, 12, 'sp4_r_v_b_24')
// (21, 13, 'sp4_r_v_b_13')
// (21, 14, 'sp4_r_v_b_0')
// (22, 10, 'sp4_h_l_37')
// (22, 10, 'sp4_v_t_37')
// (22, 11, 'sp4_v_b_37')
// (22, 12, 'sp4_v_b_24')
// (22, 13, 'sp4_v_b_13')
// (22, 14, 'sp4_v_b_0')

wire n2504;
// (17, 9, 'neigh_op_tnr_1')
// (17, 10, 'local_g3_1')
// (17, 10, 'lutff_4/in_0')
// (17, 10, 'neigh_op_rgt_1')
// (17, 11, 'neigh_op_bnr_1')
// (18, 9, 'neigh_op_top_1')
// (18, 10, 'lutff_1/out')
// (18, 11, 'neigh_op_bot_1')
// (19, 9, 'neigh_op_tnl_1')
// (19, 10, 'neigh_op_lft_1')
// (19, 11, 'neigh_op_bnl_1')

wire n2505;
// (17, 9, 'neigh_op_tnr_3')
// (17, 10, 'neigh_op_rgt_3')
// (17, 11, 'neigh_op_bnr_3')
// (18, 9, 'neigh_op_top_3')
// (18, 10, 'local_g2_3')
// (18, 10, 'lutff_2/in_3')
// (18, 10, 'lutff_3/out')
// (18, 11, 'neigh_op_bot_3')
// (19, 9, 'neigh_op_tnl_3')
// (19, 10, 'neigh_op_lft_3')
// (19, 11, 'neigh_op_bnl_3')

wire n2506;
// (17, 9, 'neigh_op_tnr_5')
// (17, 10, 'neigh_op_rgt_5')
// (17, 11, 'neigh_op_bnr_5')
// (18, 9, 'neigh_op_top_5')
// (18, 10, 'local_g1_5')
// (18, 10, 'lutff_2/in_2')
// (18, 10, 'lutff_5/out')
// (18, 11, 'neigh_op_bot_5')
// (19, 9, 'neigh_op_tnl_5')
// (19, 10, 'neigh_op_lft_5')
// (19, 11, 'neigh_op_bnl_5')

wire n2507;
// (17, 9, 'neigh_op_tnr_6')
// (17, 10, 'local_g3_6')
// (17, 10, 'lutff_0/in_1')
// (17, 10, 'lutff_6/in_1')
// (17, 10, 'neigh_op_rgt_6')
// (17, 11, 'neigh_op_bnr_6')
// (18, 9, 'neigh_op_top_6')
// (18, 10, 'lutff_6/out')
// (18, 11, 'neigh_op_bot_6')
// (19, 9, 'neigh_op_tnl_6')
// (19, 10, 'neigh_op_lft_6')
// (19, 11, 'neigh_op_bnl_6')

reg n2508 = 0;
// (17, 9, 'neigh_op_tnr_7')
// (17, 10, 'neigh_op_rgt_7')
// (17, 11, 'neigh_op_bnr_7')
// (18, 9, 'neigh_op_top_7')
// (18, 10, 'lutff_7/out')
// (18, 11, 'local_g1_7')
// (18, 11, 'lutff_3/in_3')
// (18, 11, 'neigh_op_bot_7')
// (19, 9, 'neigh_op_tnl_7')
// (19, 10, 'neigh_op_lft_7')
// (19, 11, 'neigh_op_bnl_7')

reg n2509 = 0;
// (17, 9, 'sp4_r_v_b_37')
// (17, 10, 'sp4_r_v_b_24')
// (17, 11, 'sp4_r_v_b_13')
// (17, 12, 'sp4_r_v_b_0')
// (18, 8, 'sp4_v_t_37')
// (18, 9, 'sp4_v_b_37')
// (18, 10, 'local_g2_0')
// (18, 10, 'lutff_0/in_0')
// (18, 10, 'sp4_v_b_24')
// (18, 11, 'local_g1_5')
// (18, 11, 'lutff_1/in_1')
// (18, 11, 'sp4_v_b_13')
// (18, 12, 'local_g1_0')
// (18, 12, 'lutff_1/in_2')
// (18, 12, 'lutff_7/in_2')
// (18, 12, 'sp4_h_r_0')
// (18, 12, 'sp4_v_b_0')
// (19, 12, 'sp4_h_r_13')
// (20, 12, 'local_g0_1')
// (20, 12, 'lutff_1/in_0')
// (20, 12, 'lutff_6/in_1')
// (20, 12, 'sp4_h_r_1')
// (20, 12, 'sp4_h_r_24')
// (21, 12, 'local_g1_4')
// (21, 12, 'lutff_0/in_3')
// (21, 12, 'lutff_1/in_0')
// (21, 12, 'lutff_2/in_3')
// (21, 12, 'lutff_6/in_3')
// (21, 12, 'lutff_7/in_0')
// (21, 12, 'sp4_h_r_12')
// (21, 12, 'sp4_h_r_37')
// (22, 11, 'neigh_op_tnr_2')
// (22, 12, 'local_g3_2')
// (22, 12, 'lutff_4/in_1')
// (22, 12, 'lutff_7/in_0')
// (22, 12, 'neigh_op_rgt_2')
// (22, 12, 'sp4_h_l_37')
// (22, 12, 'sp4_h_r_25')
// (22, 12, 'sp4_h_r_9')
// (22, 13, 'neigh_op_bnr_2')
// (23, 11, 'neigh_op_top_2')
// (23, 12, 'local_g2_2')
// (23, 12, 'lutff_2/in_0')
// (23, 12, 'lutff_2/out')
// (23, 12, 'sp4_h_r_20')
// (23, 12, 'sp4_h_r_36')
// (23, 13, 'neigh_op_bot_2')
// (24, 11, 'neigh_op_tnl_2')
// (24, 12, 'neigh_op_lft_2')
// (24, 12, 'sp4_h_l_36')
// (24, 12, 'sp4_h_r_33')
// (24, 13, 'neigh_op_bnl_2')
// (25, 12, 'sp4_h_r_44')

wire n2510;
// (17, 10, 'lutff_0/cout')
// (17, 10, 'lutff_1/in_3')

wire n2511;
// (17, 10, 'lutff_1/cout')
// (17, 10, 'lutff_2/in_3')

reg n2512 = 0;
// (17, 10, 'neigh_op_tnr_0')
// (17, 11, 'neigh_op_rgt_0')
// (17, 12, 'neigh_op_bnr_0')
// (18, 10, 'neigh_op_top_0')
// (18, 11, 'local_g1_0')
// (18, 11, 'lutff_0/out')
// (18, 11, 'lutff_1/in_2')
// (18, 12, 'neigh_op_bot_0')
// (19, 10, 'neigh_op_tnl_0')
// (19, 11, 'neigh_op_lft_0')
// (19, 12, 'neigh_op_bnl_0')

wire n2513;
// (17, 10, 'neigh_op_tnr_1')
// (17, 11, 'neigh_op_rgt_1')
// (17, 12, 'neigh_op_bnr_1')
// (18, 9, 'sp4_r_v_b_43')
// (18, 10, 'neigh_op_top_1')
// (18, 10, 'sp4_r_v_b_30')
// (18, 11, 'lutff_1/out')
// (18, 11, 'sp4_r_v_b_19')
// (18, 12, 'neigh_op_bot_1')
// (18, 12, 'sp4_r_v_b_6')
// (19, 8, 'sp4_v_t_43')
// (19, 9, 'sp4_v_b_43')
// (19, 10, 'neigh_op_tnl_1')
// (19, 10, 'sp4_v_b_30')
// (19, 11, 'neigh_op_lft_1')
// (19, 11, 'sp4_v_b_19')
// (19, 12, 'neigh_op_bnl_1')
// (19, 12, 'sp4_h_r_0')
// (19, 12, 'sp4_v_b_6')
// (20, 12, 'sp4_h_r_13')
// (21, 12, 'local_g3_0')
// (21, 12, 'lutff_0/in_1')
// (21, 12, 'sp4_h_r_24')
// (22, 12, 'sp4_h_r_37')
// (23, 12, 'sp4_h_l_37')

wire n2514;
// (17, 10, 'neigh_op_tnr_2')
// (17, 11, 'local_g2_2')
// (17, 11, 'lutff_7/in_1')
// (17, 11, 'neigh_op_rgt_2')
// (17, 12, 'neigh_op_bnr_2')
// (18, 10, 'neigh_op_top_2')
// (18, 11, 'lutff_2/out')
// (18, 12, 'neigh_op_bot_2')
// (19, 10, 'neigh_op_tnl_2')
// (19, 11, 'neigh_op_lft_2')
// (19, 12, 'neigh_op_bnl_2')

wire n2515;
// (17, 10, 'neigh_op_tnr_3')
// (17, 11, 'local_g3_3')
// (17, 11, 'lutff_7/in_3')
// (17, 11, 'neigh_op_rgt_3')
// (17, 12, 'neigh_op_bnr_3')
// (18, 10, 'neigh_op_top_3')
// (18, 11, 'lutff_3/out')
// (18, 12, 'neigh_op_bot_3')
// (19, 10, 'neigh_op_tnl_3')
// (19, 11, 'neigh_op_lft_3')
// (19, 12, 'neigh_op_bnl_3')

reg n2516 = 0;
// (17, 10, 'neigh_op_tnr_4')
// (17, 11, 'neigh_op_rgt_4')
// (17, 12, 'neigh_op_bnr_4')
// (18, 10, 'local_g1_4')
// (18, 10, 'lutff_0/in_1')
// (18, 10, 'neigh_op_top_4')
// (18, 11, 'lutff_4/out')
// (18, 12, 'neigh_op_bot_4')
// (19, 10, 'neigh_op_tnl_4')
// (19, 11, 'neigh_op_lft_4')
// (19, 12, 'neigh_op_bnl_4')

reg n2517 = 0;
// (17, 10, 'neigh_op_tnr_5')
// (17, 11, 'neigh_op_rgt_5')
// (17, 12, 'neigh_op_bnr_5')
// (18, 10, 'neigh_op_top_5')
// (18, 11, 'lutff_5/out')
// (18, 11, 'sp4_h_r_10')
// (18, 12, 'neigh_op_bot_5')
// (19, 10, 'neigh_op_tnl_5')
// (19, 11, 'neigh_op_lft_5')
// (19, 11, 'sp4_h_r_23')
// (19, 12, 'neigh_op_bnl_5')
// (20, 11, 'local_g2_2')
// (20, 11, 'lutff_7/in_3')
// (20, 11, 'sp4_h_r_34')
// (21, 11, 'sp4_h_r_47')
// (22, 11, 'sp4_h_l_47')

reg n2518 = 0;
// (17, 10, 'neigh_op_tnr_6')
// (17, 11, 'neigh_op_rgt_6')
// (17, 12, 'neigh_op_bnr_6')
// (18, 10, 'local_g3_0')
// (18, 10, 'lutff_0/in_3')
// (18, 10, 'neigh_op_top_6')
// (18, 10, 'sp4_r_v_b_40')
// (18, 11, 'lutff_6/out')
// (18, 11, 'sp4_r_v_b_29')
// (18, 12, 'neigh_op_bot_6')
// (18, 12, 'sp4_r_v_b_16')
// (18, 13, 'sp4_r_v_b_5')
// (19, 9, 'sp4_v_t_40')
// (19, 10, 'neigh_op_tnl_6')
// (19, 10, 'sp4_v_b_40')
// (19, 11, 'neigh_op_lft_6')
// (19, 11, 'sp4_v_b_29')
// (19, 12, 'neigh_op_bnl_6')
// (19, 12, 'sp4_v_b_16')
// (19, 13, 'sp4_v_b_5')

reg n2519 = 0;
// (17, 10, 'neigh_op_tnr_7')
// (17, 11, 'neigh_op_rgt_7')
// (17, 12, 'neigh_op_bnr_7')
// (18, 10, 'neigh_op_top_7')
// (18, 11, 'local_g0_7')
// (18, 11, 'lutff_1/in_0')
// (18, 11, 'lutff_7/out')
// (18, 12, 'neigh_op_bot_7')
// (19, 10, 'neigh_op_tnl_7')
// (19, 11, 'neigh_op_lft_7')
// (19, 12, 'neigh_op_bnl_7')

wire n2520;
// (17, 11, 'lutff_1/cout')
// (17, 11, 'lutff_2/in_3')

reg n2521 = 0;
// (17, 11, 'neigh_op_tnr_0')
// (17, 12, 'neigh_op_rgt_0')
// (17, 13, 'neigh_op_bnr_0')
// (18, 11, 'neigh_op_top_0')
// (18, 12, 'local_g2_0')
// (18, 12, 'lutff_0/out')
// (18, 12, 'lutff_7/in_3')
// (18, 13, 'neigh_op_bot_0')
// (19, 11, 'neigh_op_tnl_0')
// (19, 12, 'neigh_op_lft_0')
// (19, 13, 'neigh_op_bnl_0')

wire n2522;
// (17, 11, 'neigh_op_tnr_1')
// (17, 12, 'neigh_op_rgt_1')
// (17, 13, 'neigh_op_bnr_1')
// (18, 11, 'neigh_op_top_1')
// (18, 12, 'lutff_1/out')
// (18, 12, 'sp4_h_r_2')
// (18, 13, 'neigh_op_bot_1')
// (19, 11, 'neigh_op_tnl_1')
// (19, 12, 'neigh_op_lft_1')
// (19, 12, 'sp4_h_r_15')
// (19, 13, 'neigh_op_bnl_1')
// (20, 12, 'sp4_h_r_26')
// (21, 12, 'local_g2_7')
// (21, 12, 'lutff_7/in_2')
// (21, 12, 'sp4_h_r_39')
// (22, 12, 'sp4_h_l_39')

reg n2523 = 0;
// (17, 11, 'neigh_op_tnr_2')
// (17, 12, 'neigh_op_rgt_2')
// (17, 13, 'neigh_op_bnr_2')
// (18, 10, 'sp4_r_v_b_45')
// (18, 11, 'neigh_op_top_2')
// (18, 11, 'sp4_r_v_b_32')
// (18, 12, 'lutff_2/out')
// (18, 12, 'sp4_r_v_b_21')
// (18, 13, 'neigh_op_bot_2')
// (18, 13, 'sp4_r_v_b_8')
// (19, 9, 'sp4_v_t_45')
// (19, 10, 'sp4_v_b_45')
// (19, 11, 'neigh_op_tnl_2')
// (19, 11, 'sp4_v_b_32')
// (19, 12, 'neigh_op_lft_2')
// (19, 12, 'sp4_v_b_21')
// (19, 13, 'neigh_op_bnl_2')
// (19, 13, 'sp4_h_r_8')
// (19, 13, 'sp4_v_b_8')
// (20, 13, 'local_g1_5')
// (20, 13, 'lutff_5/in_3')
// (20, 13, 'sp4_h_r_21')
// (21, 13, 'sp4_h_r_32')
// (22, 13, 'sp4_h_r_45')
// (23, 13, 'sp4_h_l_45')

reg n2524 = 0;
// (17, 11, 'neigh_op_tnr_3')
// (17, 12, 'neigh_op_rgt_3')
// (17, 13, 'neigh_op_bnr_3')
// (18, 10, 'sp4_r_v_b_47')
// (18, 11, 'neigh_op_top_3')
// (18, 11, 'sp4_r_v_b_34')
// (18, 12, 'lutff_3/out')
// (18, 12, 'sp4_r_v_b_23')
// (18, 13, 'neigh_op_bot_3')
// (18, 13, 'sp4_r_v_b_10')
// (19, 9, 'sp4_v_t_47')
// (19, 10, 'sp4_v_b_47')
// (19, 11, 'neigh_op_tnl_3')
// (19, 11, 'sp4_v_b_34')
// (19, 12, 'neigh_op_lft_3')
// (19, 12, 'sp4_v_b_23')
// (19, 13, 'neigh_op_bnl_3')
// (19, 13, 'sp4_h_r_10')
// (19, 13, 'sp4_v_b_10')
// (20, 13, 'local_g1_7')
// (20, 13, 'lutff_4/in_0')
// (20, 13, 'sp4_h_r_23')
// (21, 13, 'sp4_h_r_34')
// (22, 13, 'sp4_h_r_47')
// (23, 13, 'sp4_h_l_47')

reg n2525 = 0;
// (17, 11, 'neigh_op_tnr_4')
// (17, 12, 'neigh_op_rgt_4')
// (17, 13, 'neigh_op_bnr_4')
// (18, 11, 'neigh_op_top_4')
// (18, 12, 'lutff_4/out')
// (18, 12, 'sp4_h_r_8')
// (18, 13, 'neigh_op_bot_4')
// (19, 11, 'neigh_op_tnl_4')
// (19, 12, 'neigh_op_lft_4')
// (19, 12, 'sp4_h_r_21')
// (19, 13, 'neigh_op_bnl_4')
// (20, 12, 'sp4_h_r_32')
// (21, 12, 'local_g3_5')
// (21, 12, 'lutff_1/in_1')
// (21, 12, 'sp4_h_r_45')
// (22, 12, 'sp4_h_l_45')

reg n2526 = 0;
// (17, 11, 'neigh_op_tnr_5')
// (17, 12, 'neigh_op_rgt_5')
// (17, 13, 'neigh_op_bnr_5')
// (18, 11, 'neigh_op_top_5')
// (18, 12, 'local_g1_5')
// (18, 12, 'lutff_1/in_1')
// (18, 12, 'lutff_5/out')
// (18, 13, 'neigh_op_bot_5')
// (19, 11, 'neigh_op_tnl_5')
// (19, 12, 'neigh_op_lft_5')
// (19, 13, 'neigh_op_bnl_5')

reg n2527 = 0;
// (17, 11, 'neigh_op_tnr_6')
// (17, 12, 'neigh_op_rgt_6')
// (17, 13, 'neigh_op_bnr_6')
// (18, 11, 'neigh_op_top_6')
// (18, 12, 'local_g0_6')
// (18, 12, 'lutff_1/in_3')
// (18, 12, 'lutff_6/out')
// (18, 13, 'neigh_op_bot_6')
// (19, 11, 'neigh_op_tnl_6')
// (19, 12, 'neigh_op_lft_6')
// (19, 13, 'neigh_op_bnl_6')

reg n2528 = 0;
// (17, 12, 'neigh_op_tnr_0')
// (17, 13, 'neigh_op_rgt_0')
// (17, 14, 'neigh_op_bnr_0')
// (18, 12, 'neigh_op_top_0')
// (18, 13, 'lutff_0/out')
// (18, 13, 'sp4_h_r_0')
// (18, 14, 'neigh_op_bot_0')
// (19, 12, 'neigh_op_tnl_0')
// (19, 13, 'neigh_op_lft_0')
// (19, 13, 'sp4_h_r_13')
// (19, 14, 'neigh_op_bnl_0')
// (20, 13, 'local_g2_0')
// (20, 13, 'lutff_4/in_2')
// (20, 13, 'sp4_h_r_24')
// (21, 13, 'sp4_h_r_37')
// (22, 13, 'sp4_h_l_37')

reg n2529 = 0;
// (17, 12, 'neigh_op_tnr_1')
// (17, 13, 'neigh_op_rgt_1')
// (17, 13, 'sp4_h_r_7')
// (17, 14, 'neigh_op_bnr_1')
// (18, 12, 'neigh_op_top_1')
// (18, 13, 'lutff_1/out')
// (18, 13, 'sp4_h_r_18')
// (18, 14, 'neigh_op_bot_1')
// (19, 12, 'neigh_op_tnl_1')
// (19, 13, 'neigh_op_lft_1')
// (19, 13, 'sp4_h_r_31')
// (19, 14, 'neigh_op_bnl_1')
// (20, 13, 'local_g2_2')
// (20, 13, 'lutff_2/in_2')
// (20, 13, 'sp4_h_r_42')
// (21, 13, 'sp4_h_l_42')

reg n2530 = 0;
// (17, 12, 'neigh_op_tnr_2')
// (17, 13, 'neigh_op_rgt_2')
// (17, 14, 'neigh_op_bnr_2')
// (18, 12, 'neigh_op_top_2')
// (18, 13, 'lutff_2/out')
// (18, 13, 'sp4_h_r_4')
// (18, 14, 'neigh_op_bot_2')
// (19, 12, 'neigh_op_tnl_2')
// (19, 13, 'neigh_op_lft_2')
// (19, 13, 'sp4_h_r_17')
// (19, 14, 'neigh_op_bnl_2')
// (20, 13, 'sp4_h_r_28')
// (21, 13, 'sp4_h_r_41')
// (22, 13, 'local_g1_0')
// (22, 13, 'lutff_2/in_1')
// (22, 13, 'sp4_h_l_41')
// (22, 13, 'sp4_h_r_0')
// (23, 13, 'sp4_h_r_13')
// (24, 13, 'sp4_h_r_24')
// (25, 13, 'sp4_h_r_37')

reg n2531 = 0;
// (17, 12, 'neigh_op_tnr_3')
// (17, 13, 'neigh_op_rgt_3')
// (17, 14, 'neigh_op_bnr_3')
// (18, 12, 'neigh_op_top_3')
// (18, 13, 'lutff_3/out')
// (18, 13, 'sp4_h_r_6')
// (18, 14, 'neigh_op_bot_3')
// (19, 12, 'neigh_op_tnl_3')
// (19, 13, 'neigh_op_lft_3')
// (19, 13, 'sp4_h_r_19')
// (19, 14, 'neigh_op_bnl_3')
// (20, 13, 'local_g3_6')
// (20, 13, 'lutff_7/in_0')
// (20, 13, 'sp4_h_r_30')
// (21, 13, 'sp4_h_r_43')
// (22, 13, 'sp4_h_l_43')

reg n2532 = 0;
// (17, 12, 'neigh_op_tnr_4')
// (17, 13, 'neigh_op_rgt_4')
// (17, 14, 'neigh_op_bnr_4')
// (18, 12, 'neigh_op_top_4')
// (18, 13, 'lutff_4/out')
// (18, 13, 'sp4_h_r_8')
// (18, 14, 'neigh_op_bot_4')
// (19, 12, 'neigh_op_tnl_4')
// (19, 13, 'neigh_op_lft_4')
// (19, 13, 'sp4_h_r_21')
// (19, 14, 'neigh_op_bnl_4')
// (20, 13, 'local_g3_0')
// (20, 13, 'lutff_1/in_2')
// (20, 13, 'sp4_h_r_32')
// (21, 13, 'sp4_h_r_45')
// (22, 13, 'sp4_h_l_45')

reg n2533 = 0;
// (17, 12, 'neigh_op_tnr_5')
// (17, 13, 'neigh_op_rgt_5')
// (17, 14, 'neigh_op_bnr_5')
// (18, 12, 'neigh_op_top_5')
// (18, 13, 'lutff_5/out')
// (18, 13, 'sp4_h_r_10')
// (18, 14, 'neigh_op_bot_5')
// (19, 12, 'neigh_op_tnl_5')
// (19, 13, 'neigh_op_lft_5')
// (19, 13, 'sp4_h_r_23')
// (19, 14, 'neigh_op_bnl_5')
// (20, 13, 'sp4_h_r_34')
// (21, 13, 'sp4_h_r_47')
// (22, 13, 'local_g0_1')
// (22, 13, 'lutff_3/in_2')
// (22, 13, 'sp4_h_l_47')
// (22, 13, 'sp4_h_r_1')
// (23, 13, 'sp4_h_r_12')
// (24, 13, 'sp4_h_r_25')
// (25, 13, 'sp4_h_r_36')

reg n2534 = 0;
// (17, 12, 'neigh_op_tnr_6')
// (17, 13, 'neigh_op_rgt_6')
// (17, 13, 'sp4_h_r_1')
// (17, 14, 'neigh_op_bnr_6')
// (18, 12, 'neigh_op_top_6')
// (18, 13, 'lutff_6/out')
// (18, 13, 'sp4_h_r_12')
// (18, 14, 'neigh_op_bot_6')
// (19, 12, 'neigh_op_tnl_6')
// (19, 13, 'neigh_op_lft_6')
// (19, 13, 'sp4_h_r_25')
// (19, 14, 'neigh_op_bnl_6')
// (20, 13, 'local_g3_4')
// (20, 13, 'lutff_1/in_0')
// (20, 13, 'sp4_h_r_36')
// (21, 13, 'sp4_h_l_36')

reg n2535 = 0;
// (17, 12, 'neigh_op_tnr_7')
// (17, 13, 'neigh_op_rgt_7')
// (17, 13, 'sp4_h_r_3')
// (17, 14, 'neigh_op_bnr_7')
// (18, 12, 'neigh_op_top_7')
// (18, 13, 'lutff_7/out')
// (18, 13, 'sp4_h_r_14')
// (18, 14, 'neigh_op_bot_7')
// (19, 12, 'neigh_op_tnl_7')
// (19, 13, 'neigh_op_lft_7')
// (19, 13, 'sp4_h_r_27')
// (19, 14, 'neigh_op_bnl_7')
// (20, 10, 'sp4_r_v_b_44')
// (20, 11, 'sp4_r_v_b_33')
// (20, 12, 'sp4_r_v_b_20')
// (20, 13, 'sp4_h_r_38')
// (20, 13, 'sp4_r_v_b_9')
// (21, 9, 'sp4_v_t_44')
// (21, 10, 'sp4_v_b_44')
// (21, 11, 'sp4_v_b_33')
// (21, 12, 'local_g0_4')
// (21, 12, 'lutff_7/in_1')
// (21, 12, 'sp4_v_b_20')
// (21, 13, 'sp4_h_l_38')
// (21, 13, 'sp4_v_b_9')

wire n2536;
// (17, 13, 'local_g3_3')
// (17, 13, 'lutff_global/cen')
// (17, 13, 'neigh_op_tnr_3')
// (17, 14, 'neigh_op_rgt_3')
// (17, 15, 'neigh_op_bnr_3')
// (18, 13, 'neigh_op_top_3')
// (18, 14, 'lutff_3/out')
// (18, 15, 'neigh_op_bot_3')
// (19, 13, 'neigh_op_tnl_3')
// (19, 14, 'neigh_op_lft_3')
// (19, 15, 'neigh_op_bnl_3')

wire n2537;
// (17, 13, 'lutff_1/cout')
// (17, 13, 'lutff_2/in_3')

wire n2538;
// (17, 13, 'lutff_2/cout')
// (17, 13, 'lutff_3/in_3')

wire n2539;
// (17, 13, 'lutff_3/cout')
// (17, 13, 'lutff_4/in_3')

wire n2540;
// (17, 13, 'lutff_4/cout')
// (17, 13, 'lutff_5/in_3')

wire n2541;
// (17, 13, 'lutff_5/cout')
// (17, 13, 'lutff_6/in_3')

reg n2542 = 0;
// (17, 13, 'neigh_op_tnr_1')
// (17, 14, 'neigh_op_rgt_1')
// (17, 14, 'sp4_h_r_7')
// (17, 15, 'neigh_op_bnr_1')
// (18, 13, 'neigh_op_top_1')
// (18, 14, 'lutff_1/out')
// (18, 14, 'sp4_h_r_18')
// (18, 15, 'neigh_op_bot_1')
// (19, 13, 'neigh_op_tnl_1')
// (19, 14, 'neigh_op_lft_1')
// (19, 14, 'sp4_h_r_31')
// (19, 15, 'neigh_op_bnl_1')
// (20, 11, 'sp4_r_v_b_36')
// (20, 12, 'sp4_r_v_b_25')
// (20, 13, 'local_g2_4')
// (20, 13, 'lutff_5/in_1')
// (20, 13, 'sp4_r_v_b_12')
// (20, 14, 'sp4_h_r_42')
// (20, 14, 'sp4_r_v_b_1')
// (21, 10, 'sp4_v_t_36')
// (21, 11, 'sp4_v_b_36')
// (21, 12, 'sp4_v_b_25')
// (21, 13, 'sp4_v_b_12')
// (21, 14, 'sp4_h_l_42')
// (21, 14, 'sp4_v_b_1')

reg n2543 = 0;
// (17, 13, 'neigh_op_tnr_2')
// (17, 14, 'neigh_op_rgt_2')
// (17, 14, 'sp4_h_r_9')
// (17, 15, 'neigh_op_bnr_2')
// (18, 13, 'neigh_op_top_2')
// (18, 14, 'lutff_2/out')
// (18, 14, 'sp4_h_r_20')
// (18, 15, 'neigh_op_bot_2')
// (19, 13, 'neigh_op_tnl_2')
// (19, 14, 'neigh_op_lft_2')
// (19, 14, 'sp4_h_r_33')
// (19, 15, 'neigh_op_bnl_2')
// (20, 11, 'sp4_r_v_b_38')
// (20, 12, 'sp4_r_v_b_27')
// (20, 13, 'local_g2_6')
// (20, 13, 'lutff_0/in_2')
// (20, 13, 'sp4_r_v_b_14')
// (20, 14, 'sp4_h_r_44')
// (20, 14, 'sp4_r_v_b_3')
// (21, 10, 'sp4_v_t_38')
// (21, 11, 'sp4_v_b_38')
// (21, 12, 'sp4_v_b_27')
// (21, 13, 'sp4_v_b_14')
// (21, 14, 'sp4_h_l_44')
// (21, 14, 'sp4_v_b_3')

reg n2544 = 0;
// (17, 13, 'neigh_op_tnr_4')
// (17, 14, 'neigh_op_rgt_4')
// (17, 15, 'neigh_op_bnr_4')
// (18, 13, 'neigh_op_top_4')
// (18, 14, 'lutff_4/out')
// (18, 14, 'sp4_r_v_b_41')
// (18, 15, 'neigh_op_bot_4')
// (18, 15, 'sp4_r_v_b_28')
// (18, 16, 'sp4_r_v_b_17')
// (18, 17, 'sp4_r_v_b_4')
// (19, 13, 'neigh_op_tnl_4')
// (19, 13, 'sp4_h_r_9')
// (19, 13, 'sp4_v_t_41')
// (19, 14, 'neigh_op_lft_4')
// (19, 14, 'sp4_v_b_41')
// (19, 15, 'neigh_op_bnl_4')
// (19, 15, 'sp4_v_b_28')
// (19, 16, 'sp4_v_b_17')
// (19, 17, 'sp4_v_b_4')
// (20, 13, 'local_g1_4')
// (20, 13, 'lutff_6/in_1')
// (20, 13, 'sp4_h_r_20')
// (21, 13, 'sp4_h_r_33')
// (22, 13, 'sp4_h_r_44')
// (23, 13, 'sp4_h_l_44')

wire n2545;
// (17, 14, 'lutff_1/cout')
// (17, 14, 'lutff_2/in_3')

wire n2546;
// (17, 14, 'lutff_2/cout')
// (17, 14, 'lutff_3/in_3')

wire n2547;
// (17, 14, 'lutff_3/cout')
// (17, 14, 'lutff_4/in_3')

wire n2548;
// (17, 14, 'lutff_4/cout')
// (17, 14, 'lutff_5/in_3')

wire n2549;
// (17, 14, 'lutff_5/cout')
// (17, 14, 'lutff_6/in_3')

reg n2550 = 0;
// (17, 14, 'neigh_op_tnr_2')
// (17, 15, 'neigh_op_rgt_2')
// (17, 16, 'neigh_op_bnr_2')
// (18, 13, 'sp4_r_v_b_45')
// (18, 14, 'neigh_op_top_2')
// (18, 14, 'sp4_r_v_b_32')
// (18, 15, 'lutff_2/out')
// (18, 15, 'sp4_r_v_b_21')
// (18, 16, 'neigh_op_bot_2')
// (18, 16, 'sp4_r_v_b_8')
// (19, 12, 'sp4_v_t_45')
// (19, 13, 'sp4_v_b_45')
// (19, 14, 'neigh_op_tnl_2')
// (19, 14, 'sp4_v_b_32')
// (19, 15, 'neigh_op_lft_2')
// (19, 15, 'sp4_v_b_21')
// (19, 16, 'neigh_op_bnl_2')
// (19, 16, 'sp4_h_r_2')
// (19, 16, 'sp4_v_b_8')
// (20, 16, 'sp4_h_r_15')
// (21, 16, 'local_g2_2')
// (21, 16, 'lutff_1/in_1')
// (21, 16, 'sp4_h_r_26')
// (22, 16, 'sp4_h_r_39')
// (23, 16, 'sp4_h_l_39')

reg n2551 = 0;
// (17, 15, 'neigh_op_tnr_0')
// (17, 16, 'neigh_op_rgt_0')
// (17, 17, 'local_g1_0')
// (17, 17, 'lutff_7/in_2')
// (17, 17, 'neigh_op_bnr_0')
// (18, 15, 'neigh_op_top_0')
// (18, 16, 'lutff_0/out')
// (18, 17, 'neigh_op_bot_0')
// (19, 15, 'neigh_op_tnl_0')
// (19, 16, 'neigh_op_lft_0')
// (19, 17, 'neigh_op_bnl_0')

reg n2552 = 0;
// (17, 15, 'neigh_op_tnr_1')
// (17, 16, 'neigh_op_rgt_1')
// (17, 17, 'local_g0_1')
// (17, 17, 'lutff_5/in_0')
// (17, 17, 'neigh_op_bnr_1')
// (18, 15, 'neigh_op_top_1')
// (18, 16, 'lutff_1/out')
// (18, 17, 'neigh_op_bot_1')
// (19, 15, 'neigh_op_tnl_1')
// (19, 16, 'neigh_op_lft_1')
// (19, 17, 'neigh_op_bnl_1')

reg n2553 = 0;
// (17, 15, 'neigh_op_tnr_3')
// (17, 16, 'neigh_op_rgt_3')
// (17, 17, 'local_g0_3')
// (17, 17, 'lutff_4/in_1')
// (17, 17, 'neigh_op_bnr_3')
// (18, 15, 'neigh_op_top_3')
// (18, 16, 'lutff_3/out')
// (18, 17, 'neigh_op_bot_3')
// (19, 15, 'neigh_op_tnl_3')
// (19, 16, 'neigh_op_lft_3')
// (19, 17, 'neigh_op_bnl_3')

reg n2554 = 0;
// (17, 15, 'neigh_op_tnr_4')
// (17, 16, 'neigh_op_rgt_4')
// (17, 17, 'local_g1_4')
// (17, 17, 'lutff_1/in_0')
// (17, 17, 'neigh_op_bnr_4')
// (18, 15, 'neigh_op_top_4')
// (18, 16, 'lutff_4/out')
// (18, 17, 'neigh_op_bot_4')
// (19, 15, 'neigh_op_tnl_4')
// (19, 16, 'neigh_op_lft_4')
// (19, 17, 'neigh_op_bnl_4')

reg n2555 = 0;
// (17, 15, 'neigh_op_tnr_5')
// (17, 16, 'neigh_op_rgt_5')
// (17, 17, 'local_g0_5')
// (17, 17, 'lutff_2/in_3')
// (17, 17, 'neigh_op_bnr_5')
// (18, 15, 'neigh_op_top_5')
// (18, 16, 'lutff_5/out')
// (18, 17, 'neigh_op_bot_5')
// (19, 15, 'neigh_op_tnl_5')
// (19, 16, 'neigh_op_lft_5')
// (19, 17, 'neigh_op_bnl_5')

reg n2556 = 0;
// (17, 15, 'neigh_op_tnr_6')
// (17, 16, 'neigh_op_rgt_6')
// (17, 17, 'local_g0_6')
// (17, 17, 'lutff_3/in_1')
// (17, 17, 'neigh_op_bnr_6')
// (18, 15, 'neigh_op_top_6')
// (18, 16, 'lutff_6/out')
// (18, 17, 'neigh_op_bot_6')
// (19, 15, 'neigh_op_tnl_6')
// (19, 16, 'neigh_op_lft_6')
// (19, 17, 'neigh_op_bnl_6')

reg n2557 = 0;
// (17, 16, 'neigh_op_tnr_0')
// (17, 17, 'neigh_op_rgt_0')
// (17, 18, 'neigh_op_bnr_0')
// (18, 16, 'neigh_op_top_0')
// (18, 17, 'local_g3_0')
// (18, 17, 'lutff_0/out')
// (18, 17, 'lutff_2/in_1')
// (18, 18, 'neigh_op_bot_0')
// (19, 16, 'neigh_op_tnl_0')
// (19, 17, 'neigh_op_lft_0')
// (19, 18, 'neigh_op_bnl_0')

wire n2558;
// (17, 16, 'neigh_op_tnr_2')
// (17, 17, 'neigh_op_rgt_2')
// (17, 18, 'neigh_op_bnr_2')
// (18, 16, 'neigh_op_top_2')
// (18, 17, 'local_g3_2')
// (18, 17, 'lutff_2/out')
// (18, 17, 'lutff_6/in_3')
// (18, 18, 'neigh_op_bot_2')
// (19, 16, 'neigh_op_tnl_2')
// (19, 17, 'neigh_op_lft_2')
// (19, 18, 'neigh_op_bnl_2')

wire n2559;
// (17, 16, 'neigh_op_tnr_3')
// (17, 17, 'neigh_op_rgt_3')
// (17, 18, 'neigh_op_bnr_3')
// (18, 16, 'neigh_op_top_3')
// (18, 17, 'local_g3_3')
// (18, 17, 'lutff_3/out')
// (18, 17, 'lutff_global/cen')
// (18, 18, 'neigh_op_bot_3')
// (19, 16, 'neigh_op_tnl_3')
// (19, 17, 'neigh_op_lft_3')
// (19, 18, 'neigh_op_bnl_3')

wire n2560;
// (17, 16, 'neigh_op_tnr_6')
// (17, 17, 'neigh_op_rgt_6')
// (17, 17, 'sp4_h_r_1')
// (17, 18, 'neigh_op_bnr_6')
// (18, 16, 'neigh_op_top_6')
// (18, 17, 'lutff_6/out')
// (18, 17, 'sp4_h_r_12')
// (18, 18, 'neigh_op_bot_6')
// (19, 16, 'neigh_op_tnl_6')
// (19, 17, 'neigh_op_lft_6')
// (19, 17, 'sp4_h_r_25')
// (19, 18, 'neigh_op_bnl_6')
// (20, 17, 'local_g2_4')
// (20, 17, 'lutff_0/in_0')
// (20, 17, 'sp4_h_r_36')
// (21, 17, 'sp4_h_l_36')

reg n2561 = 0;
// (17, 17, 'neigh_op_tnr_0')
// (17, 18, 'neigh_op_rgt_0')
// (17, 19, 'neigh_op_bnr_0')
// (18, 17, 'neigh_op_top_0')
// (18, 18, 'local_g1_0')
// (18, 18, 'lutff_0/out')
// (18, 18, 'lutff_1/in_2')
// (18, 19, 'neigh_op_bot_0')
// (19, 17, 'neigh_op_tnl_0')
// (19, 18, 'neigh_op_lft_0')
// (19, 19, 'neigh_op_bnl_0')

wire n2562;
// (17, 17, 'neigh_op_tnr_1')
// (17, 18, 'neigh_op_rgt_1')
// (17, 19, 'neigh_op_bnr_1')
// (18, 17, 'neigh_op_top_1')
// (18, 18, 'local_g0_1')
// (18, 18, 'lutff_1/out')
// (18, 18, 'lutff_7/in_2')
// (18, 19, 'neigh_op_bot_1')
// (19, 17, 'neigh_op_tnl_1')
// (19, 18, 'neigh_op_lft_1')
// (19, 19, 'neigh_op_bnl_1')

wire n2563;
// (17, 17, 'neigh_op_tnr_2')
// (17, 18, 'neigh_op_rgt_2')
// (17, 19, 'neigh_op_bnr_2')
// (18, 17, 'neigh_op_top_2')
// (18, 18, 'local_g0_2')
// (18, 18, 'lutff_2/out')
// (18, 18, 'lutff_global/cen')
// (18, 19, 'neigh_op_bot_2')
// (19, 17, 'neigh_op_tnl_2')
// (19, 18, 'neigh_op_lft_2')
// (19, 19, 'neigh_op_bnl_2')

wire n2564;
// (17, 17, 'neigh_op_tnr_6')
// (17, 18, 'neigh_op_rgt_6')
// (17, 19, 'neigh_op_bnr_6')
// (18, 17, 'local_g0_6')
// (18, 17, 'lutff_6/in_0')
// (18, 17, 'neigh_op_top_6')
// (18, 18, 'lutff_6/out')
// (18, 19, 'neigh_op_bot_6')
// (19, 17, 'neigh_op_tnl_6')
// (19, 18, 'neigh_op_lft_6')
// (19, 19, 'neigh_op_bnl_6')

wire n2565;
// (17, 17, 'neigh_op_tnr_7')
// (17, 18, 'neigh_op_rgt_7')
// (17, 18, 'sp4_h_r_3')
// (17, 19, 'neigh_op_bnr_7')
// (18, 17, 'neigh_op_top_7')
// (18, 18, 'lutff_7/out')
// (18, 18, 'sp4_h_r_14')
// (18, 19, 'neigh_op_bot_7')
// (19, 17, 'neigh_op_tnl_7')
// (19, 18, 'neigh_op_lft_7')
// (19, 18, 'sp4_h_r_27')
// (19, 19, 'neigh_op_bnl_7')
// (20, 18, 'local_g3_6')
// (20, 18, 'lutff_7/in_0')
// (20, 18, 'sp4_h_r_38')
// (21, 18, 'sp4_h_l_38')

wire n2566;
// (17, 17, 'sp4_h_r_11')
// (17, 17, 'sp4_h_r_7')
// (18, 17, 'sp4_h_r_18')
// (18, 17, 'sp4_h_r_22')
// (19, 16, 'neigh_op_tnr_7')
// (19, 17, 'neigh_op_rgt_7')
// (19, 17, 'sp4_h_r_31')
// (19, 17, 'sp4_h_r_35')
// (19, 18, 'neigh_op_bnr_7')
// (20, 16, 'neigh_op_top_7')
// (20, 17, 'local_g2_2')
// (20, 17, 'lutff_7/out')
// (20, 17, 'lutff_global/cen')
// (20, 17, 'sp4_h_r_42')
// (20, 17, 'sp4_h_r_46')
// (20, 18, 'neigh_op_bot_7')
// (21, 16, 'neigh_op_tnl_7')
// (21, 17, 'neigh_op_lft_7')
// (21, 17, 'sp4_h_l_42')
// (21, 17, 'sp4_h_l_46')
// (21, 17, 'sp4_h_r_7')
// (21, 18, 'neigh_op_bnl_7')
// (22, 17, 'sp4_h_r_18')
// (23, 17, 'sp4_h_r_31')
// (24, 17, 'sp4_h_r_42')
// (25, 17, 'sp4_h_l_42')

reg n2567 = 0;
// (17, 17, 'sp4_r_v_b_43')
// (17, 18, 'sp4_r_v_b_30')
// (17, 19, 'sp4_r_v_b_19')
// (17, 20, 'sp4_r_v_b_6')
// (17, 21, 'sp4_r_v_b_43')
// (17, 22, 'sp4_r_v_b_30')
// (17, 23, 'neigh_op_tnr_3')
// (17, 23, 'sp4_r_v_b_19')
// (17, 24, 'neigh_op_rgt_3')
// (17, 24, 'sp4_r_v_b_6')
// (17, 25, 'neigh_op_bnr_3')
// (18, 16, 'sp4_v_t_43')
// (18, 17, 'sp4_v_b_43')
// (18, 18, 'local_g3_6')
// (18, 18, 'lutff_1/in_0')
// (18, 18, 'sp4_v_b_30')
// (18, 19, 'sp4_v_b_19')
// (18, 20, 'sp4_v_b_6')
// (18, 20, 'sp4_v_t_43')
// (18, 21, 'sp4_v_b_43')
// (18, 22, 'sp4_v_b_30')
// (18, 23, 'neigh_op_top_3')
// (18, 23, 'sp4_v_b_19')
// (18, 24, 'lutff_3/out')
// (18, 24, 'sp4_v_b_6')
// (18, 25, 'neigh_op_bot_3')
// (19, 23, 'neigh_op_tnl_3')
// (19, 24, 'neigh_op_lft_3')
// (19, 25, 'neigh_op_bnl_3')

wire n2568;
// (17, 17, 'sp4_r_v_b_44')
// (17, 18, 'neigh_op_tnr_2')
// (17, 18, 'sp4_r_v_b_33')
// (17, 19, 'neigh_op_rgt_2')
// (17, 19, 'sp4_r_v_b_20')
// (17, 20, 'neigh_op_bnr_2')
// (17, 20, 'sp4_r_v_b_9')
// (18, 16, 'sp4_h_r_2')
// (18, 16, 'sp4_v_t_44')
// (18, 17, 'sp4_v_b_44')
// (18, 18, 'neigh_op_top_2')
// (18, 18, 'sp4_v_b_33')
// (18, 19, 'lutff_2/out')
// (18, 19, 'sp4_v_b_20')
// (18, 20, 'neigh_op_bot_2')
// (18, 20, 'sp4_v_b_9')
// (19, 16, 'sp4_h_r_15')
// (19, 18, 'neigh_op_tnl_2')
// (19, 19, 'neigh_op_lft_2')
// (19, 20, 'neigh_op_bnl_2')
// (20, 16, 'local_g2_2')
// (20, 16, 'lutff_global/cen')
// (20, 16, 'sp4_h_r_26')
// (21, 16, 'sp4_h_r_39')
// (22, 16, 'sp4_h_l_39')

wire n2569;
// (17, 18, 'lutff_1/cout')
// (17, 18, 'lutff_2/in_3')

wire n2570;
// (17, 18, 'lutff_2/cout')
// (17, 18, 'lutff_3/in_3')

wire n2571;
// (17, 18, 'lutff_3/cout')
// (17, 18, 'lutff_4/in_3')

wire n2572;
// (17, 18, 'lutff_4/cout')
// (17, 18, 'lutff_5/in_3')

reg n2573 = 0;
// (17, 18, 'neigh_op_tnr_0')
// (17, 19, 'neigh_op_rgt_0')
// (17, 20, 'neigh_op_bnr_0')
// (18, 18, 'local_g0_0')
// (18, 18, 'lutff_6/in_2')
// (18, 18, 'neigh_op_top_0')
// (18, 19, 'lutff_0/out')
// (18, 20, 'neigh_op_bot_0')
// (19, 18, 'neigh_op_tnl_0')
// (19, 19, 'neigh_op_lft_0')
// (19, 20, 'neigh_op_bnl_0')

wire n2574;
// (17, 18, 'neigh_op_tnr_5')
// (17, 19, 'neigh_op_rgt_5')
// (17, 20, 'neigh_op_bnr_5')
// (18, 18, 'local_g1_5')
// (18, 18, 'lutff_7/in_3')
// (18, 18, 'neigh_op_top_5')
// (18, 19, 'lutff_5/out')
// (18, 20, 'neigh_op_bot_5')
// (19, 18, 'neigh_op_tnl_5')
// (19, 19, 'neigh_op_lft_5')
// (19, 20, 'neigh_op_bnl_5')

wire n2575;
// (17, 18, 'neigh_op_tnr_7')
// (17, 19, 'neigh_op_rgt_7')
// (17, 19, 'sp4_h_r_3')
// (17, 19, 'sp4_h_r_7')
// (17, 20, 'neigh_op_bnr_7')
// (18, 18, 'neigh_op_top_7')
// (18, 19, 'local_g0_2')
// (18, 19, 'lutff_7/out')
// (18, 19, 'lutff_global/cen')
// (18, 19, 'sp4_h_r_14')
// (18, 19, 'sp4_h_r_18')
// (18, 20, 'neigh_op_bot_7')
// (19, 18, 'neigh_op_tnl_7')
// (19, 19, 'neigh_op_lft_7')
// (19, 19, 'sp4_h_r_27')
// (19, 19, 'sp4_h_r_31')
// (19, 20, 'neigh_op_bnl_7')
// (20, 19, 'sp4_h_r_38')
// (20, 19, 'sp4_h_r_42')
// (21, 19, 'sp4_h_l_38')
// (21, 19, 'sp4_h_l_42')
// (21, 19, 'sp4_h_r_11')
// (22, 19, 'sp4_h_r_22')
// (23, 19, 'sp4_h_r_35')
// (24, 19, 'sp4_h_r_46')
// (25, 19, 'sp4_h_l_46')

reg n2576 = 0;
// (17, 18, 'sp4_h_r_1')
// (18, 18, 'local_g1_4')
// (18, 18, 'lutff_6/in_3')
// (18, 18, 'sp4_h_r_12')
// (19, 17, 'neigh_op_tnr_2')
// (19, 18, 'neigh_op_rgt_2')
// (19, 18, 'sp4_h_r_25')
// (19, 19, 'neigh_op_bnr_2')
// (20, 17, 'neigh_op_top_2')
// (20, 18, 'lutff_2/out')
// (20, 18, 'sp4_h_r_36')
// (20, 19, 'neigh_op_bot_2')
// (21, 17, 'neigh_op_tnl_2')
// (21, 18, 'neigh_op_lft_2')
// (21, 18, 'sp4_h_l_36')
// (21, 19, 'neigh_op_bnl_2')

wire n2577;
// (17, 19, 'lutff_1/cout')
// (17, 19, 'lutff_2/in_3')

wire n2578;
// (17, 19, 'lutff_3/cout')
// (17, 19, 'lutff_4/in_3')

wire n2579;
// (17, 19, 'lutff_5/cout')
// (17, 19, 'lutff_6/in_3')

wire n2580;
// (17, 19, 'lutff_7/cout')
// (17, 20, 'carry_in')
// (17, 20, 'carry_in_mux')
// (17, 20, 'lutff_0/in_3')

reg n2581 = 0;
// (17, 19, 'neigh_op_tnr_3')
// (17, 20, 'neigh_op_rgt_3')
// (17, 20, 'sp4_h_r_11')
// (17, 21, 'neigh_op_bnr_3')
// (18, 19, 'neigh_op_top_3')
// (18, 20, 'lutff_3/out')
// (18, 20, 'sp4_h_r_22')
// (18, 21, 'neigh_op_bot_3')
// (19, 19, 'neigh_op_tnl_3')
// (19, 20, 'neigh_op_lft_3')
// (19, 20, 'sp4_h_r_35')
// (19, 21, 'neigh_op_bnl_3')
// (20, 17, 'sp4_r_v_b_46')
// (20, 18, 'local_g2_3')
// (20, 18, 'lutff_3/in_2')
// (20, 18, 'sp4_r_v_b_35')
// (20, 19, 'sp4_r_v_b_22')
// (20, 20, 'sp4_h_r_46')
// (20, 20, 'sp4_r_v_b_11')
// (21, 16, 'sp4_v_t_46')
// (21, 17, 'sp4_v_b_46')
// (21, 18, 'sp4_v_b_35')
// (21, 19, 'sp4_v_b_22')
// (21, 20, 'sp4_h_l_46')
// (21, 20, 'sp4_v_b_11')

wire n2582;
// (17, 19, 'sp4_r_v_b_45')
// (17, 20, 'sp4_r_v_b_32')
// (17, 21, 'neigh_op_tnr_4')
// (17, 21, 'sp4_r_v_b_21')
// (17, 22, 'neigh_op_rgt_4')
// (17, 22, 'sp4_r_v_b_8')
// (17, 23, 'neigh_op_bnr_4')
// (18, 18, 'sp4_v_t_45')
// (18, 19, 'sp4_v_b_45')
// (18, 20, 'sp4_v_b_32')
// (18, 21, 'neigh_op_top_4')
// (18, 21, 'sp4_v_b_21')
// (18, 22, 'local_g0_2')
// (18, 22, 'lutff_4/out')
// (18, 22, 'lutff_global/cen')
// (18, 22, 'sp4_h_r_2')
// (18, 22, 'sp4_v_b_8')
// (18, 23, 'neigh_op_bot_4')
// (19, 21, 'neigh_op_tnl_4')
// (19, 22, 'neigh_op_lft_4')
// (19, 22, 'sp4_h_r_15')
// (19, 23, 'neigh_op_bnl_4')
// (20, 22, 'sp4_h_r_26')
// (21, 22, 'sp4_h_r_39')
// (22, 22, 'sp4_h_l_39')

wire n2583;
// (17, 20, 'neigh_op_tnr_1')
// (17, 21, 'neigh_op_rgt_1')
// (17, 21, 'sp4_h_r_7')
// (17, 22, 'neigh_op_bnr_1')
// (18, 20, 'neigh_op_top_1')
// (18, 21, 'lutff_1/out')
// (18, 21, 'sp4_h_r_18')
// (18, 22, 'neigh_op_bot_1')
// (19, 20, 'neigh_op_tnl_1')
// (19, 21, 'neigh_op_lft_1')
// (19, 21, 'sp4_h_r_31')
// (19, 22, 'neigh_op_bnl_1')
// (20, 18, 'sp4_r_v_b_36')
// (20, 19, 'sp4_r_v_b_25')
// (20, 20, 'local_g2_4')
// (20, 20, 'lutff_3/in_1')
// (20, 20, 'sp4_r_v_b_12')
// (20, 21, 'sp4_h_r_42')
// (20, 21, 'sp4_r_v_b_1')
// (21, 17, 'sp4_v_t_36')
// (21, 18, 'sp4_v_b_36')
// (21, 19, 'sp4_v_b_25')
// (21, 20, 'sp4_v_b_12')
// (21, 21, 'sp4_h_l_42')
// (21, 21, 'sp4_v_b_1')

wire n2584;
// (17, 20, 'neigh_op_tnr_2')
// (17, 21, 'neigh_op_rgt_2')
// (17, 22, 'neigh_op_bnr_2')
// (18, 20, 'neigh_op_top_2')
// (18, 21, 'local_g2_2')
// (18, 21, 'lutff_2/out')
// (18, 21, 'lutff_global/cen')
// (18, 22, 'neigh_op_bot_2')
// (19, 20, 'neigh_op_tnl_2')
// (19, 21, 'neigh_op_lft_2')
// (19, 22, 'neigh_op_bnl_2')

reg n2585 = 0;
// (17, 20, 'neigh_op_tnr_7')
// (17, 21, 'neigh_op_rgt_7')
// (17, 22, 'neigh_op_bnr_7')
// (18, 20, 'neigh_op_top_7')
// (18, 21, 'local_g2_7')
// (18, 21, 'lutff_1/in_0')
// (18, 21, 'lutff_7/out')
// (18, 22, 'neigh_op_bot_7')
// (19, 20, 'neigh_op_tnl_7')
// (19, 21, 'neigh_op_lft_7')
// (19, 22, 'neigh_op_bnl_7')

reg n2586 = 0;
// (17, 20, 'sp4_r_v_b_40')
// (17, 21, 'sp4_r_v_b_29')
// (17, 22, 'sp4_r_v_b_16')
// (17, 23, 'sp4_r_v_b_5')
// (18, 19, 'sp4_v_t_40')
// (18, 20, 'sp4_v_b_40')
// (18, 21, 'sp4_v_b_29')
// (18, 22, 'local_g1_0')
// (18, 22, 'lutff_1/in_0')
// (18, 22, 'sp4_v_b_16')
// (18, 23, 'sp4_h_r_0')
// (18, 23, 'sp4_v_b_5')
// (19, 22, 'neigh_op_tnr_4')
// (19, 23, 'neigh_op_rgt_4')
// (19, 23, 'sp4_h_r_13')
// (19, 24, 'neigh_op_bnr_4')
// (20, 22, 'neigh_op_top_4')
// (20, 23, 'lutff_4/out')
// (20, 23, 'sp4_h_r_24')
// (20, 24, 'neigh_op_bot_4')
// (21, 22, 'neigh_op_tnl_4')
// (21, 23, 'neigh_op_lft_4')
// (21, 23, 'sp4_h_r_37')
// (21, 24, 'neigh_op_bnl_4')
// (22, 23, 'sp4_h_l_37')

wire n2587;
// (17, 21, 'neigh_op_tnr_1')
// (17, 22, 'neigh_op_rgt_1')
// (17, 23, 'neigh_op_bnr_1')
// (18, 21, 'local_g0_1')
// (18, 21, 'lutff_1/in_2')
// (18, 21, 'neigh_op_top_1')
// (18, 22, 'lutff_1/out')
// (18, 23, 'neigh_op_bot_1')
// (19, 21, 'neigh_op_tnl_1')
// (19, 22, 'neigh_op_lft_1')
// (19, 23, 'neigh_op_bnl_1')

wire n2588;
// (17, 21, 'neigh_op_tnr_2')
// (17, 22, 'neigh_op_rgt_2')
// (17, 23, 'neigh_op_bnr_2')
// (18, 19, 'sp4_r_v_b_40')
// (18, 20, 'sp4_r_v_b_29')
// (18, 21, 'neigh_op_top_2')
// (18, 21, 'sp4_r_v_b_16')
// (18, 22, 'lutff_2/out')
// (18, 22, 'sp4_r_v_b_5')
// (18, 23, 'neigh_op_bot_2')
// (19, 18, 'sp4_h_r_5')
// (19, 18, 'sp4_v_t_40')
// (19, 19, 'sp4_v_b_40')
// (19, 20, 'sp4_v_b_29')
// (19, 21, 'neigh_op_tnl_2')
// (19, 21, 'sp4_v_b_16')
// (19, 22, 'neigh_op_lft_2')
// (19, 22, 'sp4_v_b_5')
// (19, 23, 'neigh_op_bnl_2')
// (20, 18, 'local_g1_0')
// (20, 18, 'lutff_7/in_2')
// (20, 18, 'sp4_h_r_16')
// (21, 18, 'sp4_h_r_29')
// (22, 18, 'sp4_h_r_40')
// (23, 18, 'sp4_h_l_40')

reg n2589 = 0;
// (17, 21, 'neigh_op_tnr_3')
// (17, 22, 'neigh_op_rgt_3')
// (17, 23, 'neigh_op_bnr_3')
// (18, 15, 'sp4_r_v_b_38')
// (18, 16, 'sp4_r_v_b_27')
// (18, 17, 'local_g2_6')
// (18, 17, 'lutff_2/in_2')
// (18, 17, 'sp4_r_v_b_14')
// (18, 18, 'sp4_r_v_b_3')
// (18, 19, 'sp4_r_v_b_42')
// (18, 20, 'sp4_r_v_b_31')
// (18, 21, 'neigh_op_top_3')
// (18, 21, 'sp4_r_v_b_18')
// (18, 22, 'lutff_3/out')
// (18, 22, 'sp4_r_v_b_7')
// (18, 23, 'neigh_op_bot_3')
// (19, 14, 'sp4_v_t_38')
// (19, 15, 'sp4_v_b_38')
// (19, 16, 'sp4_v_b_27')
// (19, 17, 'sp4_v_b_14')
// (19, 18, 'sp4_v_b_3')
// (19, 18, 'sp4_v_t_42')
// (19, 19, 'sp4_v_b_42')
// (19, 20, 'sp4_v_b_31')
// (19, 21, 'neigh_op_tnl_3')
// (19, 21, 'sp4_v_b_18')
// (19, 22, 'neigh_op_lft_3')
// (19, 22, 'sp4_v_b_7')
// (19, 23, 'neigh_op_bnl_3')

wire n2590;
// (17, 21, 'sp4_h_r_9')
// (18, 21, 'sp4_h_r_20')
// (19, 20, 'neigh_op_tnr_6')
// (19, 21, 'neigh_op_rgt_6')
// (19, 21, 'sp4_h_r_33')
// (19, 22, 'neigh_op_bnr_6')
// (20, 18, 'sp4_r_v_b_38')
// (20, 19, 'sp4_r_v_b_27')
// (20, 20, 'neigh_op_top_6')
// (20, 20, 'sp4_r_v_b_14')
// (20, 21, 'local_g1_3')
// (20, 21, 'lutff_6/out')
// (20, 21, 'lutff_global/cen')
// (20, 21, 'sp4_h_r_44')
// (20, 21, 'sp4_r_v_b_3')
// (20, 22, 'neigh_op_bot_6')
// (21, 17, 'sp4_v_t_38')
// (21, 18, 'sp4_v_b_38')
// (21, 19, 'sp4_v_b_27')
// (21, 20, 'neigh_op_tnl_6')
// (21, 20, 'sp4_v_b_14')
// (21, 21, 'neigh_op_lft_6')
// (21, 21, 'sp4_h_l_44')
// (21, 21, 'sp4_v_b_3')
// (21, 22, 'neigh_op_bnl_6')

wire n2591;
// (17, 21, 'sp4_r_v_b_45')
// (17, 22, 'sp4_r_v_b_32')
// (17, 23, 'neigh_op_tnr_4')
// (17, 23, 'sp4_r_v_b_21')
// (17, 24, 'neigh_op_rgt_4')
// (17, 24, 'sp4_r_v_b_8')
// (17, 25, 'neigh_op_bnr_4')
// (18, 20, 'sp4_v_t_45')
// (18, 21, 'sp4_v_b_45')
// (18, 22, 'sp4_v_b_32')
// (18, 23, 'neigh_op_top_4')
// (18, 23, 'sp4_v_b_21')
// (18, 24, 'local_g0_2')
// (18, 24, 'lutff_4/out')
// (18, 24, 'lutff_global/cen')
// (18, 24, 'sp4_h_r_2')
// (18, 24, 'sp4_v_b_8')
// (18, 25, 'neigh_op_bot_4')
// (19, 23, 'neigh_op_tnl_4')
// (19, 24, 'neigh_op_lft_4')
// (19, 24, 'sp4_h_r_15')
// (19, 25, 'neigh_op_bnl_4')
// (20, 24, 'sp4_h_r_26')
// (21, 24, 'sp4_h_r_39')
// (22, 24, 'sp4_h_l_39')

reg n2592 = 0;
// (17, 22, 'neigh_op_tnr_1')
// (17, 23, 'neigh_op_rgt_1')
// (17, 24, 'neigh_op_bnr_1')
// (18, 22, 'local_g0_1')
// (18, 22, 'lutff_2/in_1')
// (18, 22, 'neigh_op_top_1')
// (18, 23, 'lutff_1/out')
// (18, 24, 'neigh_op_bot_1')
// (19, 22, 'neigh_op_tnl_1')
// (19, 23, 'neigh_op_lft_1')
// (19, 24, 'neigh_op_bnl_1')

wire n2593;
// (17, 22, 'sp4_h_r_6')
// (18, 22, 'sp4_h_r_19')
// (19, 22, 'sp4_h_r_30')
// (20, 22, 'sp4_h_r_43')
// (21, 21, 'neigh_op_tnr_7')
// (21, 22, 'neigh_op_rgt_7')
// (21, 22, 'sp4_h_l_43')
// (21, 22, 'sp4_h_r_3')
// (21, 22, 'sp4_h_r_6')
// (21, 23, 'neigh_op_bnr_7')
// (22, 21, 'neigh_op_top_7')
// (22, 22, 'local_g1_3')
// (22, 22, 'lutff_7/out')
// (22, 22, 'lutff_global/cen')
// (22, 22, 'sp4_h_r_14')
// (22, 22, 'sp4_h_r_19')
// (22, 23, 'neigh_op_bot_7')
// (23, 21, 'neigh_op_tnl_7')
// (23, 22, 'neigh_op_lft_7')
// (23, 22, 'sp4_h_r_27')
// (23, 22, 'sp4_h_r_30')
// (23, 23, 'neigh_op_bnl_7')
// (24, 22, 'sp4_h_r_38')
// (24, 22, 'sp4_h_r_43')
// (25, 22, 'sp4_h_l_38')
// (25, 22, 'sp4_h_l_43')

wire n2594;
// (17, 23, 'sp4_r_v_b_43')
// (17, 24, 'sp4_r_v_b_30')
// (17, 25, 'sp4_r_v_b_19')
// (17, 26, 'sp4_r_v_b_6')
// (18, 22, 'sp4_h_r_0')
// (18, 22, 'sp4_v_t_43')
// (18, 23, 'local_g3_3')
// (18, 23, 'lutff_global/cen')
// (18, 23, 'sp4_v_b_43')
// (18, 24, 'sp4_v_b_30')
// (18, 25, 'sp4_v_b_19')
// (18, 26, 'sp4_v_b_6')
// (19, 21, 'neigh_op_tnr_4')
// (19, 22, 'neigh_op_rgt_4')
// (19, 22, 'sp4_h_r_13')
// (19, 23, 'neigh_op_bnr_4')
// (20, 21, 'neigh_op_top_4')
// (20, 22, 'lutff_4/out')
// (20, 22, 'sp4_h_r_24')
// (20, 23, 'neigh_op_bot_4')
// (21, 21, 'neigh_op_tnl_4')
// (21, 22, 'neigh_op_lft_4')
// (21, 22, 'sp4_h_r_37')
// (21, 23, 'neigh_op_bnl_4')
// (22, 22, 'sp4_h_l_37')

reg n2595 = 0;
// (18, 1, 'local_g0_0')
// (18, 1, 'lutff_1/in_1')
// (18, 1, 'sp4_h_r_0')
// (19, 0, 'logic_op_tnr_4')
// (19, 1, 'neigh_op_rgt_4')
// (19, 1, 'sp4_h_r_13')
// (19, 2, 'neigh_op_bnr_4')
// (20, 0, 'logic_op_top_4')
// (20, 1, 'local_g3_4')
// (20, 1, 'lutff_1/in_2')
// (20, 1, 'lutff_4/in_1')
// (20, 1, 'lutff_4/out')
// (20, 1, 'sp4_h_r_24')
// (20, 2, 'neigh_op_bot_4')
// (21, 0, 'logic_op_tnl_4')
// (21, 1, 'local_g0_4')
// (21, 1, 'lutff_0/in_0')
// (21, 1, 'lutff_5/in_1')
// (21, 1, 'neigh_op_lft_4')
// (21, 1, 'sp4_h_r_37')
// (21, 2, 'neigh_op_bnl_4')
// (22, 1, 'sp4_h_l_37')

wire n2596;
// (18, 1, 'lutff_1/cout')
// (18, 1, 'lutff_2/in_3')

wire n2597;
// (18, 1, 'lutff_2/cout')
// (18, 1, 'lutff_3/in_3')

wire n2598;
// (18, 1, 'lutff_3/cout')
// (18, 1, 'lutff_4/in_3')

wire n2599;
// (18, 1, 'lutff_4/cout')
// (18, 1, 'lutff_5/in_3')

wire n2600;
// (18, 1, 'sp4_h_r_10')
// (19, 1, 'sp4_h_r_23')
// (20, 1, 'local_g2_2')
// (20, 1, 'lutff_global/cen')
// (20, 1, 'neigh_op_tnr_4')
// (20, 1, 'sp4_h_r_34')
// (20, 2, 'neigh_op_rgt_4')
// (20, 3, 'neigh_op_bnr_4')
// (21, 0, 'span12_vert_11')
// (21, 1, 'local_g3_3')
// (21, 1, 'lutff_global/cen')
// (21, 1, 'neigh_op_top_4')
// (21, 1, 'sp12_v_b_11')
// (21, 1, 'sp4_h_r_47')
// (21, 2, 'lutff_4/out')
// (21, 2, 'sp12_v_b_8')
// (21, 2, 'sp4_r_v_b_41')
// (21, 3, 'neigh_op_bot_4')
// (21, 3, 'sp12_v_b_7')
// (21, 3, 'sp4_r_v_b_28')
// (21, 4, 'sp12_v_b_4')
// (21, 4, 'sp4_r_v_b_17')
// (21, 5, 'sp12_v_b_3')
// (21, 5, 'sp4_r_v_b_4')
// (21, 6, 'sp12_v_b_0')
// (22, 1, 'neigh_op_tnl_4')
// (22, 1, 'sp4_h_l_47')
// (22, 1, 'sp4_v_t_41')
// (22, 2, 'neigh_op_lft_4')
// (22, 2, 'sp4_v_b_41')
// (22, 3, 'neigh_op_bnl_4')
// (22, 3, 'sp4_v_b_28')
// (22, 4, 'sp4_v_b_17')
// (22, 5, 'sp4_v_b_4')

reg n2601 = 0;
// (18, 3, 'local_g1_6')
// (18, 3, 'lutff_1/in_0')
// (18, 3, 'sp4_h_r_6')
// (19, 3, 'sp4_h_r_19')
// (20, 3, 'local_g2_7')
// (20, 3, 'lutff_2/in_1')
// (20, 3, 'sp4_h_r_30')
// (20, 3, 'sp4_r_v_b_39')
// (20, 4, 'sp4_r_v_b_26')
// (20, 5, 'neigh_op_tnr_1')
// (20, 5, 'sp4_r_v_b_15')
// (20, 6, 'neigh_op_rgt_1')
// (20, 6, 'sp4_r_v_b_2')
// (20, 7, 'neigh_op_bnr_1')
// (21, 2, 'sp4_v_t_39')
// (21, 3, 'sp4_h_r_43')
// (21, 3, 'sp4_v_b_39')
// (21, 4, 'sp4_r_v_b_43')
// (21, 4, 'sp4_v_b_26')
// (21, 5, 'neigh_op_top_1')
// (21, 5, 'sp4_r_v_b_30')
// (21, 5, 'sp4_v_b_15')
// (21, 6, 'lutff_1/out')
// (21, 6, 'sp4_r_v_b_19')
// (21, 6, 'sp4_v_b_2')
// (21, 7, 'neigh_op_bot_1')
// (21, 7, 'sp4_r_v_b_6')
// (22, 3, 'sp4_h_l_43')
// (22, 3, 'sp4_v_t_43')
// (22, 4, 'sp4_v_b_43')
// (22, 5, 'neigh_op_tnl_1')
// (22, 5, 'sp4_v_b_30')
// (22, 6, 'neigh_op_lft_1')
// (22, 6, 'sp4_v_b_19')
// (22, 7, 'neigh_op_bnl_1')
// (22, 7, 'sp4_v_b_6')

wire n2602;
// (18, 3, 'sp4_r_v_b_38')
// (18, 4, 'sp4_r_v_b_27')
// (18, 5, 'sp4_r_v_b_14')
// (18, 6, 'local_g1_3')
// (18, 6, 'lutff_global/cen')
// (18, 6, 'sp4_r_v_b_3')
// (19, 2, 'sp4_v_t_38')
// (19, 3, 'sp4_v_b_38')
// (19, 4, 'sp4_v_b_27')
// (19, 5, 'neigh_op_tnr_7')
// (19, 5, 'sp4_r_v_b_43')
// (19, 5, 'sp4_v_b_14')
// (19, 6, 'neigh_op_rgt_7')
// (19, 6, 'sp4_h_r_3')
// (19, 6, 'sp4_r_v_b_30')
// (19, 6, 'sp4_v_b_3')
// (19, 7, 'neigh_op_bnr_7')
// (19, 7, 'sp4_r_v_b_19')
// (19, 8, 'sp4_r_v_b_6')
// (20, 4, 'local_g1_3')
// (20, 4, 'lutff_global/cen')
// (20, 4, 'sp4_h_r_11')
// (20, 4, 'sp4_v_t_43')
// (20, 5, 'neigh_op_top_7')
// (20, 5, 'sp4_v_b_43')
// (20, 6, 'lutff_7/out')
// (20, 6, 'sp4_h_r_14')
// (20, 6, 'sp4_v_b_30')
// (20, 7, 'neigh_op_bot_7')
// (20, 7, 'sp4_v_b_19')
// (20, 8, 'sp4_v_b_6')
// (21, 4, 'sp4_h_r_22')
// (21, 5, 'neigh_op_tnl_7')
// (21, 6, 'neigh_op_lft_7')
// (21, 6, 'sp4_h_r_27')
// (21, 7, 'neigh_op_bnl_7')
// (22, 4, 'sp4_h_r_35')
// (22, 6, 'sp4_h_r_38')
// (23, 4, 'sp4_h_r_46')
// (23, 6, 'sp4_h_l_38')
// (24, 4, 'sp4_h_l_46')

wire n2603;
// (18, 4, 'local_g0_2')
// (18, 4, 'lutff_global/cen')
// (18, 4, 'sp4_h_r_2')
// (19, 3, 'neigh_op_tnr_5')
// (19, 4, 'neigh_op_rgt_5')
// (19, 4, 'sp4_h_r_15')
// (19, 5, 'neigh_op_bnr_5')
// (20, 3, 'neigh_op_top_5')
// (20, 4, 'lutff_5/out')
// (20, 4, 'sp4_h_r_26')
// (20, 5, 'neigh_op_bot_5')
// (21, 3, 'neigh_op_tnl_5')
// (21, 4, 'neigh_op_lft_5')
// (21, 4, 'sp4_h_r_39')
// (21, 5, 'neigh_op_bnl_5')
// (22, 4, 'sp4_h_l_39')

wire n2604;
// (18, 5, 'neigh_op_tnr_0')
// (18, 6, 'neigh_op_rgt_0')
// (18, 7, 'neigh_op_bnr_0')
// (19, 5, 'neigh_op_top_0')
// (19, 6, 'ram/RDATA_7')
// (19, 6, 'sp4_h_r_0')
// (19, 7, 'neigh_op_bot_0')
// (20, 5, 'neigh_op_tnl_0')
// (20, 6, 'neigh_op_lft_0')
// (20, 6, 'sp4_h_r_13')
// (20, 7, 'neigh_op_bnl_0')
// (21, 6, 'local_g3_0')
// (21, 6, 'lutff_3/in_0')
// (21, 6, 'sp4_h_r_24')
// (22, 6, 'sp4_h_r_37')
// (23, 6, 'sp4_h_l_37')

wire n2605;
// (18, 5, 'neigh_op_tnr_1')
// (18, 6, 'neigh_op_rgt_1')
// (18, 7, 'neigh_op_bnr_1')
// (19, 3, 'sp4_r_v_b_38')
// (19, 4, 'sp4_r_v_b_27')
// (19, 5, 'neigh_op_top_1')
// (19, 5, 'sp4_r_v_b_14')
// (19, 6, 'ram/RDATA_6')
// (19, 6, 'sp4_r_v_b_3')
// (19, 7, 'neigh_op_bot_1')
// (20, 2, 'sp4_v_t_38')
// (20, 3, 'sp4_v_b_38')
// (20, 4, 'sp4_v_b_27')
// (20, 5, 'neigh_op_tnl_1')
// (20, 5, 'sp4_v_b_14')
// (20, 6, 'neigh_op_lft_1')
// (20, 6, 'sp4_h_r_9')
// (20, 6, 'sp4_v_b_3')
// (20, 7, 'neigh_op_bnl_1')
// (21, 6, 'local_g0_4')
// (21, 6, 'lutff_6/in_0')
// (21, 6, 'sp4_h_r_20')
// (22, 6, 'sp4_h_r_33')
// (23, 6, 'sp4_h_r_44')
// (24, 6, 'sp4_h_l_44')

wire n2606;
// (18, 5, 'neigh_op_tnr_2')
// (18, 6, 'neigh_op_rgt_2')
// (18, 7, 'neigh_op_bnr_2')
// (19, 5, 'neigh_op_top_2')
// (19, 6, 'ram/RDATA_5')
// (19, 6, 'sp4_h_r_4')
// (19, 7, 'neigh_op_bot_2')
// (20, 5, 'neigh_op_tnl_2')
// (20, 6, 'neigh_op_lft_2')
// (20, 6, 'sp4_h_r_17')
// (20, 7, 'neigh_op_bnl_2')
// (21, 6, 'local_g2_4')
// (21, 6, 'lutff_1/in_3')
// (21, 6, 'sp4_h_r_28')
// (22, 6, 'sp4_h_r_41')
// (23, 6, 'sp4_h_l_41')

wire n2607;
// (18, 5, 'neigh_op_tnr_3')
// (18, 6, 'neigh_op_rgt_3')
// (18, 6, 'sp4_h_r_11')
// (18, 7, 'neigh_op_bnr_3')
// (19, 5, 'neigh_op_top_3')
// (19, 6, 'ram/RDATA_4')
// (19, 6, 'sp4_h_r_22')
// (19, 7, 'neigh_op_bot_3')
// (20, 5, 'neigh_op_tnl_3')
// (20, 6, 'neigh_op_lft_3')
// (20, 6, 'sp4_h_r_35')
// (20, 7, 'neigh_op_bnl_3')
// (21, 6, 'local_g2_6')
// (21, 6, 'lutff_4/in_2')
// (21, 6, 'sp4_h_r_46')
// (22, 6, 'sp4_h_l_46')

wire n2608;
// (18, 5, 'neigh_op_tnr_4')
// (18, 6, 'neigh_op_rgt_4')
// (18, 7, 'neigh_op_bnr_4')
// (19, 3, 'sp4_r_v_b_44')
// (19, 4, 'sp4_r_v_b_33')
// (19, 5, 'neigh_op_top_4')
// (19, 5, 'sp4_r_v_b_20')
// (19, 6, 'ram/RDATA_3')
// (19, 6, 'sp4_r_v_b_9')
// (19, 7, 'neigh_op_bot_4')
// (20, 2, 'sp4_v_t_44')
// (20, 3, 'sp4_v_b_44')
// (20, 4, 'sp4_v_b_33')
// (20, 5, 'neigh_op_tnl_4')
// (20, 5, 'sp4_v_b_20')
// (20, 6, 'neigh_op_lft_4')
// (20, 6, 'sp4_h_r_3')
// (20, 6, 'sp4_v_b_9')
// (20, 7, 'neigh_op_bnl_4')
// (21, 6, 'local_g1_6')
// (21, 6, 'lutff_0/in_3')
// (21, 6, 'sp4_h_r_14')
// (22, 6, 'sp4_h_r_27')
// (23, 6, 'sp4_h_r_38')
// (24, 6, 'sp4_h_l_38')

wire n2609;
// (18, 5, 'neigh_op_tnr_5')
// (18, 6, 'neigh_op_rgt_5')
// (18, 7, 'neigh_op_bnr_5')
// (19, 5, 'neigh_op_top_5')
// (19, 6, 'ram/RDATA_2')
// (19, 6, 'sp4_h_r_10')
// (19, 7, 'neigh_op_bot_5')
// (20, 5, 'neigh_op_tnl_5')
// (20, 6, 'neigh_op_lft_5')
// (20, 6, 'sp4_h_r_23')
// (20, 7, 'neigh_op_bnl_5')
// (21, 6, 'local_g3_2')
// (21, 6, 'lutff_2/in_1')
// (21, 6, 'sp4_h_r_34')
// (22, 6, 'sp4_h_r_47')
// (23, 6, 'sp4_h_l_47')

wire n2610;
// (18, 5, 'neigh_op_tnr_7')
// (18, 6, 'neigh_op_rgt_7')
// (18, 6, 'sp4_h_r_3')
// (18, 7, 'neigh_op_bnr_7')
// (19, 5, 'neigh_op_top_7')
// (19, 6, 'ram/RDATA_0')
// (19, 6, 'sp4_h_r_14')
// (19, 7, 'neigh_op_bot_7')
// (20, 5, 'neigh_op_tnl_7')
// (20, 6, 'neigh_op_lft_7')
// (20, 6, 'sp4_h_r_27')
// (20, 7, 'neigh_op_bnl_7')
// (21, 6, 'local_g3_6')
// (21, 6, 'lutff_7/in_0')
// (21, 6, 'sp4_h_r_38')
// (22, 6, 'sp4_h_l_38')

wire n2611;
// (18, 6, 'lutff_1/cout')
// (18, 6, 'lutff_2/in_3')

wire n2612;
// (18, 6, 'lutff_2/cout')
// (18, 6, 'lutff_3/in_3')

wire n2613;
// (18, 6, 'lutff_3/cout')
// (18, 6, 'lutff_4/in_3')

wire n2614;
// (18, 6, 'lutff_4/cout')
// (18, 6, 'lutff_5/in_3')

wire n2615;
// (18, 6, 'lutff_5/cout')
// (18, 6, 'lutff_6/in_3')

wire n2616;
// (18, 6, 'sp4_r_v_b_38')
// (18, 7, 'neigh_op_tnr_7')
// (18, 7, 'sp4_r_v_b_27')
// (18, 8, 'neigh_op_rgt_7')
// (18, 8, 'sp4_r_v_b_14')
// (18, 9, 'neigh_op_bnr_7')
// (18, 9, 'sp4_r_v_b_3')
// (19, 5, 'sp4_v_t_38')
// (19, 6, 'sp4_v_b_38')
// (19, 7, 'neigh_op_top_7')
// (19, 7, 'sp4_v_b_27')
// (19, 8, 'ram/RDATA_0')
// (19, 8, 'sp4_v_b_14')
// (19, 9, 'neigh_op_bot_7')
// (19, 9, 'sp4_h_r_3')
// (19, 9, 'sp4_v_b_3')
// (20, 7, 'neigh_op_tnl_7')
// (20, 8, 'neigh_op_lft_7')
// (20, 9, 'neigh_op_bnl_7')
// (20, 9, 'sp4_h_r_14')
// (21, 9, 'sp4_h_r_27')
// (22, 9, 'local_g2_6')
// (22, 9, 'lutff_3/in_3')
// (22, 9, 'sp4_h_r_38')
// (23, 9, 'sp4_h_l_38')

reg n2617 = 0;
// (18, 6, 'sp4_r_v_b_42')
// (18, 7, 'sp4_r_v_b_31')
// (18, 8, 'sp4_r_v_b_18')
// (18, 9, 'sp4_r_v_b_7')
// (19, 5, 'sp4_h_r_7')
// (19, 5, 'sp4_v_t_42')
// (19, 6, 'local_g3_2')
// (19, 6, 'ram/WDATA_5')
// (19, 6, 'sp4_v_b_42')
// (19, 7, 'sp4_v_b_31')
// (19, 8, 'sp4_v_b_18')
// (19, 9, 'sp4_v_b_7')
// (20, 5, 'sp4_h_r_18')
// (21, 4, 'neigh_op_tnr_5')
// (21, 5, 'neigh_op_rgt_5')
// (21, 5, 'sp4_h_r_31')
// (21, 6, 'neigh_op_bnr_5')
// (22, 4, 'neigh_op_top_5')
// (22, 5, 'lutff_5/out')
// (22, 5, 'sp4_h_r_42')
// (22, 6, 'neigh_op_bot_5')
// (23, 4, 'neigh_op_tnl_5')
// (23, 5, 'neigh_op_lft_5')
// (23, 5, 'sp4_h_l_42')
// (23, 6, 'neigh_op_bnl_5')

wire n2618;
// (18, 7, 'neigh_op_tnr_4')
// (18, 8, 'neigh_op_rgt_4')
// (18, 9, 'neigh_op_bnr_4')
// (19, 7, 'neigh_op_top_4')
// (19, 8, 'ram/RDATA_3')
// (19, 8, 'sp4_h_r_8')
// (19, 9, 'neigh_op_bot_4')
// (20, 7, 'neigh_op_tnl_4')
// (20, 8, 'neigh_op_lft_4')
// (20, 8, 'sp4_h_r_21')
// (20, 9, 'neigh_op_bnl_4')
// (21, 8, 'sp4_h_r_32')
// (22, 8, 'sp4_h_r_45')
// (22, 9, 'local_g3_5')
// (22, 9, 'lutff_4/in_2')
// (22, 9, 'sp4_r_v_b_45')
// (22, 10, 'sp4_r_v_b_32')
// (22, 11, 'sp4_r_v_b_21')
// (22, 12, 'sp4_r_v_b_8')
// (23, 8, 'sp4_h_l_45')
// (23, 8, 'sp4_v_t_45')
// (23, 9, 'sp4_v_b_45')
// (23, 10, 'sp4_v_b_32')
// (23, 11, 'sp4_v_b_21')
// (23, 12, 'sp4_v_b_8')

wire n2619;
// (18, 7, 'neigh_op_tnr_5')
// (18, 8, 'neigh_op_rgt_5')
// (18, 9, 'neigh_op_bnr_5')
// (19, 7, 'neigh_op_top_5')
// (19, 8, 'ram/RDATA_2')
// (19, 8, 'sp4_h_r_10')
// (19, 9, 'neigh_op_bot_5')
// (20, 7, 'neigh_op_tnl_5')
// (20, 8, 'neigh_op_lft_5')
// (20, 8, 'sp4_h_r_23')
// (20, 9, 'neigh_op_bnl_5')
// (21, 8, 'sp4_h_r_34')
// (22, 8, 'sp4_h_r_47')
// (22, 9, 'local_g3_7')
// (22, 9, 'lutff_7/in_1')
// (22, 9, 'sp4_r_v_b_47')
// (22, 10, 'sp4_r_v_b_34')
// (22, 11, 'sp4_r_v_b_23')
// (22, 12, 'sp4_r_v_b_10')
// (23, 8, 'sp4_h_l_47')
// (23, 8, 'sp4_v_t_47')
// (23, 9, 'sp4_v_b_47')
// (23, 10, 'sp4_v_b_34')
// (23, 11, 'sp4_v_b_23')
// (23, 12, 'sp4_v_b_10')

wire n2620;
// (18, 7, 'neigh_op_tnr_6')
// (18, 8, 'neigh_op_rgt_6')
// (18, 9, 'neigh_op_bnr_6')
// (19, 6, 'sp4_r_v_b_37')
// (19, 7, 'neigh_op_top_6')
// (19, 7, 'sp4_r_v_b_24')
// (19, 8, 'ram/RDATA_1')
// (19, 8, 'sp4_r_v_b_13')
// (19, 9, 'neigh_op_bot_6')
// (19, 9, 'sp4_r_v_b_0')
// (20, 5, 'sp4_v_t_37')
// (20, 6, 'sp4_v_b_37')
// (20, 7, 'neigh_op_tnl_6')
// (20, 7, 'sp4_v_b_24')
// (20, 8, 'neigh_op_lft_6')
// (20, 8, 'sp4_v_b_13')
// (20, 9, 'neigh_op_bnl_6')
// (20, 9, 'sp4_h_r_6')
// (20, 9, 'sp4_v_b_0')
// (21, 9, 'sp4_h_r_19')
// (22, 9, 'local_g3_6')
// (22, 9, 'lutff_6/in_1')
// (22, 9, 'sp4_h_r_30')
// (23, 9, 'sp4_h_r_43')
// (24, 9, 'sp4_h_l_43')

reg n2621 = 0;
// (18, 7, 'sp4_h_r_10')
// (19, 5, 'local_g1_2')
// (19, 5, 'ram/RADDR_0')
// (19, 5, 'sp4_h_r_10')
// (19, 7, 'local_g0_7')
// (19, 7, 'ram/RADDR_0')
// (19, 7, 'sp4_h_r_23')
// (20, 4, 'sp4_r_v_b_38')
// (20, 5, 'sp4_h_r_23')
// (20, 5, 'sp4_r_v_b_27')
// (20, 6, 'local_g2_6')
// (20, 6, 'lutff_0/in_2')
// (20, 6, 'lutff_1/in_3')
// (20, 6, 'sp4_r_v_b_14')
// (20, 7, 'sp4_h_r_34')
// (20, 7, 'sp4_r_v_b_3')
// (21, 3, 'sp4_v_t_38')
// (21, 4, 'sp4_v_b_38')
// (21, 5, 'sp4_h_r_34')
// (21, 5, 'sp4_v_b_27')
// (21, 6, 'sp4_v_b_14')
// (21, 7, 'sp4_h_r_10')
// (21, 7, 'sp4_h_r_47')
// (21, 7, 'sp4_v_b_3')
// (22, 5, 'sp4_h_r_47')
// (22, 6, 'neigh_op_tnr_1')
// (22, 6, 'sp4_r_v_b_47')
// (22, 7, 'neigh_op_rgt_1')
// (22, 7, 'sp4_h_l_47')
// (22, 7, 'sp4_h_r_23')
// (22, 7, 'sp4_h_r_7')
// (22, 7, 'sp4_r_v_b_34')
// (22, 8, 'neigh_op_bnr_1')
// (22, 8, 'sp4_r_v_b_23')
// (22, 9, 'sp4_r_v_b_10')
// (23, 5, 'sp4_h_l_47')
// (23, 5, 'sp4_v_t_47')
// (23, 6, 'neigh_op_top_1')
// (23, 6, 'sp4_v_b_47')
// (23, 7, 'local_g1_1')
// (23, 7, 'lutff_1/in_1')
// (23, 7, 'lutff_1/out')
// (23, 7, 'sp4_h_r_18')
// (23, 7, 'sp4_h_r_34')
// (23, 7, 'sp4_v_b_34')
// (23, 8, 'neigh_op_bot_1')
// (23, 8, 'sp4_v_b_23')
// (23, 9, 'sp4_v_b_10')
// (24, 6, 'neigh_op_tnl_1')
// (24, 7, 'neigh_op_lft_1')
// (24, 7, 'sp4_h_r_31')
// (24, 7, 'sp4_h_r_47')
// (24, 8, 'neigh_op_bnl_1')
// (25, 7, 'sp4_h_l_47')
// (25, 7, 'sp4_h_r_42')

wire n2622;
// (18, 7, 'sp4_h_r_4')
// (19, 6, 'neigh_op_tnr_6')
// (19, 7, 'neigh_op_rgt_6')
// (19, 7, 'sp4_h_r_17')
// (19, 8, 'neigh_op_bnr_6')
// (20, 6, 'neigh_op_top_6')
// (20, 7, 'lutff_6/out')
// (20, 7, 'sp4_h_r_28')
// (20, 8, 'neigh_op_bot_6')
// (21, 6, 'neigh_op_tnl_6')
// (21, 7, 'neigh_op_lft_6')
// (21, 7, 'sp4_h_r_41')
// (21, 8, 'neigh_op_bnl_6')
// (22, 7, 'local_g1_0')
// (22, 7, 'lutff_3/in_0')
// (22, 7, 'sp4_h_l_41')
// (22, 7, 'sp4_h_r_0')
// (23, 7, 'sp4_h_r_13')
// (24, 7, 'sp4_h_r_24')
// (25, 7, 'sp4_h_r_37')

wire n2623;
// (18, 7, 'sp4_h_r_7')
// (19, 5, 'local_g0_2')
// (19, 5, 'ram/RCLKE')
// (19, 5, 'sp4_h_r_2')
// (19, 7, 'local_g0_2')
// (19, 7, 'ram/RCLKE')
// (19, 7, 'sp4_h_r_18')
// (20, 5, 'sp4_h_r_15')
// (20, 7, 'sp4_h_r_31')
// (21, 5, 'sp4_h_r_26')
// (21, 7, 'neigh_op_tnr_2')
// (21, 7, 'sp4_h_r_42')
// (21, 8, 'local_g3_2')
// (21, 8, 'lutff_5/in_2')
// (21, 8, 'neigh_op_rgt_2')
// (21, 8, 'sp4_r_v_b_36')
// (21, 9, 'neigh_op_bnr_2')
// (21, 9, 'sp4_r_v_b_25')
// (21, 10, 'sp4_r_v_b_12')
// (21, 11, 'sp4_r_v_b_1')
// (22, 5, 'sp4_h_r_39')
// (22, 6, 'sp4_r_v_b_45')
// (22, 7, 'neigh_op_top_2')
// (22, 7, 'sp4_h_l_42')
// (22, 7, 'sp4_r_v_b_32')
// (22, 7, 'sp4_v_t_36')
// (22, 8, 'lutff_2/out')
// (22, 8, 'sp4_r_v_b_21')
// (22, 8, 'sp4_v_b_36')
// (22, 9, 'neigh_op_bot_2')
// (22, 9, 'sp4_r_v_b_8')
// (22, 9, 'sp4_v_b_25')
// (22, 10, 'sp4_v_b_12')
// (22, 11, 'sp4_v_b_1')
// (23, 5, 'sp4_h_l_39')
// (23, 5, 'sp4_v_t_45')
// (23, 6, 'sp4_v_b_45')
// (23, 7, 'neigh_op_tnl_2')
// (23, 7, 'sp4_v_b_32')
// (23, 8, 'neigh_op_lft_2')
// (23, 8, 'sp4_v_b_21')
// (23, 9, 'neigh_op_bnl_2')
// (23, 9, 'sp4_v_b_8')

reg n2624 = 0;
// (18, 9, 'local_g1_4')
// (18, 9, 'lutff_4/in_3')
// (18, 9, 'sp4_h_r_4')
// (19, 8, 'neigh_op_tnr_6')
// (19, 9, 'neigh_op_rgt_6')
// (19, 9, 'sp4_h_r_17')
// (19, 10, 'neigh_op_bnr_6')
// (20, 8, 'neigh_op_top_6')
// (20, 9, 'lutff_6/out')
// (20, 9, 'sp4_h_r_28')
// (20, 10, 'neigh_op_bot_6')
// (21, 8, 'neigh_op_tnl_6')
// (21, 9, 'neigh_op_lft_6')
// (21, 9, 'sp4_h_r_41')
// (21, 10, 'neigh_op_bnl_6')
// (22, 9, 'sp4_h_l_41')

wire n2625;
// (18, 9, 'neigh_op_tnr_4')
// (18, 10, 'neigh_op_rgt_4')
// (18, 11, 'neigh_op_bnr_4')
// (19, 7, 'sp4_r_v_b_44')
// (19, 8, 'sp4_r_v_b_33')
// (19, 9, 'neigh_op_top_4')
// (19, 9, 'sp4_r_v_b_20')
// (19, 10, 'ram/RDATA_3')
// (19, 10, 'sp4_r_v_b_9')
// (19, 11, 'neigh_op_bot_4')
// (20, 6, 'sp4_v_t_44')
// (20, 7, 'sp4_v_b_44')
// (20, 8, 'sp4_v_b_33')
// (20, 9, 'neigh_op_tnl_4')
// (20, 9, 'sp4_v_b_20')
// (20, 10, 'neigh_op_lft_4')
// (20, 10, 'sp4_h_r_3')
// (20, 10, 'sp4_v_b_9')
// (20, 11, 'neigh_op_bnl_4')
// (21, 10, 'local_g1_6')
// (21, 10, 'lutff_2/in_3')
// (21, 10, 'sp4_h_r_14')
// (22, 10, 'sp4_h_r_27')
// (23, 10, 'sp4_h_r_38')
// (24, 10, 'sp4_h_l_38')

wire n2626;
// (18, 9, 'neigh_op_tnr_5')
// (18, 9, 'sp4_r_v_b_39')
// (18, 10, 'neigh_op_rgt_5')
// (18, 10, 'sp4_r_v_b_26')
// (18, 11, 'neigh_op_bnr_5')
// (18, 11, 'sp4_r_v_b_15')
// (18, 12, 'local_g1_2')
// (18, 12, 'lutff_2/in_3')
// (18, 12, 'sp4_r_v_b_2')
// (19, 8, 'sp4_v_t_39')
// (19, 9, 'neigh_op_top_5')
// (19, 9, 'sp4_v_b_39')
// (19, 10, 'ram/RDATA_2')
// (19, 10, 'sp4_v_b_26')
// (19, 11, 'neigh_op_bot_5')
// (19, 11, 'sp4_v_b_15')
// (19, 12, 'sp4_v_b_2')
// (20, 9, 'neigh_op_tnl_5')
// (20, 10, 'neigh_op_lft_5')
// (20, 11, 'neigh_op_bnl_5')

wire n2627;
// (18, 9, 'neigh_op_tnr_6')
// (18, 10, 'neigh_op_rgt_6')
// (18, 10, 'sp4_r_v_b_44')
// (18, 11, 'neigh_op_bnr_6')
// (18, 11, 'sp4_r_v_b_33')
// (18, 12, 'local_g3_4')
// (18, 12, 'lutff_3/in_0')
// (18, 12, 'sp4_r_v_b_20')
// (18, 13, 'sp4_r_v_b_9')
// (19, 9, 'neigh_op_top_6')
// (19, 9, 'sp4_v_t_44')
// (19, 10, 'ram/RDATA_1')
// (19, 10, 'sp4_v_b_44')
// (19, 11, 'neigh_op_bot_6')
// (19, 11, 'sp4_v_b_33')
// (19, 12, 'sp4_v_b_20')
// (19, 13, 'sp4_v_b_9')
// (20, 9, 'neigh_op_tnl_6')
// (20, 10, 'neigh_op_lft_6')
// (20, 11, 'neigh_op_bnl_6')

wire n2628;
// (18, 9, 'neigh_op_tnr_7')
// (18, 10, 'neigh_op_rgt_7')
// (18, 10, 'sp4_h_r_3')
// (18, 11, 'neigh_op_bnr_7')
// (19, 9, 'neigh_op_top_7')
// (19, 10, 'ram/RDATA_0')
// (19, 10, 'sp4_h_r_14')
// (19, 11, 'neigh_op_bot_7')
// (20, 9, 'neigh_op_tnl_7')
// (20, 10, 'neigh_op_lft_7')
// (20, 10, 'sp4_h_r_27')
// (20, 11, 'neigh_op_bnl_7')
// (21, 10, 'local_g2_6')
// (21, 10, 'lutff_5/in_1')
// (21, 10, 'sp4_h_r_38')
// (22, 10, 'sp4_h_l_38')

reg n2629 = 0;
// (18, 10, 'local_g0_0')
// (18, 10, 'lutff_5/in_1')
// (18, 10, 'sp4_h_r_8')
// (19, 10, 'sp4_h_r_21')
// (20, 10, 'neigh_op_tnr_3')
// (20, 10, 'sp4_h_r_32')
// (20, 11, 'neigh_op_rgt_3')
// (20, 12, 'neigh_op_bnr_3')
// (21, 10, 'neigh_op_top_3')
// (21, 10, 'sp4_h_r_45')
// (21, 11, 'lutff_3/out')
// (21, 11, 'sp4_r_v_b_39')
// (21, 12, 'neigh_op_bot_3')
// (21, 12, 'sp4_r_v_b_26')
// (21, 13, 'sp4_r_v_b_15')
// (21, 14, 'sp4_r_v_b_2')
// (22, 10, 'neigh_op_tnl_3')
// (22, 10, 'sp4_h_l_45')
// (22, 10, 'sp4_v_t_39')
// (22, 11, 'neigh_op_lft_3')
// (22, 11, 'sp4_v_b_39')
// (22, 12, 'neigh_op_bnl_3')
// (22, 12, 'sp4_v_b_26')
// (22, 13, 'sp4_v_b_15')
// (22, 14, 'sp4_v_b_2')

reg n2630 = 0;
// (18, 10, 'local_g0_2')
// (18, 10, 'lutff_1/in_3')
// (18, 10, 'sp4_h_r_2')
// (19, 9, 'neigh_op_tnr_5')
// (19, 10, 'neigh_op_rgt_5')
// (19, 10, 'sp4_h_r_15')
// (19, 11, 'neigh_op_bnr_5')
// (20, 9, 'neigh_op_top_5')
// (20, 10, 'lutff_5/out')
// (20, 10, 'sp4_h_r_26')
// (20, 11, 'neigh_op_bot_5')
// (21, 9, 'neigh_op_tnl_5')
// (21, 10, 'neigh_op_lft_5')
// (21, 10, 'sp4_h_r_39')
// (21, 11, 'neigh_op_bnl_5')
// (22, 10, 'sp4_h_l_39')

reg n2631 = 0;
// (18, 10, 'local_g0_6')
// (18, 10, 'lutff_3/in_3')
// (18, 10, 'sp4_h_r_6')
// (19, 9, 'neigh_op_tnr_7')
// (19, 10, 'neigh_op_rgt_7')
// (19, 10, 'sp4_h_r_19')
// (19, 11, 'neigh_op_bnr_7')
// (20, 9, 'neigh_op_top_7')
// (20, 10, 'lutff_7/out')
// (20, 10, 'sp4_h_r_30')
// (20, 11, 'neigh_op_bot_7')
// (21, 9, 'neigh_op_tnl_7')
// (21, 10, 'neigh_op_lft_7')
// (21, 10, 'sp4_h_r_43')
// (21, 11, 'neigh_op_bnl_7')
// (22, 10, 'sp4_h_l_43')

wire n2632;
// (18, 10, 'neigh_op_tnr_0')
// (18, 11, 'neigh_op_rgt_0')
// (18, 12, 'neigh_op_bnr_0')
// (19, 10, 'neigh_op_top_0')
// (19, 11, 'ram/RDATA_15')
// (19, 12, 'neigh_op_bot_0')
// (20, 10, 'neigh_op_tnl_0')
// (20, 11, 'local_g1_0')
// (20, 11, 'lutff_1/in_0')
// (20, 11, 'neigh_op_lft_0')
// (20, 12, 'neigh_op_bnl_0')

wire n2633;
// (18, 10, 'neigh_op_tnr_2')
// (18, 11, 'neigh_op_rgt_2')
// (18, 12, 'local_g0_2')
// (18, 12, 'lutff_0/in_2')
// (18, 12, 'neigh_op_bnr_2')
// (19, 10, 'neigh_op_top_2')
// (19, 11, 'ram/RDATA_13')
// (19, 12, 'neigh_op_bot_2')
// (20, 10, 'neigh_op_tnl_2')
// (20, 11, 'neigh_op_lft_2')
// (20, 12, 'neigh_op_bnl_2')

wire n2634;
// (18, 10, 'neigh_op_tnr_3')
// (18, 11, 'local_g3_3')
// (18, 11, 'lutff_0/in_0')
// (18, 11, 'neigh_op_rgt_3')
// (18, 12, 'neigh_op_bnr_3')
// (19, 10, 'neigh_op_top_3')
// (19, 11, 'ram/RDATA_12')
// (19, 12, 'neigh_op_bot_3')
// (20, 10, 'neigh_op_tnl_3')
// (20, 11, 'neigh_op_lft_3')
// (20, 12, 'neigh_op_bnl_3')

wire n2635;
// (18, 10, 'neigh_op_tnr_4')
// (18, 11, 'neigh_op_rgt_4')
// (18, 12, 'neigh_op_bnr_4')
// (19, 10, 'neigh_op_top_4')
// (19, 11, 'ram/RDATA_11')
// (19, 12, 'neigh_op_bot_4')
// (20, 10, 'neigh_op_tnl_4')
// (20, 11, 'local_g1_4')
// (20, 11, 'lutff_4/in_1')
// (20, 11, 'neigh_op_lft_4')
// (20, 12, 'neigh_op_bnl_4')

wire n2636;
// (18, 10, 'neigh_op_tnr_5')
// (18, 11, 'neigh_op_rgt_5')
// (18, 12, 'local_g0_5')
// (18, 12, 'lutff_6/in_3')
// (18, 12, 'neigh_op_bnr_5')
// (19, 10, 'neigh_op_top_5')
// (19, 11, 'ram/RDATA_10')
// (19, 12, 'neigh_op_bot_5')
// (20, 10, 'neigh_op_tnl_5')
// (20, 11, 'neigh_op_lft_5')
// (20, 12, 'neigh_op_bnl_5')

wire n2637;
// (18, 10, 'neigh_op_tnr_6')
// (18, 11, 'local_g0_1')
// (18, 11, 'lutff_6/in_1')
// (18, 11, 'neigh_op_rgt_6')
// (18, 11, 'sp4_h_r_1')
// (18, 12, 'neigh_op_bnr_6')
// (19, 10, 'neigh_op_top_6')
// (19, 11, 'ram/RDATA_9')
// (19, 11, 'sp4_h_r_12')
// (19, 12, 'neigh_op_bot_6')
// (20, 10, 'neigh_op_tnl_6')
// (20, 11, 'neigh_op_lft_6')
// (20, 11, 'sp4_h_r_25')
// (20, 12, 'neigh_op_bnl_6')
// (21, 11, 'sp4_h_r_36')
// (22, 11, 'sp4_h_l_36')

wire n2638;
// (18, 10, 'neigh_op_tnr_7')
// (18, 11, 'local_g2_7')
// (18, 11, 'lutff_5/in_0')
// (18, 11, 'neigh_op_rgt_7')
// (18, 12, 'neigh_op_bnr_7')
// (19, 10, 'neigh_op_top_7')
// (19, 11, 'ram/RDATA_8')
// (19, 12, 'neigh_op_bot_7')
// (20, 10, 'neigh_op_tnl_7')
// (20, 11, 'neigh_op_lft_7')
// (20, 12, 'neigh_op_bnl_7')

reg n2639 = 0;
// (18, 11, 'local_g1_1')
// (18, 11, 'lutff_3/in_1')
// (18, 11, 'sp4_h_r_9')
// (19, 11, 'sp4_h_r_20')
// (20, 10, 'neigh_op_tnr_6')
// (20, 11, 'neigh_op_rgt_6')
// (20, 11, 'sp4_h_r_33')
// (20, 12, 'neigh_op_bnr_6')
// (21, 10, 'neigh_op_top_6')
// (21, 11, 'lutff_6/out')
// (21, 11, 'sp4_h_r_44')
// (21, 12, 'neigh_op_bot_6')
// (22, 10, 'neigh_op_tnl_6')
// (22, 11, 'neigh_op_lft_6')
// (22, 11, 'sp4_h_l_44')
// (22, 12, 'neigh_op_bnl_6')

wire n2640;
// (18, 11, 'local_g2_3')
// (18, 11, 'lutff_7/in_0')
// (18, 11, 'neigh_op_tnr_3')
// (18, 12, 'neigh_op_rgt_3')
// (18, 13, 'neigh_op_bnr_3')
// (19, 11, 'neigh_op_top_3')
// (19, 12, 'ram/RDATA_4')
// (19, 13, 'neigh_op_bot_3')
// (20, 11, 'neigh_op_tnl_3')
// (20, 12, 'neigh_op_lft_3')
// (20, 13, 'neigh_op_bnl_3')

wire n2641;
// (18, 11, 'local_g2_6')
// (18, 11, 'lutff_4/in_2')
// (18, 11, 'neigh_op_tnr_6')
// (18, 12, 'neigh_op_rgt_6')
// (18, 13, 'neigh_op_bnr_6')
// (19, 11, 'neigh_op_top_6')
// (19, 12, 'ram/RDATA_1')
// (19, 13, 'neigh_op_bot_6')
// (20, 11, 'neigh_op_tnl_6')
// (20, 12, 'neigh_op_lft_6')
// (20, 13, 'neigh_op_bnl_6')

wire n2642;
// (18, 11, 'neigh_op_tnr_0')
// (18, 12, 'neigh_op_rgt_0')
// (18, 13, 'neigh_op_bnr_0')
// (19, 11, 'neigh_op_top_0')
// (19, 12, 'ram/RDATA_7')
// (19, 13, 'neigh_op_bot_0')
// (20, 11, 'local_g2_0')
// (20, 11, 'lutff_3/in_1')
// (20, 11, 'neigh_op_tnl_0')
// (20, 12, 'neigh_op_lft_0')
// (20, 13, 'neigh_op_bnl_0')

wire n2643;
// (18, 11, 'neigh_op_tnr_1')
// (18, 12, 'neigh_op_rgt_1')
// (18, 13, 'neigh_op_bnr_1')
// (19, 11, 'neigh_op_top_1')
// (19, 12, 'ram/RDATA_6')
// (19, 13, 'neigh_op_bot_1')
// (20, 11, 'local_g3_1')
// (20, 11, 'lutff_2/in_0')
// (20, 11, 'neigh_op_tnl_1')
// (20, 12, 'neigh_op_lft_1')
// (20, 13, 'neigh_op_bnl_1')

wire n2644;
// (18, 11, 'neigh_op_tnr_4')
// (18, 12, 'neigh_op_rgt_4')
// (18, 13, 'neigh_op_bnr_4')
// (19, 11, 'neigh_op_top_4')
// (19, 12, 'ram/RDATA_3')
// (19, 13, 'neigh_op_bot_4')
// (20, 11, 'local_g3_4')
// (20, 11, 'lutff_6/in_3')
// (20, 11, 'neigh_op_tnl_4')
// (20, 12, 'neigh_op_lft_4')
// (20, 13, 'neigh_op_bnl_4')

wire n2645;
// (18, 11, 'neigh_op_tnr_5')
// (18, 12, 'local_g3_5')
// (18, 12, 'lutff_5/in_3')
// (18, 12, 'neigh_op_rgt_5')
// (18, 13, 'neigh_op_bnr_5')
// (19, 11, 'neigh_op_top_5')
// (19, 12, 'ram/RDATA_2')
// (19, 13, 'neigh_op_bot_5')
// (20, 11, 'neigh_op_tnl_5')
// (20, 12, 'neigh_op_lft_5')
// (20, 13, 'neigh_op_bnl_5')

wire n2646;
// (18, 11, 'neigh_op_tnr_7')
// (18, 12, 'neigh_op_rgt_7')
// (18, 13, 'neigh_op_bnr_7')
// (19, 11, 'neigh_op_top_7')
// (19, 12, 'ram/RDATA_0')
// (19, 13, 'neigh_op_bot_7')
// (20, 11, 'local_g2_7')
// (20, 11, 'lutff_0/in_1')
// (20, 11, 'neigh_op_tnl_7')
// (20, 12, 'neigh_op_lft_7')
// (20, 13, 'neigh_op_bnl_7')

wire n2647;
// (18, 12, 'local_g3_2')
// (18, 12, 'lutff_4/in_1')
// (18, 12, 'neigh_op_tnr_2')
// (18, 13, 'neigh_op_rgt_2')
// (18, 14, 'neigh_op_bnr_2')
// (19, 12, 'neigh_op_top_2')
// (19, 13, 'ram/RDATA_13')
// (19, 14, 'neigh_op_bot_2')
// (20, 12, 'neigh_op_tnl_2')
// (20, 13, 'neigh_op_lft_2')
// (20, 14, 'neigh_op_bnl_2')

wire n2648;
// (18, 12, 'neigh_op_tnr_0')
// (18, 13, 'local_g2_0')
// (18, 13, 'lutff_4/in_2')
// (18, 13, 'neigh_op_rgt_0')
// (18, 14, 'neigh_op_bnr_0')
// (19, 12, 'neigh_op_top_0')
// (19, 13, 'ram/RDATA_15')
// (19, 14, 'neigh_op_bot_0')
// (20, 12, 'neigh_op_tnl_0')
// (20, 13, 'neigh_op_lft_0')
// (20, 14, 'neigh_op_bnl_0')

wire n2649;
// (18, 12, 'neigh_op_tnr_1')
// (18, 13, 'local_g3_1')
// (18, 13, 'lutff_1/in_3')
// (18, 13, 'neigh_op_rgt_1')
// (18, 14, 'neigh_op_bnr_1')
// (19, 12, 'neigh_op_top_1')
// (19, 13, 'ram/RDATA_14')
// (19, 14, 'neigh_op_bot_1')
// (20, 12, 'neigh_op_tnl_1')
// (20, 13, 'neigh_op_lft_1')
// (20, 14, 'neigh_op_bnl_1')

wire n2650;
// (18, 12, 'neigh_op_tnr_3')
// (18, 13, 'neigh_op_rgt_3')
// (18, 14, 'neigh_op_bnr_3')
// (19, 12, 'neigh_op_top_3')
// (19, 13, 'ram/RDATA_12')
// (19, 13, 'sp4_r_v_b_39')
// (19, 14, 'neigh_op_bot_3')
// (19, 14, 'sp4_r_v_b_26')
// (19, 15, 'sp4_r_v_b_15')
// (19, 16, 'sp4_r_v_b_2')
// (20, 12, 'neigh_op_tnl_3')
// (20, 12, 'sp4_h_r_2')
// (20, 12, 'sp4_v_t_39')
// (20, 13, 'neigh_op_lft_3')
// (20, 13, 'sp4_v_b_39')
// (20, 14, 'neigh_op_bnl_3')
// (20, 14, 'sp4_v_b_26')
// (20, 15, 'sp4_v_b_15')
// (20, 16, 'sp4_v_b_2')
// (21, 12, 'sp4_h_r_15')
// (22, 12, 'local_g2_2')
// (22, 12, 'lutff_0/in_0')
// (22, 12, 'sp4_h_r_26')
// (23, 12, 'sp4_h_r_39')
// (24, 12, 'sp4_h_l_39')

wire n2651;
// (18, 12, 'neigh_op_tnr_4')
// (18, 13, 'neigh_op_rgt_4')
// (18, 14, 'local_g0_4')
// (18, 14, 'lutff_4/in_0')
// (18, 14, 'neigh_op_bnr_4')
// (19, 12, 'neigh_op_top_4')
// (19, 13, 'ram/RDATA_11')
// (19, 14, 'neigh_op_bot_4')
// (20, 12, 'neigh_op_tnl_4')
// (20, 13, 'neigh_op_lft_4')
// (20, 14, 'neigh_op_bnl_4')

wire n2652;
// (18, 12, 'neigh_op_tnr_5')
// (18, 13, 'local_g3_5')
// (18, 13, 'lutff_7/in_1')
// (18, 13, 'neigh_op_rgt_5')
// (18, 14, 'neigh_op_bnr_5')
// (19, 12, 'neigh_op_top_5')
// (19, 13, 'ram/RDATA_10')
// (19, 14, 'neigh_op_bot_5')
// (20, 12, 'neigh_op_tnl_5')
// (20, 13, 'neigh_op_lft_5')
// (20, 14, 'neigh_op_bnl_5')

wire n2653;
// (18, 12, 'neigh_op_tnr_6')
// (18, 13, 'neigh_op_rgt_6')
// (18, 14, 'neigh_op_bnr_6')
// (19, 12, 'neigh_op_top_6')
// (19, 13, 'ram/RDATA_9')
// (19, 14, 'neigh_op_bot_6')
// (20, 12, 'neigh_op_tnl_6')
// (20, 13, 'neigh_op_lft_6')
// (20, 14, 'local_g2_6')
// (20, 14, 'lutff_6/in_2')
// (20, 14, 'neigh_op_bnl_6')

wire n2654;
// (18, 12, 'neigh_op_tnr_7')
// (18, 13, 'local_g2_7')
// (18, 13, 'lutff_3/in_0')
// (18, 13, 'neigh_op_rgt_7')
// (18, 14, 'neigh_op_bnr_7')
// (19, 12, 'neigh_op_top_7')
// (19, 13, 'ram/RDATA_8')
// (19, 14, 'neigh_op_bot_7')
// (20, 12, 'neigh_op_tnl_7')
// (20, 13, 'neigh_op_lft_7')
// (20, 14, 'neigh_op_bnl_7')

wire n2655;
// (18, 13, 'local_g2_3')
// (18, 13, 'lutff_5/in_0')
// (18, 13, 'neigh_op_tnr_3')
// (18, 14, 'neigh_op_rgt_3')
// (18, 15, 'neigh_op_bnr_3')
// (19, 13, 'neigh_op_top_3')
// (19, 14, 'ram/RDATA_4')
// (19, 15, 'neigh_op_bot_3')
// (20, 13, 'neigh_op_tnl_3')
// (20, 14, 'neigh_op_lft_3')
// (20, 15, 'neigh_op_bnl_3')

wire n2656;
// (18, 13, 'local_g2_6')
// (18, 13, 'lutff_0/in_2')
// (18, 13, 'neigh_op_tnr_6')
// (18, 14, 'neigh_op_rgt_6')
// (18, 15, 'neigh_op_bnr_6')
// (19, 13, 'neigh_op_top_6')
// (19, 14, 'ram/RDATA_1')
// (19, 15, 'neigh_op_bot_6')
// (20, 13, 'neigh_op_tnl_6')
// (20, 14, 'neigh_op_lft_6')
// (20, 15, 'neigh_op_bnl_6')

wire n2657;
// (18, 13, 'local_g3_0')
// (18, 13, 'lutff_6/in_3')
// (18, 13, 'neigh_op_tnr_0')
// (18, 14, 'neigh_op_rgt_0')
// (18, 15, 'neigh_op_bnr_0')
// (19, 13, 'neigh_op_top_0')
// (19, 14, 'ram/RDATA_7')
// (19, 15, 'neigh_op_bot_0')
// (20, 13, 'neigh_op_tnl_0')
// (20, 14, 'neigh_op_lft_0')
// (20, 15, 'neigh_op_bnl_0')

wire n2658;
// (18, 13, 'local_g3_7')
// (18, 13, 'lutff_2/in_0')
// (18, 13, 'neigh_op_tnr_7')
// (18, 14, 'neigh_op_rgt_7')
// (18, 15, 'neigh_op_bnr_7')
// (19, 13, 'neigh_op_top_7')
// (19, 14, 'ram/RDATA_0')
// (19, 15, 'neigh_op_bot_7')
// (20, 13, 'neigh_op_tnl_7')
// (20, 14, 'neigh_op_lft_7')
// (20, 15, 'neigh_op_bnl_7')

wire n2659;
// (18, 13, 'neigh_op_tnr_1')
// (18, 14, 'local_g3_1')
// (18, 14, 'lutff_2/in_0')
// (18, 14, 'neigh_op_rgt_1')
// (18, 15, 'neigh_op_bnr_1')
// (19, 13, 'neigh_op_top_1')
// (19, 14, 'ram/RDATA_6')
// (19, 15, 'neigh_op_bot_1')
// (20, 13, 'neigh_op_tnl_1')
// (20, 14, 'neigh_op_lft_1')
// (20, 15, 'neigh_op_bnl_1')

wire n2660;
// (18, 13, 'neigh_op_tnr_2')
// (18, 14, 'neigh_op_rgt_2')
// (18, 15, 'neigh_op_bnr_2')
// (19, 13, 'neigh_op_top_2')
// (19, 14, 'ram/RDATA_5')
// (19, 15, 'neigh_op_bot_2')
// (20, 13, 'neigh_op_tnl_2')
// (20, 14, 'local_g1_2')
// (20, 14, 'lutff_4/in_3')
// (20, 14, 'neigh_op_lft_2')
// (20, 15, 'neigh_op_bnl_2')

wire n2661;
// (18, 13, 'neigh_op_tnr_4')
// (18, 14, 'neigh_op_rgt_4')
// (18, 15, 'neigh_op_bnr_4')
// (19, 13, 'neigh_op_top_4')
// (19, 14, 'ram/RDATA_3')
// (19, 15, 'neigh_op_bot_4')
// (20, 13, 'neigh_op_tnl_4')
// (20, 14, 'local_g0_4')
// (20, 14, 'lutff_5/in_3')
// (20, 14, 'neigh_op_lft_4')
// (20, 15, 'neigh_op_bnl_4')

wire n2662;
// (18, 13, 'neigh_op_tnr_5')
// (18, 14, 'local_g2_5')
// (18, 14, 'lutff_1/in_2')
// (18, 14, 'neigh_op_rgt_5')
// (18, 15, 'neigh_op_bnr_5')
// (19, 13, 'neigh_op_top_5')
// (19, 14, 'ram/RDATA_2')
// (19, 15, 'neigh_op_bot_5')
// (20, 13, 'neigh_op_tnl_5')
// (20, 14, 'neigh_op_lft_5')
// (20, 15, 'neigh_op_bnl_5')

wire n2663;
// (18, 13, 'sp4_h_r_11')
// (19, 12, 'sp4_h_r_10')
// (19, 13, 'sp4_h_r_22')
// (20, 12, 'sp4_h_r_23')
// (20, 13, 'local_g3_3')
// (20, 13, 'lutff_global/cen')
// (20, 13, 'sp4_h_r_35')
// (21, 10, 'sp4_r_v_b_45')
// (21, 11, 'sp4_r_v_b_32')
// (21, 12, 'local_g2_2')
// (21, 12, 'lutff_global/cen')
// (21, 12, 'neigh_op_tnr_4')
// (21, 12, 'sp4_h_r_34')
// (21, 12, 'sp4_r_v_b_21')
// (21, 13, 'neigh_op_rgt_4')
// (21, 13, 'sp4_h_r_46')
// (21, 13, 'sp4_r_v_b_8')
// (21, 14, 'neigh_op_bnr_4')
// (22, 9, 'sp4_v_t_45')
// (22, 10, 'sp4_v_b_45')
// (22, 11, 'sp4_v_b_32')
// (22, 12, 'local_g0_4')
// (22, 12, 'lutff_1/in_1')
// (22, 12, 'neigh_op_top_4')
// (22, 12, 'sp4_h_r_47')
// (22, 12, 'sp4_v_b_21')
// (22, 13, 'local_g0_2')
// (22, 13, 'lutff_4/out')
// (22, 13, 'lutff_global/cen')
// (22, 13, 'sp4_h_l_46')
// (22, 13, 'sp4_h_r_2')
// (22, 13, 'sp4_h_r_8')
// (22, 13, 'sp4_r_v_b_41')
// (22, 13, 'sp4_v_b_8')
// (22, 14, 'neigh_op_bot_4')
// (22, 14, 'sp4_r_v_b_28')
// (22, 15, 'sp4_r_v_b_17')
// (22, 16, 'sp4_r_v_b_4')
// (23, 12, 'neigh_op_tnl_4')
// (23, 12, 'sp4_h_l_47')
// (23, 12, 'sp4_v_t_41')
// (23, 13, 'neigh_op_lft_4')
// (23, 13, 'sp4_h_r_15')
// (23, 13, 'sp4_h_r_21')
// (23, 13, 'sp4_v_b_41')
// (23, 14, 'neigh_op_bnl_4')
// (23, 14, 'sp4_v_b_28')
// (23, 15, 'sp4_v_b_17')
// (23, 16, 'sp4_v_b_4')
// (24, 13, 'sp4_h_r_26')
// (24, 13, 'sp4_h_r_32')
// (25, 13, 'sp4_h_r_39')
// (25, 13, 'sp4_h_r_45')

wire n2664;
// (18, 13, 'sp4_r_v_b_40')
// (18, 14, 'sp4_r_v_b_29')
// (18, 15, 'sp4_r_v_b_16')
// (18, 16, 'sp4_r_v_b_5')
// (19, 9, 'sp4_r_v_b_43')
// (19, 10, 'local_g0_6')
// (19, 10, 'local_g1_6')
// (19, 10, 'ram/MASK_0')
// (19, 10, 'ram/MASK_1')
// (19, 10, 'ram/MASK_2')
// (19, 10, 'ram/MASK_3')
// (19, 10, 'sp4_r_v_b_30')
// (19, 11, 'local_g2_3')
// (19, 11, 'local_g3_3')
// (19, 11, 'neigh_op_tnr_3')
// (19, 11, 'ram/MASK_10')
// (19, 11, 'ram/MASK_11')
// (19, 11, 'ram/MASK_12')
// (19, 11, 'ram/MASK_13')
// (19, 11, 'ram/MASK_14')
// (19, 11, 'ram/MASK_15')
// (19, 11, 'ram/MASK_8')
// (19, 11, 'ram/MASK_9')
// (19, 11, 'sp4_r_v_b_19')
// (19, 12, 'local_g2_3')
// (19, 12, 'local_g3_3')
// (19, 12, 'neigh_op_rgt_3')
// (19, 12, 'ram/MASK_0')
// (19, 12, 'ram/MASK_1')
// (19, 12, 'ram/MASK_2')
// (19, 12, 'ram/MASK_3')
// (19, 12, 'ram/MASK_4')
// (19, 12, 'ram/MASK_5')
// (19, 12, 'ram/MASK_6')
// (19, 12, 'ram/MASK_7')
// (19, 12, 'sp4_h_r_11')
// (19, 12, 'sp4_r_v_b_38')
// (19, 12, 'sp4_r_v_b_6')
// (19, 12, 'sp4_v_t_40')
// (19, 13, 'local_g0_3')
// (19, 13, 'local_g1_3')
// (19, 13, 'neigh_op_bnr_3')
// (19, 13, 'ram/MASK_10')
// (19, 13, 'ram/MASK_11')
// (19, 13, 'ram/MASK_12')
// (19, 13, 'ram/MASK_13')
// (19, 13, 'ram/MASK_14')
// (19, 13, 'ram/MASK_15')
// (19, 13, 'ram/MASK_8')
// (19, 13, 'ram/MASK_9')
// (19, 13, 'sp4_r_v_b_27')
// (19, 13, 'sp4_v_b_40')
// (19, 14, 'local_g2_5')
// (19, 14, 'local_g2_6')
// (19, 14, 'ram/MASK_0')
// (19, 14, 'ram/MASK_1')
// (19, 14, 'ram/MASK_2')
// (19, 14, 'ram/MASK_3')
// (19, 14, 'ram/MASK_4')
// (19, 14, 'ram/MASK_5')
// (19, 14, 'ram/MASK_6')
// (19, 14, 'ram/MASK_7')
// (19, 14, 'sp4_r_v_b_14')
// (19, 14, 'sp4_v_b_29')
// (19, 15, 'sp4_r_v_b_3')
// (19, 15, 'sp4_v_b_16')
// (19, 16, 'sp4_v_b_5')
// (20, 8, 'sp4_v_t_43')
// (20, 9, 'sp4_v_b_43')
// (20, 10, 'sp4_v_b_30')
// (20, 11, 'neigh_op_top_3')
// (20, 11, 'sp4_v_b_19')
// (20, 11, 'sp4_v_t_38')
// (20, 12, 'lutff_3/out')
// (20, 12, 'sp4_h_r_22')
// (20, 12, 'sp4_v_b_38')
// (20, 12, 'sp4_v_b_6')
// (20, 13, 'neigh_op_bot_3')
// (20, 13, 'sp4_v_b_27')
// (20, 14, 'sp4_v_b_14')
// (20, 15, 'sp4_v_b_3')
// (21, 11, 'neigh_op_tnl_3')
// (21, 12, 'neigh_op_lft_3')
// (21, 12, 'sp4_h_r_35')
// (21, 13, 'neigh_op_bnl_3')
// (22, 12, 'sp4_h_r_46')
// (23, 12, 'sp4_h_l_46')

wire io_19_31_1;
// (18, 16, 'sp4_r_v_b_38')
// (18, 17, 'sp4_r_v_b_27')
// (18, 18, 'sp4_r_v_b_14')
// (18, 19, 'sp4_r_v_b_3')
// (18, 20, 'sp4_r_v_b_38')
// (18, 21, 'sp4_r_v_b_27')
// (18, 22, 'sp4_r_v_b_14')
// (18, 23, 'sp4_r_v_b_3')
// (18, 24, 'sp4_r_v_b_43')
// (18, 25, 'sp4_r_v_b_30')
// (18, 26, 'sp4_r_v_b_19')
// (18, 27, 'sp4_r_v_b_6')
// (18, 28, 'sp4_r_v_b_39')
// (18, 29, 'sp4_r_v_b_26')
// (18, 30, 'sp4_r_v_b_15')
// (19, 14, 'neigh_op_tnr_7')
// (19, 15, 'neigh_op_rgt_7')
// (19, 15, 'sp4_h_r_3')
// (19, 15, 'sp4_v_t_38')
// (19, 16, 'neigh_op_bnr_7')
// (19, 16, 'sp4_v_b_38')
// (19, 17, 'sp4_v_b_27')
// (19, 18, 'sp4_v_b_14')
// (19, 19, 'sp4_v_b_3')
// (19, 19, 'sp4_v_t_38')
// (19, 20, 'sp4_v_b_38')
// (19, 21, 'sp4_v_b_27')
// (19, 22, 'sp4_v_b_14')
// (19, 23, 'sp4_v_b_3')
// (19, 23, 'sp4_v_t_43')
// (19, 24, 'sp4_v_b_43')
// (19, 25, 'sp4_v_b_30')
// (19, 26, 'sp4_v_b_19')
// (19, 27, 'sp4_v_b_6')
// (19, 27, 'sp4_v_t_39')
// (19, 28, 'sp4_v_b_39')
// (19, 29, 'sp4_v_b_26')
// (19, 30, 'sp4_v_b_15')
// (19, 31, 'io_1/D_OUT_0')
// (19, 31, 'io_1/PAD')
// (19, 31, 'local_g1_2')
// (19, 31, 'span4_vert_2')
// (20, 14, 'neigh_op_top_7')
// (20, 15, 'lutff_7/out')
// (20, 15, 'sp4_h_r_14')
// (20, 16, 'neigh_op_bot_7')
// (21, 14, 'neigh_op_tnl_7')
// (21, 15, 'neigh_op_lft_7')
// (21, 15, 'sp4_h_r_27')
// (21, 16, 'neigh_op_bnl_7')
// (22, 15, 'sp4_h_r_38')
// (23, 15, 'sp4_h_l_38')

wire n2666;
// (18, 18, 'sp4_h_r_9')
// (19, 18, 'sp4_h_r_20')
// (20, 17, 'neigh_op_tnr_6')
// (20, 18, 'neigh_op_rgt_6')
// (20, 18, 'sp4_h_r_33')
// (20, 19, 'neigh_op_bnr_6')
// (21, 15, 'sp4_r_v_b_38')
// (21, 16, 'sp4_r_v_b_27')
// (21, 17, 'neigh_op_top_6')
// (21, 17, 'sp4_r_v_b_14')
// (21, 18, 'local_g1_3')
// (21, 18, 'lutff_6/out')
// (21, 18, 'lutff_global/cen')
// (21, 18, 'sp4_h_r_44')
// (21, 18, 'sp4_r_v_b_3')
// (21, 19, 'neigh_op_bot_6')
// (22, 14, 'sp4_v_t_38')
// (22, 15, 'sp4_v_b_38')
// (22, 16, 'sp4_v_b_27')
// (22, 17, 'neigh_op_tnl_6')
// (22, 17, 'sp4_v_b_14')
// (22, 18, 'neigh_op_lft_6')
// (22, 18, 'sp4_h_l_44')
// (22, 18, 'sp4_v_b_3')
// (22, 19, 'neigh_op_bnl_6')

reg n2667 = 0;
// (18, 19, 'local_g0_4')
// (18, 19, 'lutff_5/in_3')
// (18, 19, 'sp4_h_r_4')
// (19, 18, 'neigh_op_tnr_6')
// (19, 19, 'neigh_op_rgt_6')
// (19, 19, 'sp4_h_r_17')
// (19, 20, 'neigh_op_bnr_6')
// (20, 18, 'neigh_op_top_6')
// (20, 19, 'lutff_6/out')
// (20, 19, 'sp4_h_r_28')
// (20, 20, 'neigh_op_bot_6')
// (21, 18, 'neigh_op_tnl_6')
// (21, 19, 'neigh_op_lft_6')
// (21, 19, 'sp4_h_r_41')
// (21, 20, 'neigh_op_bnl_6')
// (22, 19, 'sp4_h_l_41')

reg n2668 = 0;
// (19, 1, 'neigh_op_tnr_0')
// (19, 2, 'neigh_op_rgt_0')
// (19, 3, 'neigh_op_bnr_0')
// (20, 1, 'neigh_op_top_0')
// (20, 2, 'local_g0_0')
// (20, 2, 'lutff_0/out')
// (20, 2, 'lutff_4/in_2')
// (20, 3, 'neigh_op_bot_0')
// (21, 1, 'neigh_op_tnl_0')
// (21, 2, 'neigh_op_lft_0')
// (21, 3, 'neigh_op_bnl_0')

reg n2669 = 0;
// (19, 1, 'neigh_op_tnr_6')
// (19, 2, 'neigh_op_rgt_6')
// (19, 3, 'neigh_op_bnr_6')
// (20, 1, 'neigh_op_top_6')
// (20, 2, 'local_g0_6')
// (20, 2, 'lutff_4/in_0')
// (20, 2, 'lutff_6/out')
// (20, 3, 'neigh_op_bot_6')
// (21, 1, 'neigh_op_tnl_6')
// (21, 2, 'neigh_op_lft_6')
// (21, 3, 'neigh_op_bnl_6')

wire n2670;
// (19, 3, 'neigh_op_tnr_1')
// (19, 4, 'neigh_op_rgt_1')
// (19, 5, 'neigh_op_bnr_1')
// (20, 3, 'neigh_op_top_1')
// (20, 4, 'lutff_1/out')
// (20, 5, 'neigh_op_bot_1')
// (21, 3, 'neigh_op_tnl_1')
// (21, 4, 'local_g0_1')
// (21, 4, 'lutff_4/in_1')
// (21, 4, 'neigh_op_lft_1')
// (21, 5, 'neigh_op_bnl_1')

wire n2671;
// (19, 3, 'neigh_op_tnr_3')
// (19, 4, 'neigh_op_rgt_3')
// (19, 5, 'neigh_op_bnr_3')
// (20, 3, 'neigh_op_top_3')
// (20, 4, 'lutff_3/out')
// (20, 5, 'neigh_op_bot_3')
// (21, 3, 'neigh_op_tnl_3')
// (21, 4, 'local_g0_3')
// (21, 4, 'lutff_7/in_2')
// (21, 4, 'neigh_op_lft_3')
// (21, 5, 'neigh_op_bnl_3')

wire n2672;
// (19, 3, 'neigh_op_tnr_7')
// (19, 4, 'neigh_op_rgt_7')
// (19, 5, 'neigh_op_bnr_7')
// (20, 3, 'neigh_op_top_7')
// (20, 4, 'lutff_7/out')
// (20, 5, 'neigh_op_bot_7')
// (21, 3, 'neigh_op_tnl_7')
// (21, 4, 'local_g0_7')
// (21, 4, 'lutff_0/in_1')
// (21, 4, 'neigh_op_lft_7')
// (21, 5, 'neigh_op_bnl_7')

reg n2673 = 0;
// (19, 4, 'neigh_op_tnr_2')
// (19, 5, 'neigh_op_rgt_2')
// (19, 5, 'sp4_h_r_9')
// (19, 6, 'neigh_op_bnr_2')
// (20, 4, 'local_g1_2')
// (20, 4, 'lutff_4/in_3')
// (20, 4, 'lutff_5/in_2')
// (20, 4, 'neigh_op_top_2')
// (20, 5, 'local_g3_2')
// (20, 5, 'lutff_2/in_1')
// (20, 5, 'lutff_2/out')
// (20, 5, 'lutff_7/in_2')
// (20, 5, 'sp4_h_r_20')
// (20, 5, 'sp4_h_r_4')
// (20, 6, 'neigh_op_bot_2')
// (21, 4, 'neigh_op_tnl_2')
// (21, 5, 'neigh_op_lft_2')
// (21, 5, 'sp4_h_r_17')
// (21, 5, 'sp4_h_r_33')
// (21, 6, 'neigh_op_bnl_2')
// (22, 2, 'sp4_r_v_b_38')
// (22, 3, 'sp4_r_v_b_27')
// (22, 4, 'local_g2_6')
// (22, 4, 'lutff_3/in_1')
// (22, 4, 'sp4_r_v_b_14')
// (22, 5, 'local_g3_4')
// (22, 5, 'lutff_0/in_1')
// (22, 5, 'lutff_2/in_3')
// (22, 5, 'sp4_h_r_28')
// (22, 5, 'sp4_h_r_44')
// (22, 5, 'sp4_r_v_b_3')
// (23, 1, 'sp4_v_t_38')
// (23, 2, 'sp4_v_b_38')
// (23, 3, 'sp4_v_b_27')
// (23, 4, 'sp4_v_b_14')
// (23, 5, 'sp4_h_l_44')
// (23, 5, 'sp4_h_r_41')
// (23, 5, 'sp4_v_b_3')
// (24, 5, 'sp4_h_l_41')

reg n2674 = 0;
// (19, 4, 'neigh_op_tnr_3')
// (19, 5, 'neigh_op_rgt_3')
// (19, 5, 'sp4_h_r_11')
// (19, 6, 'neigh_op_bnr_3')
// (20, 4, 'local_g0_3')
// (20, 4, 'lutff_4/in_1')
// (20, 4, 'lutff_5/in_0')
// (20, 4, 'neigh_op_top_3')
// (20, 5, 'local_g0_3')
// (20, 5, 'lutff_1/in_2')
// (20, 5, 'lutff_3/in_2')
// (20, 5, 'lutff_3/out')
// (20, 5, 'lutff_7/in_0')
// (20, 5, 'sp4_h_r_22')
// (20, 5, 'sp4_h_r_6')
// (20, 6, 'neigh_op_bot_3')
// (21, 4, 'neigh_op_tnl_3')
// (21, 5, 'neigh_op_lft_3')
// (21, 5, 'sp4_h_r_19')
// (21, 5, 'sp4_h_r_35')
// (21, 6, 'neigh_op_bnl_3')
// (22, 2, 'sp4_r_v_b_40')
// (22, 3, 'sp4_r_v_b_29')
// (22, 4, 'local_g3_0')
// (22, 4, 'lutff_3/in_0')
// (22, 4, 'sp4_r_v_b_16')
// (22, 5, 'local_g2_6')
// (22, 5, 'lutff_0/in_0')
// (22, 5, 'lutff_2/in_0')
// (22, 5, 'sp4_h_r_30')
// (22, 5, 'sp4_h_r_46')
// (22, 5, 'sp4_r_v_b_5')
// (23, 1, 'sp4_v_t_40')
// (23, 2, 'sp4_v_b_40')
// (23, 3, 'sp4_v_b_29')
// (23, 4, 'sp4_v_b_16')
// (23, 5, 'sp4_h_l_46')
// (23, 5, 'sp4_h_r_43')
// (23, 5, 'sp4_v_b_5')
// (24, 5, 'sp4_h_l_43')

reg n2675 = 0;
// (19, 4, 'neigh_op_tnr_5')
// (19, 5, 'neigh_op_rgt_5')
// (19, 5, 'sp4_r_v_b_42')
// (19, 6, 'neigh_op_bnr_5')
// (19, 6, 'sp4_r_v_b_31')
// (19, 7, 'sp4_r_v_b_18')
// (19, 8, 'sp4_r_v_b_7')
// (20, 4, 'local_g1_5')
// (20, 4, 'lutff_4/in_2')
// (20, 4, 'lutff_5/in_1')
// (20, 4, 'neigh_op_top_5')
// (20, 4, 'sp4_h_r_0')
// (20, 4, 'sp4_v_t_42')
// (20, 5, 'local_g3_5')
// (20, 5, 'lutff_0/in_2')
// (20, 5, 'lutff_3/in_3')
// (20, 5, 'lutff_5/in_1')
// (20, 5, 'lutff_5/out')
// (20, 5, 'lutff_7/in_1')
// (20, 5, 'sp4_h_r_10')
// (20, 5, 'sp4_v_b_42')
// (20, 6, 'neigh_op_bot_5')
// (20, 6, 'sp4_v_b_31')
// (20, 7, 'sp4_v_b_18')
// (20, 8, 'sp4_v_b_7')
// (21, 4, 'neigh_op_tnl_5')
// (21, 4, 'sp4_h_r_13')
// (21, 5, 'neigh_op_lft_5')
// (21, 5, 'sp4_h_r_23')
// (21, 6, 'neigh_op_bnl_5')
// (22, 4, 'local_g2_0')
// (22, 4, 'lutff_3/in_3')
// (22, 4, 'sp4_h_r_24')
// (22, 5, 'local_g3_2')
// (22, 5, 'lutff_0/in_3')
// (22, 5, 'lutff_2/in_1')
// (22, 5, 'sp4_h_r_34')
// (23, 4, 'sp4_h_r_37')
// (23, 5, 'sp4_h_r_47')
// (24, 4, 'sp4_h_l_37')
// (24, 5, 'sp4_h_l_47')

wire n2676;
// (19, 4, 'sp4_r_v_b_43')
// (19, 5, 'sp4_r_v_b_30')
// (19, 6, 'sp4_r_v_b_19')
// (19, 7, 'sp4_r_v_b_6')
// (20, 3, 'sp4_v_t_43')
// (20, 4, 'sp4_v_b_43')
// (20, 5, 'sp4_v_b_30')
// (20, 6, 'local_g1_3')
// (20, 6, 'lutff_global/cen')
// (20, 6, 'sp4_v_b_19')
// (20, 7, 'sp4_h_r_1')
// (20, 7, 'sp4_v_b_6')
// (21, 7, 'sp4_h_r_12')
// (22, 6, 'neigh_op_tnr_2')
// (22, 7, 'neigh_op_rgt_2')
// (22, 7, 'sp4_h_r_25')
// (22, 8, 'neigh_op_bnr_2')
// (23, 6, 'neigh_op_top_2')
// (23, 7, 'local_g2_2')
// (23, 7, 'lutff_2/out')
// (23, 7, 'lutff_global/cen')
// (23, 7, 'sp4_h_r_36')
// (23, 8, 'neigh_op_bot_2')
// (24, 6, 'neigh_op_tnl_2')
// (24, 7, 'neigh_op_lft_2')
// (24, 7, 'sp4_h_l_36')
// (24, 8, 'neigh_op_bnl_2')

reg n2677 = 0;
// (19, 5, 'local_g3_1')
// (19, 5, 'neigh_op_tnr_1')
// (19, 5, 'ram/RADDR_1')
// (19, 6, 'neigh_op_rgt_1')
// (19, 7, 'local_g1_1')
// (19, 7, 'neigh_op_bnr_1')
// (19, 7, 'ram/RADDR_1')
// (20, 5, 'neigh_op_top_1')
// (20, 6, 'local_g0_1')
// (20, 6, 'lutff_1/in_2')
// (20, 6, 'lutff_1/out')
// (20, 7, 'neigh_op_bot_1')
// (21, 5, 'neigh_op_tnl_1')
// (21, 6, 'neigh_op_lft_1')
// (21, 7, 'neigh_op_bnl_1')

reg n2678 = 0;
// (19, 5, 'local_g3_2')
// (19, 5, 'neigh_op_tnr_2')
// (19, 5, 'ram/RADDR_2')
// (19, 6, 'neigh_op_rgt_2')
// (19, 7, 'local_g1_2')
// (19, 7, 'neigh_op_bnr_2')
// (19, 7, 'ram/RADDR_2')
// (20, 5, 'neigh_op_top_2')
// (20, 6, 'local_g0_2')
// (20, 6, 'lutff_2/in_2')
// (20, 6, 'lutff_2/out')
// (20, 7, 'neigh_op_bot_2')
// (21, 5, 'neigh_op_tnl_2')
// (21, 6, 'neigh_op_lft_2')
// (21, 7, 'neigh_op_bnl_2')

reg n2679 = 0;
// (19, 5, 'local_g3_3')
// (19, 5, 'neigh_op_tnr_3')
// (19, 5, 'ram/RADDR_3')
// (19, 6, 'neigh_op_rgt_3')
// (19, 7, 'local_g1_3')
// (19, 7, 'neigh_op_bnr_3')
// (19, 7, 'ram/RADDR_3')
// (20, 5, 'neigh_op_top_3')
// (20, 6, 'local_g3_3')
// (20, 6, 'lutff_3/in_1')
// (20, 6, 'lutff_3/out')
// (20, 7, 'neigh_op_bot_3')
// (21, 5, 'neigh_op_tnl_3')
// (21, 6, 'neigh_op_lft_3')
// (21, 7, 'neigh_op_bnl_3')

reg n2680 = 0;
// (19, 5, 'local_g3_4')
// (19, 5, 'neigh_op_tnr_4')
// (19, 5, 'ram/RADDR_4')
// (19, 6, 'neigh_op_rgt_4')
// (19, 7, 'local_g1_4')
// (19, 7, 'neigh_op_bnr_4')
// (19, 7, 'ram/RADDR_4')
// (20, 5, 'neigh_op_top_4')
// (20, 6, 'local_g2_4')
// (20, 6, 'lutff_4/in_2')
// (20, 6, 'lutff_4/out')
// (20, 7, 'neigh_op_bot_4')
// (21, 5, 'neigh_op_tnl_4')
// (21, 6, 'neigh_op_lft_4')
// (21, 7, 'neigh_op_bnl_4')

reg n2681 = 0;
// (19, 5, 'local_g3_5')
// (19, 5, 'neigh_op_tnr_5')
// (19, 5, 'ram/RADDR_5')
// (19, 6, 'neigh_op_rgt_5')
// (19, 7, 'local_g1_5')
// (19, 7, 'neigh_op_bnr_5')
// (19, 7, 'ram/RADDR_5')
// (20, 5, 'neigh_op_top_5')
// (20, 6, 'local_g0_5')
// (20, 6, 'lutff_5/in_2')
// (20, 6, 'lutff_5/out')
// (20, 7, 'neigh_op_bot_5')
// (21, 5, 'neigh_op_tnl_5')
// (21, 6, 'neigh_op_lft_5')
// (21, 7, 'neigh_op_bnl_5')

reg n2682 = 0;
// (19, 5, 'local_g3_6')
// (19, 5, 'neigh_op_tnr_6')
// (19, 5, 'ram/RADDR_6')
// (19, 6, 'neigh_op_rgt_6')
// (19, 7, 'local_g1_6')
// (19, 7, 'neigh_op_bnr_6')
// (19, 7, 'ram/RADDR_6')
// (20, 5, 'neigh_op_top_6')
// (20, 6, 'local_g3_6')
// (20, 6, 'lutff_6/in_1')
// (20, 6, 'lutff_6/out')
// (20, 7, 'neigh_op_bot_6')
// (21, 5, 'neigh_op_tnl_6')
// (21, 6, 'neigh_op_lft_6')
// (21, 7, 'neigh_op_bnl_6')

wire n2683;
// (19, 5, 'sp4_r_v_b_47')
// (19, 6, 'local_g2_2')
// (19, 6, 'ram/WCLKE')
// (19, 6, 'sp4_r_v_b_34')
// (19, 7, 'neigh_op_tnr_5')
// (19, 7, 'sp4_r_v_b_23')
// (19, 8, 'local_g2_2')
// (19, 8, 'neigh_op_rgt_5')
// (19, 8, 'ram/WCLKE')
// (19, 8, 'sp4_r_v_b_10')
// (19, 9, 'neigh_op_bnr_5')
// (20, 4, 'sp4_v_t_47')
// (20, 5, 'local_g2_7')
// (20, 5, 'lutff_6/in_1')
// (20, 5, 'sp4_v_b_47')
// (20, 6, 'sp4_v_b_34')
// (20, 7, 'neigh_op_top_5')
// (20, 7, 'sp4_v_b_23')
// (20, 8, 'lutff_5/out')
// (20, 8, 'sp4_v_b_10')
// (20, 9, 'neigh_op_bot_5')
// (21, 7, 'neigh_op_tnl_5')
// (21, 8, 'neigh_op_lft_5')
// (21, 9, 'neigh_op_bnl_5')

wire n2684;
// (19, 6, 'neigh_op_tnr_2')
// (19, 7, 'neigh_op_rgt_2')
// (19, 8, 'neigh_op_bnr_2')
// (20, 6, 'neigh_op_top_2')
// (20, 7, 'lutff_2/out')
// (20, 7, 'sp4_h_r_4')
// (20, 8, 'neigh_op_bot_2')
// (21, 6, 'neigh_op_tnl_2')
// (21, 7, 'neigh_op_lft_2')
// (21, 7, 'sp4_h_r_17')
// (21, 8, 'neigh_op_bnl_2')
// (22, 7, 'local_g3_4')
// (22, 7, 'lutff_2/in_3')
// (22, 7, 'sp4_h_r_28')
// (23, 7, 'sp4_h_r_41')
// (24, 7, 'sp4_h_l_41')

wire n2685;
// (19, 6, 'neigh_op_tnr_4')
// (19, 7, 'neigh_op_rgt_4')
// (19, 8, 'neigh_op_bnr_4')
// (20, 4, 'sp4_r_v_b_44')
// (20, 5, 'sp4_r_v_b_33')
// (20, 6, 'neigh_op_top_4')
// (20, 6, 'sp4_r_v_b_20')
// (20, 7, 'lutff_4/out')
// (20, 7, 'sp4_r_v_b_9')
// (20, 8, 'neigh_op_bot_4')
// (21, 3, 'sp4_v_t_44')
// (21, 4, 'sp4_v_b_44')
// (21, 5, 'sp4_v_b_33')
// (21, 6, 'neigh_op_tnl_4')
// (21, 6, 'sp4_v_b_20')
// (21, 7, 'neigh_op_lft_4')
// (21, 7, 'sp4_h_r_3')
// (21, 7, 'sp4_v_b_9')
// (21, 8, 'neigh_op_bnl_4')
// (22, 7, 'local_g1_6')
// (22, 7, 'lutff_6/in_1')
// (22, 7, 'sp4_h_r_14')
// (23, 7, 'sp4_h_r_27')
// (24, 7, 'sp4_h_r_38')
// (25, 7, 'sp4_h_l_38')

wire n2686;
// (19, 6, 'sp4_h_r_11')
// (20, 6, 'sp4_h_r_22')
// (21, 6, 'local_g3_3')
// (21, 6, 'lutff_global/cen')
// (21, 6, 'sp4_h_r_35')
// (21, 7, 'neigh_op_tnr_6')
// (21, 8, 'neigh_op_rgt_6')
// (21, 9, 'neigh_op_bnr_6')
// (22, 2, 'sp12_v_t_23')
// (22, 3, 'sp12_v_b_23')
// (22, 4, 'sp12_v_b_20')
// (22, 5, 'sp12_v_b_19')
// (22, 6, 'sp12_v_b_16')
// (22, 6, 'sp4_h_r_46')
// (22, 7, 'neigh_op_top_6')
// (22, 7, 'sp12_v_b_15')
// (22, 7, 'sp4_r_v_b_40')
// (22, 8, 'lutff_6/out')
// (22, 8, 'sp12_v_b_12')
// (22, 8, 'sp4_r_v_b_29')
// (22, 9, 'local_g3_3')
// (22, 9, 'lutff_global/cen')
// (22, 9, 'neigh_op_bot_6')
// (22, 9, 'sp12_v_b_11')
// (22, 9, 'sp4_r_v_b_16')
// (22, 10, 'sp12_v_b_8')
// (22, 10, 'sp4_r_v_b_5')
// (22, 11, 'sp12_v_b_7')
// (22, 12, 'sp12_v_b_4')
// (22, 13, 'sp12_v_b_3')
// (22, 14, 'sp12_v_b_0')
// (23, 6, 'sp4_h_l_46')
// (23, 6, 'sp4_v_t_40')
// (23, 7, 'neigh_op_tnl_6')
// (23, 7, 'sp4_v_b_40')
// (23, 8, 'local_g0_6')
// (23, 8, 'lutff_1/in_3')
// (23, 8, 'neigh_op_lft_6')
// (23, 8, 'sp4_v_b_29')
// (23, 9, 'neigh_op_bnl_6')
// (23, 9, 'sp4_v_b_16')
// (23, 10, 'sp4_v_b_5')

wire n2687;
// (19, 7, 'neigh_op_tnr_0')
// (19, 8, 'neigh_op_rgt_0')
// (19, 9, 'neigh_op_bnr_0')
// (20, 7, 'neigh_op_top_0')
// (20, 8, 'lutff_0/out')
// (20, 9, 'neigh_op_bot_0')
// (21, 7, 'neigh_op_tnl_0')
// (21, 8, 'local_g1_0')
// (21, 8, 'lutff_7/in_0')
// (21, 8, 'neigh_op_lft_0')
// (21, 9, 'neigh_op_bnl_0')

wire n2688;
// (19, 7, 'neigh_op_tnr_2')
// (19, 8, 'neigh_op_rgt_2')
// (19, 9, 'neigh_op_bnr_2')
// (20, 7, 'neigh_op_top_2')
// (20, 8, 'lutff_2/out')
// (20, 9, 'neigh_op_bot_2')
// (21, 7, 'neigh_op_tnl_2')
// (21, 8, 'local_g1_2')
// (21, 8, 'lutff_6/in_1')
// (21, 8, 'neigh_op_lft_2')
// (21, 9, 'neigh_op_bnl_2')

wire n2689;
// (19, 7, 'neigh_op_tnr_4')
// (19, 8, 'neigh_op_rgt_4')
// (19, 9, 'neigh_op_bnr_4')
// (20, 7, 'neigh_op_top_4')
// (20, 8, 'lutff_4/out')
// (20, 9, 'neigh_op_bot_4')
// (21, 7, 'neigh_op_tnl_4')
// (21, 8, 'local_g0_4')
// (21, 8, 'lutff_4/in_0')
// (21, 8, 'neigh_op_lft_4')
// (21, 9, 'neigh_op_bnl_4')

reg n2690 = 0;
// (19, 7, 'sp4_h_r_1')
// (20, 7, 'local_g0_4')
// (20, 7, 'lutff_3/in_1')
// (20, 7, 'sp4_h_r_12')
// (21, 6, 'neigh_op_tnr_2')
// (21, 7, 'local_g3_2')
// (21, 7, 'lutff_3/in_2')
// (21, 7, 'neigh_op_rgt_2')
// (21, 7, 'sp4_h_r_25')
// (21, 8, 'neigh_op_bnr_2')
// (22, 6, 'neigh_op_top_2')
// (22, 7, 'local_g2_2')
// (22, 7, 'lutff_2/in_0')
// (22, 7, 'lutff_2/out')
// (22, 7, 'lutff_7/in_1')
// (22, 7, 'sp4_h_r_36')
// (22, 8, 'neigh_op_bot_2')
// (23, 6, 'neigh_op_tnl_2')
// (23, 7, 'neigh_op_lft_2')
// (23, 7, 'sp4_h_l_36')
// (23, 8, 'neigh_op_bnl_2')

reg n2691 = 0;
// (19, 7, 'sp4_h_r_3')
// (20, 7, 'local_g1_6')
// (20, 7, 'lutff_7/in_2')
// (20, 7, 'sp4_h_r_14')
// (21, 6, 'neigh_op_tnr_3')
// (21, 7, 'local_g2_3')
// (21, 7, 'lutff_7/in_2')
// (21, 7, 'neigh_op_rgt_3')
// (21, 7, 'sp4_h_r_27')
// (21, 8, 'neigh_op_bnr_3')
// (22, 6, 'neigh_op_top_3')
// (22, 7, 'local_g2_3')
// (22, 7, 'lutff_3/in_2')
// (22, 7, 'lutff_3/out')
// (22, 7, 'lutff_7/in_2')
// (22, 7, 'sp4_h_r_38')
// (22, 8, 'neigh_op_bot_3')
// (23, 6, 'neigh_op_tnl_3')
// (23, 7, 'neigh_op_lft_3')
// (23, 7, 'sp4_h_l_38')
// (23, 8, 'neigh_op_bnl_3')

reg n2692 = 0;
// (19, 7, 'sp4_h_r_9')
// (20, 7, 'local_g1_4')
// (20, 7, 'lutff_5/in_2')
// (20, 7, 'sp4_h_r_20')
// (21, 6, 'neigh_op_tnr_6')
// (21, 7, 'local_g2_6')
// (21, 7, 'lutff_5/in_1')
// (21, 7, 'neigh_op_rgt_6')
// (21, 7, 'sp4_h_r_33')
// (21, 8, 'neigh_op_bnr_6')
// (22, 6, 'neigh_op_top_6')
// (22, 7, 'local_g2_6')
// (22, 7, 'local_g3_6')
// (22, 7, 'lutff_6/in_2')
// (22, 7, 'lutff_6/out')
// (22, 7, 'lutff_7/in_0')
// (22, 7, 'sp4_h_r_44')
// (22, 8, 'neigh_op_bot_6')
// (23, 6, 'neigh_op_tnl_6')
// (23, 7, 'neigh_op_lft_6')
// (23, 7, 'sp4_h_l_44')
// (23, 8, 'neigh_op_bnl_6')

reg n2693 = 0;
// (19, 7, 'sp4_r_v_b_36')
// (19, 8, 'sp4_r_v_b_25')
// (19, 9, 'sp4_r_v_b_12')
// (19, 10, 'sp4_r_v_b_1')
// (20, 6, 'local_g1_1')
// (20, 6, 'lutff_7/in_3')
// (20, 6, 'sp4_h_r_1')
// (20, 6, 'sp4_v_t_36')
// (20, 7, 'sp4_v_b_36')
// (20, 8, 'local_g2_1')
// (20, 8, 'lutff_5/in_2')
// (20, 8, 'sp4_v_b_25')
// (20, 9, 'sp4_v_b_12')
// (20, 10, 'sp4_v_b_1')
// (21, 6, 'sp4_h_r_12')
// (22, 5, 'neigh_op_tnr_2')
// (22, 6, 'neigh_op_rgt_2')
// (22, 6, 'sp4_h_r_25')
// (22, 6, 'sp4_r_v_b_36')
// (22, 7, 'local_g0_2')
// (22, 7, 'lutff_5/in_3')
// (22, 7, 'neigh_op_bnr_2')
// (22, 7, 'sp4_r_v_b_25')
// (22, 8, 'local_g2_4')
// (22, 8, 'lutff_4/in_0')
// (22, 8, 'sp4_r_v_b_12')
// (22, 9, 'sp4_r_v_b_1')
// (23, 5, 'neigh_op_top_2')
// (23, 5, 'sp4_v_t_36')
// (23, 6, 'lutff_2/out')
// (23, 6, 'sp4_h_r_36')
// (23, 6, 'sp4_v_b_36')
// (23, 7, 'neigh_op_bot_2')
// (23, 7, 'sp4_v_b_25')
// (23, 8, 'sp4_v_b_12')
// (23, 9, 'sp4_v_b_1')
// (24, 5, 'neigh_op_tnl_2')
// (24, 6, 'neigh_op_lft_2')
// (24, 6, 'sp4_h_l_36')
// (24, 7, 'neigh_op_bnl_2')

wire n2694;
// (19, 8, 'sp4_h_r_11')
// (20, 8, 'sp4_h_r_22')
// (21, 6, 'neigh_op_tnr_1')
// (21, 6, 'sp4_r_v_b_47')
// (21, 7, 'local_g2_2')
// (21, 7, 'lutff_global/cen')
// (21, 7, 'neigh_op_rgt_1')
// (21, 7, 'sp4_r_v_b_34')
// (21, 8, 'local_g3_3')
// (21, 8, 'lutff_global/cen')
// (21, 8, 'neigh_op_bnr_1')
// (21, 8, 'sp4_h_r_35')
// (21, 8, 'sp4_r_v_b_23')
// (21, 9, 'sp4_r_v_b_10')
// (22, 5, 'sp4_r_v_b_43')
// (22, 5, 'sp4_v_t_47')
// (22, 6, 'neigh_op_top_1')
// (22, 6, 'sp4_r_v_b_30')
// (22, 6, 'sp4_v_b_47')
// (22, 7, 'local_g3_3')
// (22, 7, 'lutff_1/out')
// (22, 7, 'lutff_global/cen')
// (22, 7, 'sp4_r_v_b_19')
// (22, 7, 'sp4_v_b_34')
// (22, 8, 'neigh_op_bot_1')
// (22, 8, 'sp4_h_r_46')
// (22, 8, 'sp4_r_v_b_6')
// (22, 8, 'sp4_v_b_23')
// (22, 9, 'sp4_v_b_10')
// (23, 4, 'sp4_v_t_43')
// (23, 5, 'sp4_v_b_43')
// (23, 6, 'neigh_op_tnl_1')
// (23, 6, 'sp4_v_b_30')
// (23, 7, 'neigh_op_lft_1')
// (23, 7, 'sp4_v_b_19')
// (23, 8, 'neigh_op_bnl_1')
// (23, 8, 'sp4_h_l_46')
// (23, 8, 'sp4_v_b_6')

reg n2695 = 0;
// (19, 10, 'neigh_op_tnr_0')
// (19, 11, 'neigh_op_rgt_0')
// (19, 12, 'neigh_op_bnr_0')
// (20, 10, 'neigh_op_top_0')
// (20, 11, 'local_g3_0')
// (20, 11, 'lutff_0/out')
// (20, 11, 'lutff_7/in_0')
// (20, 12, 'neigh_op_bot_0')
// (21, 10, 'neigh_op_tnl_0')
// (21, 11, 'neigh_op_lft_0')
// (21, 12, 'neigh_op_bnl_0')

reg n2696 = 0;
// (19, 10, 'neigh_op_tnr_1')
// (19, 11, 'neigh_op_rgt_1')
// (19, 12, 'neigh_op_bnr_1')
// (20, 10, 'neigh_op_top_1')
// (20, 10, 'sp4_r_v_b_46')
// (20, 11, 'lutff_1/out')
// (20, 11, 'sp4_r_v_b_35')
// (20, 12, 'neigh_op_bot_1')
// (20, 12, 'sp4_r_v_b_22')
// (20, 13, 'local_g2_3')
// (20, 13, 'lutff_3/in_2')
// (20, 13, 'sp4_r_v_b_11')
// (21, 9, 'sp4_v_t_46')
// (21, 10, 'neigh_op_tnl_1')
// (21, 10, 'sp4_v_b_46')
// (21, 11, 'neigh_op_lft_1')
// (21, 11, 'sp4_v_b_35')
// (21, 12, 'neigh_op_bnl_1')
// (21, 12, 'sp4_v_b_22')
// (21, 13, 'sp4_v_b_11')

reg n2697 = 0;
// (19, 10, 'neigh_op_tnr_2')
// (19, 11, 'neigh_op_rgt_2')
// (19, 12, 'neigh_op_bnr_2')
// (20, 10, 'neigh_op_top_2')
// (20, 11, 'lutff_2/out')
// (20, 12, 'local_g1_2')
// (20, 12, 'lutff_0/in_3')
// (20, 12, 'neigh_op_bot_2')
// (21, 10, 'neigh_op_tnl_2')
// (21, 11, 'neigh_op_lft_2')
// (21, 12, 'neigh_op_bnl_2')

reg n2698 = 0;
// (19, 10, 'neigh_op_tnr_3')
// (19, 11, 'neigh_op_rgt_3')
// (19, 12, 'neigh_op_bnr_3')
// (20, 10, 'neigh_op_top_3')
// (20, 11, 'lutff_3/out')
// (20, 12, 'neigh_op_bot_3')
// (21, 10, 'neigh_op_tnl_3')
// (21, 11, 'neigh_op_lft_3')
// (21, 12, 'local_g3_3')
// (21, 12, 'lutff_4/in_2')
// (21, 12, 'neigh_op_bnl_3')

reg n2699 = 0;
// (19, 10, 'neigh_op_tnr_4')
// (19, 11, 'neigh_op_rgt_4')
// (19, 12, 'neigh_op_bnr_4')
// (20, 10, 'neigh_op_top_4')
// (20, 11, 'local_g2_4')
// (20, 11, 'lutff_4/out')
// (20, 11, 'lutff_5/in_1')
// (20, 12, 'neigh_op_bot_4')
// (21, 10, 'neigh_op_tnl_4')
// (21, 11, 'neigh_op_lft_4')
// (21, 12, 'neigh_op_bnl_4')

wire n2700;
// (19, 10, 'neigh_op_tnr_5')
// (19, 10, 'sp4_r_v_b_39')
// (19, 11, 'neigh_op_rgt_5')
// (19, 11, 'sp4_r_v_b_26')
// (19, 12, 'neigh_op_bnr_5')
// (19, 12, 'sp4_r_v_b_15')
// (19, 13, 'sp4_r_v_b_2')
// (20, 9, 'sp4_v_t_39')
// (20, 10, 'neigh_op_top_5')
// (20, 10, 'sp4_v_b_39')
// (20, 11, 'lutff_5/out')
// (20, 11, 'sp4_v_b_26')
// (20, 12, 'neigh_op_bot_5')
// (20, 12, 'sp4_v_b_15')
// (20, 13, 'local_g0_2')
// (20, 13, 'lutff_6/in_0')
// (20, 13, 'sp4_v_b_2')
// (21, 10, 'neigh_op_tnl_5')
// (21, 11, 'neigh_op_lft_5')
// (21, 12, 'neigh_op_bnl_5')

reg n2701 = 0;
// (19, 10, 'neigh_op_tnr_6')
// (19, 11, 'neigh_op_rgt_6')
// (19, 12, 'neigh_op_bnr_6')
// (20, 10, 'neigh_op_top_6')
// (20, 11, 'local_g3_6')
// (20, 11, 'lutff_5/in_0')
// (20, 11, 'lutff_6/out')
// (20, 12, 'neigh_op_bot_6')
// (21, 10, 'neigh_op_tnl_6')
// (21, 11, 'neigh_op_lft_6')
// (21, 12, 'neigh_op_bnl_6')

wire n2702;
// (19, 10, 'neigh_op_tnr_7')
// (19, 11, 'neigh_op_rgt_7')
// (19, 12, 'neigh_op_bnr_7')
// (20, 10, 'neigh_op_top_7')
// (20, 11, 'lutff_7/out')
// (20, 11, 'sp4_r_v_b_47')
// (20, 12, 'neigh_op_bot_7')
// (20, 12, 'sp4_r_v_b_34')
// (20, 13, 'local_g3_7')
// (20, 13, 'lutff_7/in_3')
// (20, 13, 'sp4_r_v_b_23')
// (20, 14, 'sp4_r_v_b_10')
// (21, 10, 'neigh_op_tnl_7')
// (21, 10, 'sp4_v_t_47')
// (21, 11, 'neigh_op_lft_7')
// (21, 11, 'sp4_v_b_47')
// (21, 12, 'neigh_op_bnl_7')
// (21, 12, 'sp4_v_b_34')
// (21, 13, 'sp4_v_b_23')
// (21, 14, 'sp4_v_b_10')

wire n2703;
// (19, 11, 'neigh_op_tnr_0')
// (19, 12, 'neigh_op_rgt_0')
// (19, 13, 'neigh_op_bnr_0')
// (20, 11, 'neigh_op_top_0')
// (20, 12, 'lutff_0/out')
// (20, 13, 'local_g1_0')
// (20, 13, 'lutff_2/in_1')
// (20, 13, 'neigh_op_bot_0')
// (21, 11, 'neigh_op_tnl_0')
// (21, 12, 'neigh_op_lft_0')
// (21, 13, 'neigh_op_bnl_0')

wire n2704;
// (19, 11, 'neigh_op_tnr_1')
// (19, 12, 'neigh_op_rgt_1')
// (19, 13, 'neigh_op_bnr_1')
// (20, 11, 'local_g1_1')
// (20, 11, 'lutff_5/in_3')
// (20, 11, 'lutff_7/in_1')
// (20, 11, 'neigh_op_top_1')
// (20, 12, 'local_g2_1')
// (20, 12, 'lutff_0/in_1')
// (20, 12, 'lutff_1/out')
// (20, 13, 'neigh_op_bot_1')
// (21, 11, 'neigh_op_tnl_1')
// (21, 12, 'local_g1_1')
// (21, 12, 'lutff_4/in_0')
// (21, 12, 'neigh_op_lft_1')
// (21, 13, 'neigh_op_bnl_1')

wire n2705;
// (19, 11, 'neigh_op_tnr_6')
// (19, 12, 'neigh_op_rgt_6')
// (19, 13, 'neigh_op_bnr_6')
// (20, 11, 'local_g1_6')
// (20, 11, 'lutff_5/in_2')
// (20, 11, 'lutff_7/in_2')
// (20, 11, 'neigh_op_top_6')
// (20, 12, 'local_g2_6')
// (20, 12, 'lutff_0/in_0')
// (20, 12, 'lutff_6/out')
// (20, 13, 'local_g1_6')
// (20, 13, 'lutff_3/in_0')
// (20, 13, 'neigh_op_bot_6')
// (21, 11, 'neigh_op_tnl_6')
// (21, 12, 'neigh_op_lft_6')
// (21, 13, 'neigh_op_bnl_6')

reg n2706 = 0;
// (19, 12, 'neigh_op_tnr_0')
// (19, 13, 'neigh_op_rgt_0')
// (19, 14, 'neigh_op_bnr_0')
// (20, 12, 'neigh_op_top_0')
// (20, 13, 'lutff_0/out')
// (20, 14, 'neigh_op_bot_0')
// (21, 12, 'neigh_op_tnl_0')
// (21, 13, 'neigh_op_lft_0')
// (21, 14, 'local_g3_0')
// (21, 14, 'lutff_4/in_1')
// (21, 14, 'neigh_op_bnl_0')

wire n2707;
// (19, 12, 'neigh_op_tnr_1')
// (19, 13, 'neigh_op_rgt_1')
// (19, 14, 'neigh_op_bnr_1')
// (20, 12, 'neigh_op_top_1')
// (20, 13, 'local_g1_1')
// (20, 13, 'lutff_1/out')
// (20, 13, 'lutff_3/in_1')
// (20, 14, 'neigh_op_bot_1')
// (21, 12, 'neigh_op_tnl_1')
// (21, 13, 'neigh_op_lft_1')
// (21, 14, 'neigh_op_bnl_1')

reg n2708 = 0;
// (19, 12, 'neigh_op_tnr_2')
// (19, 13, 'neigh_op_rgt_2')
// (19, 14, 'neigh_op_bnr_2')
// (20, 12, 'neigh_op_top_2')
// (20, 13, 'lutff_2/out')
// (20, 14, 'neigh_op_bot_2')
// (21, 12, 'neigh_op_tnl_2')
// (21, 13, 'neigh_op_lft_2')
// (21, 14, 'local_g3_2')
// (21, 14, 'lutff_4/in_3')
// (21, 14, 'neigh_op_bnl_2')

reg n2709 = 0;
// (19, 12, 'neigh_op_tnr_3')
// (19, 13, 'neigh_op_rgt_3')
// (19, 14, 'neigh_op_bnr_3')
// (20, 12, 'neigh_op_top_3')
// (20, 13, 'lutff_3/out')
// (20, 14, 'neigh_op_bot_3')
// (21, 12, 'neigh_op_tnl_3')
// (21, 13, 'neigh_op_lft_3')
// (21, 14, 'local_g3_3')
// (21, 14, 'lutff_7/in_3')
// (21, 14, 'neigh_op_bnl_3')

reg n2710 = 0;
// (19, 12, 'neigh_op_tnr_4')
// (19, 13, 'neigh_op_rgt_4')
// (19, 14, 'neigh_op_bnr_4')
// (20, 12, 'neigh_op_top_4')
// (20, 13, 'lutff_4/out')
// (20, 14, 'neigh_op_bot_4')
// (21, 12, 'neigh_op_tnl_4')
// (21, 13, 'neigh_op_lft_4')
// (21, 14, 'local_g3_4')
// (21, 14, 'lutff_0/in_1')
// (21, 14, 'neigh_op_bnl_4')

reg n2711 = 0;
// (19, 12, 'neigh_op_tnr_5')
// (19, 13, 'neigh_op_rgt_5')
// (19, 14, 'neigh_op_bnr_5')
// (20, 12, 'neigh_op_top_5')
// (20, 13, 'lutff_5/out')
// (20, 13, 'sp4_h_r_10')
// (20, 14, 'neigh_op_bot_5')
// (21, 12, 'neigh_op_tnl_5')
// (21, 13, 'neigh_op_lft_5')
// (21, 13, 'sp4_h_r_23')
// (21, 14, 'neigh_op_bnl_5')
// (22, 13, 'sp4_h_r_34')
// (23, 13, 'local_g2_7')
// (23, 13, 'lutff_6/in_1')
// (23, 13, 'sp4_h_r_47')
// (24, 13, 'sp4_h_l_47')

reg n2712 = 0;
// (19, 12, 'neigh_op_tnr_6')
// (19, 13, 'neigh_op_rgt_6')
// (19, 14, 'neigh_op_bnr_6')
// (20, 12, 'neigh_op_top_6')
// (20, 13, 'lutff_6/out')
// (20, 14, 'neigh_op_bot_6')
// (21, 12, 'neigh_op_tnl_6')
// (21, 13, 'neigh_op_lft_6')
// (21, 14, 'local_g3_6')
// (21, 14, 'lutff_2/in_1')
// (21, 14, 'neigh_op_bnl_6')

reg n2713 = 0;
// (19, 12, 'neigh_op_tnr_7')
// (19, 13, 'neigh_op_rgt_7')
// (19, 13, 'sp4_h_r_3')
// (19, 14, 'neigh_op_bnr_7')
// (20, 12, 'neigh_op_top_7')
// (20, 13, 'lutff_7/out')
// (20, 13, 'sp4_h_r_14')
// (20, 14, 'neigh_op_bot_7')
// (21, 12, 'neigh_op_tnl_7')
// (21, 13, 'neigh_op_lft_7')
// (21, 13, 'sp4_h_r_27')
// (21, 14, 'neigh_op_bnl_7')
// (22, 13, 'sp4_h_r_38')
// (23, 13, 'local_g0_3')
// (23, 13, 'lutff_0/in_3')
// (23, 13, 'sp4_h_l_38')
// (23, 13, 'sp4_h_r_11')
// (24, 13, 'sp4_h_r_22')
// (25, 13, 'sp4_h_r_35')

wire n2714;
// (19, 13, 'neigh_op_tnr_2')
// (19, 14, 'neigh_op_rgt_2')
// (19, 15, 'neigh_op_bnr_2')
// (20, 13, 'neigh_op_top_2')
// (20, 14, 'local_g3_2')
// (20, 14, 'lutff_2/out')
// (20, 14, 'lutff_3/in_0')
// (20, 15, 'neigh_op_bot_2')
// (21, 13, 'neigh_op_tnl_2')
// (21, 14, 'neigh_op_lft_2')
// (21, 15, 'neigh_op_bnl_2')

wire n2715;
// (19, 13, 'neigh_op_tnr_3')
// (19, 14, 'neigh_op_rgt_3')
// (19, 15, 'neigh_op_bnr_3')
// (20, 13, 'neigh_op_top_3')
// (20, 14, 'lutff_3/out')
// (20, 15, 'local_g1_3')
// (20, 15, 'lutff_7/in_1')
// (20, 15, 'neigh_op_bot_3')
// (21, 13, 'neigh_op_tnl_3')
// (21, 14, 'neigh_op_lft_3')
// (21, 15, 'neigh_op_bnl_3')

reg n2716 = 0;
// (19, 13, 'neigh_op_tnr_4')
// (19, 14, 'neigh_op_rgt_4')
// (19, 14, 'sp4_r_v_b_40')
// (19, 15, 'neigh_op_bnr_4')
// (19, 15, 'sp4_r_v_b_29')
// (19, 16, 'sp4_r_v_b_16')
// (19, 17, 'sp4_r_v_b_5')
// (20, 13, 'neigh_op_top_4')
// (20, 13, 'sp4_h_r_5')
// (20, 13, 'sp4_v_t_40')
// (20, 14, 'lutff_4/out')
// (20, 14, 'sp4_v_b_40')
// (20, 15, 'neigh_op_bot_4')
// (20, 15, 'sp4_v_b_29')
// (20, 16, 'sp4_v_b_16')
// (20, 17, 'sp4_v_b_5')
// (21, 13, 'neigh_op_tnl_4')
// (21, 13, 'sp4_h_r_16')
// (21, 14, 'neigh_op_lft_4')
// (21, 15, 'neigh_op_bnl_4')
// (22, 13, 'local_g2_5')
// (22, 13, 'lutff_0/in_3')
// (22, 13, 'sp4_h_r_29')
// (23, 13, 'sp4_h_r_40')
// (24, 13, 'sp4_h_l_40')

reg n2717 = 0;
// (19, 13, 'neigh_op_tnr_5')
// (19, 14, 'neigh_op_rgt_5')
// (19, 15, 'neigh_op_bnr_5')
// (20, 11, 'sp4_r_v_b_46')
// (20, 12, 'sp4_r_v_b_35')
// (20, 13, 'neigh_op_top_5')
// (20, 13, 'sp4_r_v_b_22')
// (20, 14, 'lutff_5/out')
// (20, 14, 'sp4_r_v_b_11')
// (20, 15, 'neigh_op_bot_5')
// (21, 10, 'sp4_v_t_46')
// (21, 11, 'sp4_v_b_46')
// (21, 12, 'local_g2_3')
// (21, 12, 'lutff_5/in_0')
// (21, 12, 'sp4_v_b_35')
// (21, 13, 'neigh_op_tnl_5')
// (21, 13, 'sp4_v_b_22')
// (21, 14, 'neigh_op_lft_5')
// (21, 14, 'sp4_v_b_11')
// (21, 15, 'neigh_op_bnl_5')

reg n2718 = 0;
// (19, 13, 'neigh_op_tnr_6')
// (19, 14, 'neigh_op_rgt_6')
// (19, 15, 'neigh_op_bnr_6')
// (20, 13, 'neigh_op_top_6')
// (20, 13, 'sp4_r_v_b_40')
// (20, 14, 'lutff_6/out')
// (20, 14, 'sp4_r_v_b_29')
// (20, 15, 'neigh_op_bot_6')
// (20, 15, 'sp4_r_v_b_16')
// (20, 16, 'sp4_r_v_b_5')
// (21, 12, 'local_g1_5')
// (21, 12, 'lutff_2/in_2')
// (21, 12, 'sp4_h_r_5')
// (21, 12, 'sp4_v_t_40')
// (21, 13, 'neigh_op_tnl_6')
// (21, 13, 'sp4_v_b_40')
// (21, 14, 'neigh_op_lft_6')
// (21, 14, 'sp4_v_b_29')
// (21, 15, 'neigh_op_bnl_6')
// (21, 15, 'sp4_v_b_16')
// (21, 16, 'sp4_v_b_5')
// (22, 12, 'sp4_h_r_16')
// (23, 12, 'sp4_h_r_29')
// (24, 12, 'sp4_h_r_40')
// (25, 12, 'sp4_h_l_40')

wire n2719;
// (19, 13, 'neigh_op_tnr_7')
// (19, 14, 'neigh_op_rgt_7')
// (19, 15, 'neigh_op_bnr_7')
// (20, 13, 'neigh_op_top_7')
// (20, 14, 'local_g3_7')
// (20, 14, 'lutff_3/in_1')
// (20, 14, 'lutff_7/out')
// (20, 15, 'neigh_op_bot_7')
// (21, 13, 'neigh_op_tnl_7')
// (21, 14, 'neigh_op_lft_7')
// (21, 15, 'neigh_op_bnl_7')

wire n2720;
// (19, 13, 'sp4_r_v_b_37')
// (19, 14, 'sp4_r_v_b_24')
// (19, 15, 'sp4_r_v_b_13')
// (19, 16, 'sp4_r_v_b_0')
// (20, 12, 'sp4_h_r_0')
// (20, 12, 'sp4_v_t_37')
// (20, 13, 'local_g2_5')
// (20, 13, 'lutff_4/in_3')
// (20, 13, 'lutff_5/in_0')
// (20, 13, 'sp4_v_b_37')
// (20, 14, 'sp4_v_b_24')
// (20, 15, 'sp4_v_b_13')
// (20, 16, 'sp4_v_b_0')
// (21, 11, 'neigh_op_tnr_4')
// (21, 12, 'local_g2_4')
// (21, 12, 'lutff_5/in_3')
// (21, 12, 'neigh_op_rgt_4')
// (21, 12, 'sp4_h_r_13')
// (21, 13, 'neigh_op_bnr_4')
// (22, 11, 'neigh_op_top_4')
// (22, 12, 'lutff_4/out')
// (22, 12, 'sp4_h_r_24')
// (22, 13, 'local_g1_4')
// (22, 13, 'lutff_2/in_3')
// (22, 13, 'neigh_op_bot_4')
// (23, 11, 'neigh_op_tnl_4')
// (23, 12, 'neigh_op_lft_4')
// (23, 12, 'sp4_h_r_37')
// (23, 13, 'neigh_op_bnl_4')
// (24, 12, 'sp4_h_l_37')

reg n2721 = 0;
// (19, 14, 'neigh_op_tnr_1')
// (19, 15, 'neigh_op_rgt_1')
// (19, 16, 'neigh_op_bnr_1')
// (19, 16, 'sp4_r_v_b_39')
// (19, 17, 'sp4_r_v_b_26')
// (19, 18, 'sp4_r_v_b_15')
// (19, 19, 'sp4_r_v_b_2')
// (20, 14, 'neigh_op_top_1')
// (20, 15, 'lutff_1/out')
// (20, 15, 'sp4_h_r_2')
// (20, 15, 'sp4_v_t_39')
// (20, 16, 'neigh_op_bot_1')
// (20, 16, 'sp4_v_b_39')
// (20, 17, 'sp4_v_b_26')
// (20, 18, 'local_g1_7')
// (20, 18, 'lutff_3/in_3')
// (20, 18, 'sp4_v_b_15')
// (20, 19, 'sp4_v_b_2')
// (21, 14, 'neigh_op_tnl_1')
// (21, 15, 'neigh_op_lft_1')
// (21, 15, 'sp4_h_r_15')
// (21, 16, 'neigh_op_bnl_1')
// (22, 15, 'sp4_h_r_26')
// (23, 15, 'sp4_h_r_39')
// (24, 15, 'sp4_h_l_39')

wire n2722;
// (19, 14, 'neigh_op_tnr_5')
// (19, 15, 'neigh_op_rgt_5')
// (19, 16, 'neigh_op_bnr_5')
// (20, 14, 'neigh_op_top_5')
// (20, 15, 'local_g0_2')
// (20, 15, 'lutff_5/out')
// (20, 15, 'lutff_global/cen')
// (20, 15, 'sp4_h_r_10')
// (20, 16, 'neigh_op_bot_5')
// (21, 14, 'neigh_op_tnl_5')
// (21, 15, 'neigh_op_lft_5')
// (21, 15, 'sp4_h_r_23')
// (21, 16, 'neigh_op_bnl_5')
// (22, 15, 'sp4_h_r_34')
// (23, 15, 'sp4_h_r_47')
// (24, 15, 'sp4_h_l_47')

reg n2723 = 0;
// (19, 15, 'neigh_op_tnr_3')
// (19, 16, 'neigh_op_rgt_3')
// (19, 17, 'neigh_op_bnr_3')
// (20, 15, 'neigh_op_top_3')
// (20, 16, 'lutff_3/out')
// (20, 17, 'neigh_op_bot_3')
// (21, 15, 'neigh_op_tnl_3')
// (21, 16, 'local_g1_3')
// (21, 16, 'lutff_4/in_2')
// (21, 16, 'neigh_op_lft_3')
// (21, 17, 'neigh_op_bnl_3')

wire n2724;
// (19, 16, 'neigh_op_tnr_0')
// (19, 17, 'neigh_op_rgt_0')
// (19, 18, 'neigh_op_bnr_0')
// (20, 16, 'neigh_op_top_0')
// (20, 17, 'lutff_0/out')
// (20, 18, 'local_g0_0')
// (20, 18, 'lutff_1/in_1')
// (20, 18, 'neigh_op_bot_0')
// (21, 16, 'neigh_op_tnl_0')
// (21, 17, 'neigh_op_lft_0')
// (21, 18, 'neigh_op_bnl_0')

reg n2725 = 0;
// (19, 16, 'neigh_op_tnr_4')
// (19, 17, 'neigh_op_rgt_4')
// (19, 18, 'neigh_op_bnr_4')
// (20, 16, 'neigh_op_top_4')
// (20, 17, 'lutff_4/out')
// (20, 18, 'local_g0_4')
// (20, 18, 'lutff_4/in_2')
// (20, 18, 'neigh_op_bot_4')
// (21, 16, 'neigh_op_tnl_4')
// (21, 17, 'neigh_op_lft_4')
// (21, 18, 'neigh_op_bnl_4')

wire n2726;
// (19, 16, 'neigh_op_tnr_5')
// (19, 17, 'neigh_op_rgt_5')
// (19, 18, 'neigh_op_bnr_5')
// (20, 16, 'neigh_op_top_5')
// (20, 17, 'local_g0_5')
// (20, 17, 'lutff_0/in_3')
// (20, 17, 'lutff_5/out')
// (20, 18, 'neigh_op_bot_5')
// (21, 16, 'neigh_op_tnl_5')
// (21, 17, 'neigh_op_lft_5')
// (21, 18, 'neigh_op_bnl_5')

wire n2727;
// (19, 16, 'sp4_r_v_b_46')
// (19, 17, 'sp4_r_v_b_35')
// (19, 18, 'sp4_r_v_b_22')
// (19, 19, 'sp4_r_v_b_11')
// (19, 20, 'sp4_r_v_b_38')
// (19, 21, 'neigh_op_tnr_7')
// (19, 21, 'sp4_r_v_b_27')
// (19, 22, 'neigh_op_rgt_7')
// (19, 22, 'sp4_r_v_b_14')
// (19, 23, 'neigh_op_bnr_7')
// (19, 23, 'sp4_r_v_b_3')
// (20, 15, 'sp4_v_t_46')
// (20, 16, 'sp4_v_b_46')
// (20, 17, 'local_g3_3')
// (20, 17, 'lutff_5/in_3')
// (20, 17, 'sp4_v_b_35')
// (20, 18, 'sp4_v_b_22')
// (20, 19, 'sp4_v_b_11')
// (20, 19, 'sp4_v_t_38')
// (20, 20, 'sp4_v_b_38')
// (20, 21, 'neigh_op_top_7')
// (20, 21, 'sp4_v_b_27')
// (20, 22, 'lutff_7/out')
// (20, 22, 'sp4_v_b_14')
// (20, 23, 'neigh_op_bot_7')
// (20, 23, 'sp4_v_b_3')
// (21, 21, 'neigh_op_tnl_7')
// (21, 22, 'neigh_op_lft_7')
// (21, 23, 'neigh_op_bnl_7')

reg n2728 = 0;
// (19, 16, 'sp4_r_v_b_47')
// (19, 17, 'sp4_r_v_b_34')
// (19, 18, 'sp4_r_v_b_23')
// (19, 19, 'sp4_r_v_b_10')
// (20, 15, 'sp4_v_t_47')
// (20, 16, 'sp4_v_b_47')
// (20, 17, 'sp4_v_b_34')
// (20, 18, 'local_g0_7')
// (20, 18, 'lutff_4/in_1')
// (20, 18, 'sp4_v_b_23')
// (20, 19, 'sp4_h_r_10')
// (20, 19, 'sp4_v_b_10')
// (21, 18, 'neigh_op_tnr_1')
// (21, 19, 'neigh_op_rgt_1')
// (21, 19, 'sp4_h_r_23')
// (21, 20, 'neigh_op_bnr_1')
// (22, 18, 'neigh_op_top_1')
// (22, 19, 'lutff_1/out')
// (22, 19, 'sp4_h_r_34')
// (22, 20, 'neigh_op_bot_1')
// (23, 18, 'neigh_op_tnl_1')
// (23, 19, 'neigh_op_lft_1')
// (23, 19, 'sp4_h_r_47')
// (23, 20, 'neigh_op_bnl_1')
// (24, 19, 'sp4_h_l_47')

wire n2729;
// (19, 17, 'neigh_op_tnr_1')
// (19, 18, 'neigh_op_rgt_1')
// (19, 19, 'neigh_op_bnr_1')
// (20, 17, 'neigh_op_top_1')
// (20, 18, 'local_g0_1')
// (20, 18, 'lutff_0/in_1')
// (20, 18, 'lutff_1/out')
// (20, 19, 'neigh_op_bot_1')
// (21, 17, 'neigh_op_tnl_1')
// (21, 18, 'neigh_op_lft_1')
// (21, 19, 'neigh_op_bnl_1')

wire n2730;
// (19, 17, 'neigh_op_tnr_3')
// (19, 18, 'neigh_op_rgt_3')
// (19, 19, 'neigh_op_bnr_3')
// (20, 17, 'neigh_op_top_3')
// (20, 18, 'local_g0_3')
// (20, 18, 'lutff_3/out')
// (20, 18, 'lutff_6/in_1')
// (20, 19, 'neigh_op_bot_3')
// (21, 17, 'neigh_op_tnl_3')
// (21, 18, 'neigh_op_lft_3')
// (21, 19, 'neigh_op_bnl_3')

wire n2731;
// (19, 17, 'neigh_op_tnr_4')
// (19, 18, 'neigh_op_rgt_4')
// (19, 19, 'neigh_op_bnr_4')
// (20, 17, 'neigh_op_top_4')
// (20, 18, 'local_g2_4')
// (20, 18, 'lutff_4/out')
// (20, 18, 'lutff_7/in_3')
// (20, 19, 'neigh_op_bot_4')
// (21, 17, 'neigh_op_tnl_4')
// (21, 18, 'neigh_op_lft_4')
// (21, 19, 'neigh_op_bnl_4')

wire n2732;
// (19, 17, 'neigh_op_tnr_5')
// (19, 18, 'neigh_op_rgt_5')
// (19, 19, 'neigh_op_bnr_5')
// (20, 17, 'neigh_op_top_5')
// (20, 18, 'local_g0_2')
// (20, 18, 'lutff_5/out')
// (20, 18, 'lutff_global/cen')
// (20, 18, 'sp4_h_r_10')
// (20, 19, 'neigh_op_bot_5')
// (21, 17, 'neigh_op_tnl_5')
// (21, 18, 'neigh_op_lft_5')
// (21, 18, 'sp4_h_r_23')
// (21, 19, 'neigh_op_bnl_5')
// (22, 18, 'sp4_h_r_34')
// (23, 18, 'sp4_h_r_47')
// (24, 18, 'sp4_h_l_47')

wire n2733;
// (19, 17, 'neigh_op_tnr_6')
// (19, 18, 'neigh_op_rgt_6')
// (19, 19, 'neigh_op_bnr_6')
// (20, 17, 'neigh_op_top_6')
// (20, 18, 'local_g1_6')
// (20, 18, 'lutff_1/in_2')
// (20, 18, 'lutff_6/out')
// (20, 19, 'neigh_op_bot_6')
// (21, 17, 'neigh_op_tnl_6')
// (21, 18, 'neigh_op_lft_6')
// (21, 19, 'neigh_op_bnl_6')

wire n2734;
// (19, 17, 'neigh_op_tnr_7')
// (19, 18, 'neigh_op_rgt_7')
// (19, 19, 'neigh_op_bnr_7')
// (20, 17, 'neigh_op_top_7')
// (20, 18, 'lutff_7/out')
// (20, 19, 'local_g0_7')
// (20, 19, 'lutff_1/in_0')
// (20, 19, 'neigh_op_bot_7')
// (21, 17, 'neigh_op_tnl_7')
// (21, 18, 'neigh_op_lft_7')
// (21, 19, 'neigh_op_bnl_7')

wire n2735;
// (19, 17, 'sp4_h_r_10')
// (20, 16, 'neigh_op_tnr_1')
// (20, 17, 'neigh_op_rgt_1')
// (20, 17, 'sp4_h_r_23')
// (20, 18, 'neigh_op_bnr_1')
// (21, 16, 'neigh_op_top_1')
// (21, 17, 'local_g2_2')
// (21, 17, 'lutff_1/out')
// (21, 17, 'lutff_global/cen')
// (21, 17, 'sp4_h_r_34')
// (21, 18, 'neigh_op_bot_1')
// (22, 16, 'neigh_op_tnl_1')
// (22, 17, 'neigh_op_lft_1')
// (22, 17, 'sp4_h_r_47')
// (22, 18, 'neigh_op_bnl_1')
// (23, 17, 'sp4_h_l_47')

wire n2736;
// (19, 17, 'sp4_h_r_3')
// (20, 17, 'sp4_h_r_14')
// (21, 16, 'neigh_op_tnr_3')
// (21, 17, 'neigh_op_rgt_3')
// (21, 17, 'sp4_h_r_27')
// (21, 18, 'neigh_op_bnr_3')
// (22, 16, 'neigh_op_top_3')
// (22, 17, 'lutff_3/out')
// (22, 17, 'sp4_h_r_38')
// (22, 18, 'neigh_op_bot_3')
// (23, 16, 'neigh_op_tnl_3')
// (23, 17, 'neigh_op_lft_3')
// (23, 17, 'sp4_h_l_38')
// (23, 17, 'sp4_h_r_6')
// (23, 18, 'neigh_op_bnl_3')
// (24, 17, 'local_g1_3')
// (24, 17, 'lutff_global/cen')
// (24, 17, 'sp4_h_r_19')
// (25, 17, 'sp4_h_r_30')

wire n2737;
// (19, 17, 'sp4_h_r_9')
// (20, 17, 'sp4_h_r_20')
// (21, 16, 'neigh_op_tnr_6')
// (21, 17, 'neigh_op_rgt_6')
// (21, 17, 'sp4_h_r_33')
// (21, 18, 'neigh_op_bnr_6')
// (22, 14, 'sp4_r_v_b_38')
// (22, 15, 'sp4_r_v_b_27')
// (22, 16, 'neigh_op_top_6')
// (22, 16, 'sp4_r_v_b_14')
// (22, 17, 'local_g1_3')
// (22, 17, 'lutff_6/out')
// (22, 17, 'lutff_global/cen')
// (22, 17, 'sp4_h_r_44')
// (22, 17, 'sp4_r_v_b_3')
// (22, 18, 'neigh_op_bot_6')
// (23, 13, 'sp4_v_t_38')
// (23, 14, 'sp4_v_b_38')
// (23, 15, 'sp4_v_b_27')
// (23, 16, 'neigh_op_tnl_6')
// (23, 16, 'sp4_v_b_14')
// (23, 17, 'neigh_op_lft_6')
// (23, 17, 'sp4_h_l_44')
// (23, 17, 'sp4_v_b_3')
// (23, 18, 'neigh_op_bnl_6')

wire n2738;
// (19, 17, 'sp4_r_v_b_45')
// (19, 18, 'sp4_r_v_b_32')
// (19, 19, 'neigh_op_tnr_4')
// (19, 19, 'sp4_r_v_b_21')
// (19, 20, 'neigh_op_rgt_4')
// (19, 20, 'sp4_r_v_b_8')
// (19, 21, 'neigh_op_bnr_4')
// (20, 16, 'sp4_v_t_45')
// (20, 17, 'sp4_v_b_45')
// (20, 18, 'sp4_v_b_32')
// (20, 19, 'neigh_op_top_4')
// (20, 19, 'sp4_v_b_21')
// (20, 20, 'local_g0_2')
// (20, 20, 'lutff_4/out')
// (20, 20, 'lutff_global/cen')
// (20, 20, 'sp4_h_r_2')
// (20, 20, 'sp4_v_b_8')
// (20, 21, 'neigh_op_bot_4')
// (21, 19, 'neigh_op_tnl_4')
// (21, 20, 'neigh_op_lft_4')
// (21, 20, 'sp4_h_r_15')
// (21, 21, 'neigh_op_bnl_4')
// (22, 20, 'sp4_h_r_26')
// (23, 20, 'sp4_h_r_39')
// (24, 20, 'sp4_h_l_39')

wire n2739;
// (19, 18, 'neigh_op_tnr_1')
// (19, 19, 'neigh_op_rgt_1')
// (19, 20, 'neigh_op_bnr_1')
// (20, 18, 'local_g1_1')
// (20, 18, 'lutff_0/in_2')
// (20, 18, 'neigh_op_top_1')
// (20, 19, 'lutff_1/out')
// (20, 20, 'neigh_op_bot_1')
// (21, 18, 'neigh_op_tnl_1')
// (21, 19, 'neigh_op_lft_1')
// (21, 20, 'neigh_op_bnl_1')

wire n2740;
// (19, 19, 'neigh_op_tnr_0')
// (19, 19, 'sp4_r_v_b_45')
// (19, 20, 'neigh_op_rgt_0')
// (19, 20, 'sp4_r_v_b_32')
// (19, 21, 'neigh_op_bnr_0')
// (19, 21, 'sp4_r_v_b_21')
// (19, 22, 'sp4_r_v_b_8')
// (20, 18, 'sp4_v_t_45')
// (20, 19, 'neigh_op_top_0')
// (20, 19, 'sp4_v_b_45')
// (20, 20, 'lutff_0/out')
// (20, 20, 'sp4_v_b_32')
// (20, 21, 'neigh_op_bot_0')
// (20, 21, 'sp4_v_b_21')
// (20, 22, 'local_g0_2')
// (20, 22, 'lutff_global/cen')
// (20, 22, 'sp4_h_r_2')
// (20, 22, 'sp4_v_b_8')
// (21, 19, 'neigh_op_tnl_0')
// (21, 20, 'neigh_op_lft_0')
// (21, 21, 'neigh_op_bnl_0')
// (21, 22, 'sp4_h_r_15')
// (22, 22, 'sp4_h_r_26')
// (23, 22, 'sp4_h_r_39')
// (24, 22, 'sp4_h_l_39')

wire n2741;
// (19, 19, 'neigh_op_tnr_1')
// (19, 20, 'neigh_op_rgt_1')
// (19, 21, 'neigh_op_bnr_1')
// (20, 19, 'local_g1_1')
// (20, 19, 'lutff_1/in_1')
// (20, 19, 'neigh_op_top_1')
// (20, 20, 'lutff_1/out')
// (20, 21, 'neigh_op_bot_1')
// (21, 19, 'neigh_op_tnl_1')
// (21, 20, 'neigh_op_lft_1')
// (21, 21, 'neigh_op_bnl_1')

reg n2742 = 0;
// (19, 19, 'neigh_op_tnr_2')
// (19, 20, 'neigh_op_rgt_2')
// (19, 21, 'neigh_op_bnr_2')
// (20, 19, 'neigh_op_top_2')
// (20, 20, 'local_g2_2')
// (20, 20, 'lutff_2/out')
// (20, 20, 'lutff_5/in_3')
// (20, 21, 'neigh_op_bot_2')
// (21, 19, 'neigh_op_tnl_2')
// (21, 20, 'neigh_op_lft_2')
// (21, 21, 'neigh_op_bnl_2')

wire n2743;
// (19, 19, 'neigh_op_tnr_3')
// (19, 20, 'neigh_op_rgt_3')
// (19, 21, 'neigh_op_bnr_3')
// (20, 19, 'local_g0_3')
// (20, 19, 'lutff_1/in_2')
// (20, 19, 'neigh_op_top_3')
// (20, 20, 'lutff_3/out')
// (20, 21, 'neigh_op_bot_3')
// (21, 19, 'neigh_op_tnl_3')
// (21, 20, 'neigh_op_lft_3')
// (21, 21, 'neigh_op_bnl_3')

wire n2744;
// (19, 19, 'neigh_op_tnr_5')
// (19, 20, 'neigh_op_rgt_5')
// (19, 21, 'neigh_op_bnr_5')
// (20, 19, 'neigh_op_top_5')
// (20, 20, 'local_g0_5')
// (20, 20, 'lutff_5/out')
// (20, 20, 'lutff_7/in_2')
// (20, 21, 'neigh_op_bot_5')
// (21, 19, 'neigh_op_tnl_5')
// (21, 20, 'neigh_op_lft_5')
// (21, 21, 'neigh_op_bnl_5')

wire n2745;
// (19, 19, 'neigh_op_tnr_6')
// (19, 20, 'neigh_op_rgt_6')
// (19, 20, 'sp4_r_v_b_44')
// (19, 21, 'neigh_op_bnr_6')
// (19, 21, 'sp4_r_v_b_33')
// (19, 22, 'sp4_r_v_b_20')
// (19, 23, 'sp4_r_v_b_9')
// (20, 19, 'local_g0_2')
// (20, 19, 'lutff_global/cen')
// (20, 19, 'neigh_op_top_6')
// (20, 19, 'sp4_h_r_2')
// (20, 19, 'sp4_v_t_44')
// (20, 20, 'lutff_6/out')
// (20, 20, 'sp4_v_b_44')
// (20, 21, 'neigh_op_bot_6')
// (20, 21, 'sp4_v_b_33')
// (20, 22, 'sp4_v_b_20')
// (20, 23, 'sp4_v_b_9')
// (21, 19, 'neigh_op_tnl_6')
// (21, 19, 'sp4_h_r_15')
// (21, 20, 'neigh_op_lft_6')
// (21, 21, 'neigh_op_bnl_6')
// (22, 19, 'sp4_h_r_26')
// (23, 19, 'sp4_h_r_39')
// (24, 19, 'sp4_h_l_39')

wire n2746;
// (19, 19, 'neigh_op_tnr_7')
// (19, 20, 'neigh_op_rgt_7')
// (19, 21, 'neigh_op_bnr_7')
// (20, 18, 'sp4_r_v_b_39')
// (20, 19, 'neigh_op_top_7')
// (20, 19, 'sp4_r_v_b_26')
// (20, 20, 'lutff_7/out')
// (20, 20, 'sp4_r_v_b_15')
// (20, 21, 'neigh_op_bot_7')
// (20, 21, 'sp4_r_v_b_2')
// (21, 17, 'sp4_v_t_39')
// (21, 18, 'local_g3_7')
// (21, 18, 'lutff_3/in_3')
// (21, 18, 'sp4_v_b_39')
// (21, 19, 'neigh_op_tnl_7')
// (21, 19, 'sp4_v_b_26')
// (21, 20, 'neigh_op_lft_7')
// (21, 20, 'sp4_v_b_15')
// (21, 21, 'neigh_op_bnl_7')
// (21, 21, 'sp4_v_b_2')

wire n2747;
// (19, 19, 'sp4_h_r_9')
// (20, 19, 'sp4_h_r_20')
// (21, 18, 'neigh_op_tnr_6')
// (21, 19, 'neigh_op_rgt_6')
// (21, 19, 'sp4_h_r_33')
// (21, 20, 'neigh_op_bnr_6')
// (22, 16, 'sp4_r_v_b_38')
// (22, 17, 'sp4_r_v_b_27')
// (22, 18, 'neigh_op_top_6')
// (22, 18, 'sp4_r_v_b_14')
// (22, 19, 'local_g1_3')
// (22, 19, 'lutff_6/out')
// (22, 19, 'lutff_global/cen')
// (22, 19, 'sp4_h_r_44')
// (22, 19, 'sp4_r_v_b_3')
// (22, 20, 'neigh_op_bot_6')
// (23, 15, 'sp4_v_t_38')
// (23, 16, 'sp4_v_b_38')
// (23, 17, 'sp4_v_b_27')
// (23, 18, 'neigh_op_tnl_6')
// (23, 18, 'sp4_v_b_14')
// (23, 19, 'neigh_op_lft_6')
// (23, 19, 'sp4_h_l_44')
// (23, 19, 'sp4_v_b_3')
// (23, 20, 'neigh_op_bnl_6')

reg n2748 = 0;
// (19, 20, 'neigh_op_tnr_2')
// (19, 21, 'neigh_op_rgt_2')
// (19, 22, 'neigh_op_bnr_2')
// (20, 20, 'neigh_op_top_2')
// (20, 21, 'local_g1_2')
// (20, 21, 'lutff_2/out')
// (20, 21, 'lutff_3/in_2')
// (20, 22, 'neigh_op_bot_2')
// (21, 20, 'neigh_op_tnl_2')
// (21, 21, 'neigh_op_lft_2')
// (21, 22, 'neigh_op_bnl_2')

wire n2749;
// (19, 20, 'neigh_op_tnr_3')
// (19, 21, 'neigh_op_rgt_3')
// (19, 22, 'neigh_op_bnr_3')
// (20, 20, 'neigh_op_top_3')
// (20, 21, 'local_g3_3')
// (20, 21, 'lutff_3/out')
// (20, 21, 'lutff_7/in_1')
// (20, 22, 'neigh_op_bot_3')
// (21, 20, 'neigh_op_tnl_3')
// (21, 21, 'neigh_op_lft_3')
// (21, 22, 'neigh_op_bnl_3')

wire n2750;
// (19, 20, 'neigh_op_tnr_7')
// (19, 21, 'neigh_op_rgt_7')
// (19, 22, 'neigh_op_bnr_7')
// (20, 20, 'local_g1_7')
// (20, 20, 'lutff_1/in_1')
// (20, 20, 'neigh_op_top_7')
// (20, 21, 'lutff_7/out')
// (20, 22, 'neigh_op_bot_7')
// (21, 20, 'neigh_op_tnl_7')
// (21, 21, 'neigh_op_lft_7')
// (21, 22, 'neigh_op_bnl_7')

wire n2751;
// (19, 20, 'sp4_h_r_5')
// (20, 20, 'sp4_h_r_16')
// (21, 19, 'neigh_op_tnr_4')
// (21, 20, 'neigh_op_rgt_4')
// (21, 20, 'sp4_h_r_29')
// (21, 21, 'neigh_op_bnr_4')
// (22, 19, 'neigh_op_top_4')
// (22, 20, 'lutff_4/out')
// (22, 20, 'sp4_h_r_40')
// (22, 21, 'neigh_op_bot_4')
// (22, 21, 'sp4_r_v_b_42')
// (22, 22, 'sp4_r_v_b_31')
// (22, 23, 'sp4_r_v_b_18')
// (22, 24, 'sp4_r_v_b_7')
// (23, 19, 'neigh_op_tnl_4')
// (23, 20, 'neigh_op_lft_4')
// (23, 20, 'sp4_h_l_40')
// (23, 20, 'sp4_h_r_1')
// (23, 20, 'sp4_v_t_42')
// (23, 21, 'local_g2_2')
// (23, 21, 'lutff_global/cen')
// (23, 21, 'neigh_op_bnl_4')
// (23, 21, 'sp4_v_b_42')
// (23, 22, 'sp4_v_b_31')
// (23, 23, 'sp4_v_b_18')
// (23, 24, 'sp4_v_b_7')
// (24, 20, 'sp4_h_r_12')
// (25, 20, 'sp4_h_r_25')

reg n2752 = 0;
// (19, 21, 'neigh_op_tnr_0')
// (19, 22, 'neigh_op_rgt_0')
// (19, 23, 'neigh_op_bnr_0')
// (20, 21, 'neigh_op_top_0')
// (20, 22, 'local_g2_0')
// (20, 22, 'lutff_0/out')
// (20, 22, 'lutff_7/in_3')
// (20, 23, 'neigh_op_bot_0')
// (21, 21, 'neigh_op_tnl_0')
// (21, 22, 'neigh_op_lft_0')
// (21, 23, 'neigh_op_bnl_0')

wire n2753;
// (19, 21, 'neigh_op_tnr_5')
// (19, 22, 'neigh_op_rgt_5')
// (19, 23, 'neigh_op_bnr_5')
// (20, 21, 'local_g0_5')
// (20, 21, 'lutff_7/in_2')
// (20, 21, 'neigh_op_top_5')
// (20, 22, 'lutff_5/out')
// (20, 23, 'neigh_op_bot_5')
// (21, 21, 'neigh_op_tnl_5')
// (21, 22, 'neigh_op_lft_5')
// (21, 23, 'neigh_op_bnl_5')

wire n2754;
// (19, 22, 'neigh_op_tnr_3')
// (19, 23, 'neigh_op_rgt_3')
// (19, 24, 'neigh_op_bnr_3')
// (20, 22, 'neigh_op_top_3')
// (20, 23, 'local_g3_3')
// (20, 23, 'lutff_3/out')
// (20, 23, 'lutff_global/cen')
// (20, 24, 'neigh_op_bot_3')
// (21, 22, 'neigh_op_tnl_3')
// (21, 23, 'neigh_op_lft_3')
// (21, 24, 'neigh_op_bnl_3')

reg n2755 = 0;
// (19, 22, 'sp4_h_r_3')
// (20, 22, 'local_g1_6')
// (20, 22, 'lutff_5/in_0')
// (20, 22, 'sp4_h_r_14')
// (21, 22, 'sp4_h_r_27')
// (22, 21, 'neigh_op_tnr_0')
// (22, 22, 'neigh_op_rgt_0')
// (22, 22, 'sp4_h_r_38')
// (22, 23, 'neigh_op_bnr_0')
// (23, 21, 'neigh_op_top_0')
// (23, 22, 'lutff_0/out')
// (23, 22, 'sp4_h_l_38')
// (23, 22, 'sp4_h_r_0')
// (23, 23, 'neigh_op_bot_0')
// (24, 21, 'neigh_op_tnl_0')
// (24, 22, 'neigh_op_lft_0')
// (24, 22, 'sp4_h_r_13')
// (24, 23, 'neigh_op_bnl_0')
// (25, 22, 'sp4_h_r_24')

wire n2756;
// (20, 0, 'logic_op_tnr_0')
// (20, 1, 'neigh_op_rgt_0')
// (20, 2, 'neigh_op_bnr_0')
// (21, 0, 'logic_op_top_0')
// (21, 1, 'lutff_0/out')
// (21, 1, 'sp4_r_v_b_33')
// (21, 2, 'local_g1_0')
// (21, 2, 'lutff_0/in_3')
// (21, 2, 'lutff_5/in_0')
// (21, 2, 'neigh_op_bot_0')
// (21, 2, 'sp4_r_v_b_20')
// (21, 3, 'sp4_r_v_b_9')
// (22, 0, 'logic_op_tnl_0')
// (22, 0, 'span4_vert_33')
// (22, 1, 'neigh_op_lft_0')
// (22, 1, 'sp4_v_b_33')
// (22, 2, 'neigh_op_bnl_0')
// (22, 2, 'sp4_v_b_20')
// (22, 3, 'local_g0_1')
// (22, 3, 'local_g1_1')
// (22, 3, 'lutff_2/in_1')
// (22, 3, 'lutff_4/in_0')
// (22, 3, 'lutff_6/in_0')
// (22, 3, 'sp4_v_b_9')

wire n2757;
// (20, 0, 'logic_op_tnr_5')
// (20, 1, 'neigh_op_rgt_5')
// (20, 1, 'sp4_r_v_b_26')
// (20, 2, 'neigh_op_bnr_5')
// (20, 2, 'sp4_r_v_b_15')
// (20, 3, 'sp4_r_v_b_2')
// (21, 0, 'logic_op_top_5')
// (21, 0, 'span4_vert_26')
// (21, 1, 'local_g3_5')
// (21, 1, 'lutff_5/out')
// (21, 1, 'lutff_global/s_r')
// (21, 1, 'sp4_r_v_b_27')
// (21, 1, 'sp4_v_b_26')
// (21, 2, 'local_g0_5')
// (21, 2, 'lutff_4/in_3')
// (21, 2, 'lutff_5/in_2')
// (21, 2, 'neigh_op_bot_5')
// (21, 2, 'sp4_r_v_b_14')
// (21, 2, 'sp4_v_b_15')
// (21, 3, 'sp4_h_r_8')
// (21, 3, 'sp4_r_v_b_3')
// (21, 3, 'sp4_v_b_2')
// (22, 0, 'logic_op_tnl_5')
// (22, 0, 'span4_vert_27')
// (22, 1, 'neigh_op_lft_5')
// (22, 1, 'sp4_v_b_27')
// (22, 2, 'local_g0_6')
// (22, 2, 'lutff_0/in_0')
// (22, 2, 'lutff_1/in_3')
// (22, 2, 'lutff_2/in_2')
// (22, 2, 'lutff_6/in_2')
// (22, 2, 'neigh_op_bnl_5')
// (22, 2, 'sp4_v_b_14')
// (22, 3, 'local_g1_5')
// (22, 3, 'lutff_global/s_r')
// (22, 3, 'sp4_h_r_21')
// (22, 3, 'sp4_v_b_3')
// (23, 3, 'sp4_h_r_32')
// (24, 3, 'sp4_h_r_45')
// (25, 3, 'sp4_h_l_45')

wire n2758;
// (20, 1, 'local_g3_5')
// (20, 1, 'lutff_global/s_r')
// (20, 1, 'neigh_op_tnr_5')
// (20, 2, 'neigh_op_rgt_5')
// (20, 3, 'neigh_op_bnr_5')
// (21, 1, 'neigh_op_top_5')
// (21, 2, 'local_g2_5')
// (21, 2, 'lutff_3/in_0')
// (21, 2, 'lutff_5/out')
// (21, 3, 'neigh_op_bot_5')
// (22, 1, 'neigh_op_tnl_5')
// (22, 2, 'neigh_op_lft_5')
// (22, 3, 'neigh_op_bnl_5')

wire n2759;
// (20, 1, 'lutff_1/cout')
// (20, 1, 'lutff_2/in_3')

wire n2760;
// (20, 1, 'lutff_2/cout')
// (20, 1, 'lutff_3/in_3')

wire n2761;
// (20, 1, 'neigh_op_tnr_0')
// (20, 1, 'sp4_r_v_b_16')
// (20, 2, 'neigh_op_rgt_0')
// (20, 2, 'sp4_r_v_b_5')
// (20, 3, 'neigh_op_bnr_0')
// (21, 0, 'span4_vert_16')
// (21, 1, 'neigh_op_top_0')
// (21, 1, 'sp4_v_b_16')
// (21, 2, 'local_g1_5')
// (21, 2, 'lutff_0/out')
// (21, 2, 'lutff_global/s_r')
// (21, 2, 'sp4_h_r_0')
// (21, 2, 'sp4_v_b_5')
// (21, 3, 'neigh_op_bot_0')
// (22, 1, 'neigh_op_tnl_0')
// (22, 2, 'neigh_op_lft_0')
// (22, 2, 'sp4_h_r_13')
// (22, 3, 'neigh_op_bnl_0')
// (23, 2, 'sp4_h_r_24')
// (24, 2, 'sp4_h_r_37')
// (25, 2, 'sp4_h_l_37')

reg n2762 = 0;
// (20, 2, 'neigh_op_tnr_2')
// (20, 3, 'neigh_op_rgt_2')
// (20, 4, 'neigh_op_bnr_2')
// (21, 2, 'neigh_op_top_2')
// (21, 3, 'local_g1_2')
// (21, 3, 'lutff_2/in_1')
// (21, 3, 'lutff_2/out')
// (21, 4, 'neigh_op_bot_2')
// (22, 2, 'neigh_op_tnl_2')
// (22, 3, 'local_g0_2')
// (22, 3, 'lutff_5/in_3')
// (22, 3, 'neigh_op_lft_2')
// (22, 4, 'neigh_op_bnl_2')

reg n2763 = 0;
// (20, 2, 'neigh_op_tnr_3')
// (20, 3, 'neigh_op_rgt_3')
// (20, 4, 'neigh_op_bnr_3')
// (21, 1, 'sp4_r_v_b_47')
// (21, 2, 'neigh_op_top_3')
// (21, 2, 'sp4_r_v_b_34')
// (21, 3, 'local_g1_3')
// (21, 3, 'lutff_3/in_1')
// (21, 3, 'lutff_3/out')
// (21, 3, 'sp4_r_v_b_23')
// (21, 4, 'neigh_op_bot_3')
// (21, 4, 'sp4_r_v_b_10')
// (22, 0, 'span4_vert_47')
// (22, 1, 'sp4_v_b_47')
// (22, 2, 'neigh_op_tnl_3')
// (22, 2, 'sp4_v_b_34')
// (22, 3, 'local_g1_7')
// (22, 3, 'lutff_5/in_1')
// (22, 3, 'neigh_op_lft_3')
// (22, 3, 'sp4_v_b_23')
// (22, 4, 'neigh_op_bnl_3')
// (22, 4, 'sp4_v_b_10')

reg n2764 = 0;
// (20, 2, 'neigh_op_tnr_4')
// (20, 3, 'neigh_op_rgt_4')
// (20, 4, 'neigh_op_bnr_4')
// (21, 2, 'neigh_op_top_4')
// (21, 3, 'local_g3_4')
// (21, 3, 'lutff_4/in_1')
// (21, 3, 'lutff_4/out')
// (21, 4, 'neigh_op_bot_4')
// (22, 2, 'neigh_op_tnl_4')
// (22, 3, 'neigh_op_lft_4')
// (22, 4, 'local_g3_4')
// (22, 4, 'lutff_5/in_2')
// (22, 4, 'neigh_op_bnl_4')

reg n2765 = 0;
// (20, 2, 'neigh_op_tnr_5')
// (20, 3, 'neigh_op_rgt_5')
// (20, 4, 'neigh_op_bnr_5')
// (21, 2, 'neigh_op_top_5')
// (21, 3, 'local_g1_5')
// (21, 3, 'lutff_5/in_1')
// (21, 3, 'lutff_5/out')
// (21, 4, 'neigh_op_bot_5')
// (22, 2, 'neigh_op_tnl_5')
// (22, 3, 'local_g0_5')
// (22, 3, 'lutff_5/in_2')
// (22, 3, 'neigh_op_lft_5')
// (22, 4, 'neigh_op_bnl_5')

reg n2766 = 0;
// (20, 2, 'neigh_op_tnr_6')
// (20, 3, 'neigh_op_rgt_6')
// (20, 4, 'neigh_op_bnr_6')
// (21, 2, 'neigh_op_top_6')
// (21, 3, 'local_g2_6')
// (21, 3, 'lutff_6/in_2')
// (21, 3, 'lutff_6/out')
// (21, 4, 'neigh_op_bot_6')
// (22, 2, 'neigh_op_tnl_6')
// (22, 3, 'local_g1_6')
// (22, 3, 'lutff_7/in_0')
// (22, 3, 'neigh_op_lft_6')
// (22, 4, 'neigh_op_bnl_6')

reg n2767 = 0;
// (20, 2, 'neigh_op_tnr_7')
// (20, 3, 'neigh_op_rgt_7')
// (20, 4, 'neigh_op_bnr_7')
// (21, 2, 'neigh_op_top_7')
// (21, 3, 'local_g2_7')
// (21, 3, 'lutff_7/in_2')
// (21, 3, 'lutff_7/out')
// (21, 4, 'neigh_op_bot_7')
// (22, 2, 'neigh_op_tnl_7')
// (22, 3, 'local_g0_7')
// (22, 3, 'lutff_7/in_2')
// (22, 3, 'neigh_op_lft_7')
// (22, 4, 'neigh_op_bnl_7')

reg n2768 = 0;
// (20, 3, 'neigh_op_tnr_0')
// (20, 4, 'local_g3_0')
// (20, 4, 'lutff_7/in_2')
// (20, 4, 'neigh_op_rgt_0')
// (20, 5, 'neigh_op_bnr_0')
// (21, 3, 'neigh_op_top_0')
// (21, 4, 'lutff_0/out')
// (21, 5, 'neigh_op_bot_0')
// (22, 3, 'neigh_op_tnl_0')
// (22, 4, 'local_g1_0')
// (22, 4, 'lutff_5/in_0')
// (22, 4, 'neigh_op_lft_0')
// (22, 5, 'neigh_op_bnl_0')

reg n2769 = 0;
// (20, 3, 'neigh_op_tnr_1')
// (20, 4, 'neigh_op_rgt_1')
// (20, 5, 'neigh_op_bnr_1')
// (21, 3, 'neigh_op_top_1')
// (21, 4, 'lutff_1/out')
// (21, 5, 'neigh_op_bot_1')
// (22, 3, 'neigh_op_tnl_1')
// (22, 4, 'local_g0_1')
// (22, 4, 'lutff_1/in_0')
// (22, 4, 'lutff_7/in_2')
// (22, 4, 'neigh_op_lft_1')
// (22, 5, 'neigh_op_bnl_1')

reg n2770 = 0;
// (20, 3, 'neigh_op_tnr_2')
// (20, 4, 'neigh_op_rgt_2')
// (20, 5, 'neigh_op_bnr_2')
// (21, 3, 'neigh_op_top_2')
// (21, 4, 'lutff_2/out')
// (21, 5, 'neigh_op_bot_2')
// (22, 3, 'neigh_op_tnl_2')
// (22, 4, 'local_g0_2')
// (22, 4, 'lutff_1/in_1')
// (22, 4, 'lutff_6/in_0')
// (22, 4, 'neigh_op_lft_2')
// (22, 5, 'neigh_op_bnl_2')

reg n2771 = 0;
// (20, 3, 'neigh_op_tnr_3')
// (20, 4, 'neigh_op_rgt_3')
// (20, 5, 'neigh_op_bnr_3')
// (21, 3, 'neigh_op_top_3')
// (21, 4, 'lutff_3/out')
// (21, 5, 'neigh_op_bot_3')
// (22, 3, 'neigh_op_tnl_3')
// (22, 4, 'local_g1_3')
// (22, 4, 'lutff_1/in_3')
// (22, 4, 'lutff_4/in_2')
// (22, 4, 'neigh_op_lft_3')
// (22, 5, 'neigh_op_bnl_3')

reg n2772 = 0;
// (20, 3, 'neigh_op_tnr_4')
// (20, 4, 'local_g2_4')
// (20, 4, 'lutff_1/in_3')
// (20, 4, 'neigh_op_rgt_4')
// (20, 5, 'neigh_op_bnr_4')
// (21, 3, 'neigh_op_top_4')
// (21, 4, 'lutff_4/out')
// (21, 5, 'neigh_op_bot_4')
// (22, 3, 'neigh_op_tnl_4')
// (22, 4, 'local_g1_4')
// (22, 4, 'lutff_1/in_2')
// (22, 4, 'neigh_op_lft_4')
// (22, 5, 'neigh_op_bnl_4')

reg n2773 = 0;
// (20, 3, 'neigh_op_tnr_5')
// (20, 4, 'neigh_op_rgt_5')
// (20, 5, 'neigh_op_bnr_5')
// (21, 3, 'neigh_op_top_5')
// (21, 4, 'local_g2_5')
// (21, 4, 'lutff_5/in_2')
// (21, 4, 'lutff_5/out')
// (21, 5, 'neigh_op_bot_5')
// (22, 3, 'neigh_op_tnl_5')
// (22, 4, 'local_g1_5')
// (22, 4, 'lutff_5/in_1')
// (22, 4, 'neigh_op_lft_5')
// (22, 5, 'neigh_op_bnl_5')

reg n2774 = 0;
// (20, 3, 'neigh_op_tnr_6')
// (20, 4, 'neigh_op_rgt_6')
// (20, 5, 'neigh_op_bnr_6')
// (21, 3, 'neigh_op_top_6')
// (21, 4, 'local_g0_6')
// (21, 4, 'lutff_6/in_2')
// (21, 4, 'lutff_6/out')
// (21, 5, 'neigh_op_bot_6')
// (22, 3, 'neigh_op_tnl_6')
// (22, 4, 'local_g0_6')
// (22, 4, 'lutff_5/in_3')
// (22, 4, 'neigh_op_lft_6')
// (22, 5, 'neigh_op_bnl_6')

reg n2775 = 0;
// (20, 3, 'neigh_op_tnr_7')
// (20, 4, 'local_g3_7')
// (20, 4, 'lutff_3/in_1')
// (20, 4, 'neigh_op_rgt_7')
// (20, 5, 'neigh_op_bnr_7')
// (21, 3, 'neigh_op_top_7')
// (21, 4, 'lutff_7/out')
// (21, 5, 'neigh_op_bot_7')
// (22, 3, 'neigh_op_tnl_7')
// (22, 4, 'neigh_op_lft_7')
// (22, 5, 'local_g2_7')
// (22, 5, 'lutff_3/in_2')
// (22, 5, 'neigh_op_bnl_7')

reg n2776 = 0;
// (20, 4, 'neigh_op_tnr_0')
// (20, 5, 'neigh_op_rgt_0')
// (20, 6, 'neigh_op_bnr_0')
// (21, 4, 'neigh_op_top_0')
// (21, 5, 'local_g1_0')
// (21, 5, 'lutff_0/in_1')
// (21, 5, 'lutff_0/out')
// (21, 5, 'lutff_7/in_2')
// (21, 6, 'neigh_op_bot_0')
// (22, 4, 'neigh_op_tnl_0')
// (22, 5, 'neigh_op_lft_0')
// (22, 6, 'neigh_op_bnl_0')

reg n2777 = 0;
// (20, 4, 'neigh_op_tnr_1')
// (20, 5, 'neigh_op_rgt_1')
// (20, 6, 'neigh_op_bnr_1')
// (21, 4, 'neigh_op_top_1')
// (21, 5, 'local_g3_1')
// (21, 5, 'lutff_1/in_1')
// (21, 5, 'lutff_1/out')
// (21, 5, 'lutff_7/in_1')
// (21, 6, 'neigh_op_bot_1')
// (22, 4, 'neigh_op_tnl_1')
// (22, 5, 'neigh_op_lft_1')
// (22, 6, 'neigh_op_bnl_1')

reg n2778 = 0;
// (20, 4, 'neigh_op_tnr_2')
// (20, 5, 'neigh_op_rgt_2')
// (20, 6, 'neigh_op_bnr_2')
// (21, 4, 'neigh_op_top_2')
// (21, 5, 'lutff_2/out')
// (21, 6, 'neigh_op_bot_2')
// (22, 4, 'neigh_op_tnl_2')
// (22, 5, 'local_g1_2')
// (22, 5, 'lutff_1/in_2')
// (22, 5, 'lutff_3/in_0')
// (22, 5, 'neigh_op_lft_2')
// (22, 6, 'neigh_op_bnl_2')

reg n2779 = 0;
// (20, 4, 'neigh_op_tnr_3')
// (20, 5, 'neigh_op_rgt_3')
// (20, 6, 'neigh_op_bnr_3')
// (21, 2, 'sp4_r_v_b_42')
// (21, 3, 'sp4_r_v_b_31')
// (21, 4, 'neigh_op_top_3')
// (21, 4, 'sp4_r_v_b_18')
// (21, 5, 'local_g3_3')
// (21, 5, 'lutff_3/in_1')
// (21, 5, 'lutff_3/out')
// (21, 5, 'sp4_r_v_b_7')
// (21, 6, 'neigh_op_bot_3')
// (22, 1, 'sp4_v_t_42')
// (22, 2, 'sp4_v_b_42')
// (22, 3, 'local_g3_7')
// (22, 3, 'lutff_7/in_3')
// (22, 3, 'sp4_v_b_31')
// (22, 4, 'neigh_op_tnl_3')
// (22, 4, 'sp4_v_b_18')
// (22, 5, 'neigh_op_lft_3')
// (22, 5, 'sp4_v_b_7')
// (22, 6, 'neigh_op_bnl_3')

reg n2780 = 0;
// (20, 4, 'neigh_op_tnr_4')
// (20, 5, 'neigh_op_rgt_4')
// (20, 6, 'neigh_op_bnr_4')
// (21, 4, 'neigh_op_top_4')
// (21, 5, 'local_g0_4')
// (21, 5, 'lutff_4/in_2')
// (21, 5, 'lutff_4/out')
// (21, 5, 'lutff_7/in_3')
// (21, 6, 'neigh_op_bot_4')
// (22, 4, 'neigh_op_tnl_4')
// (22, 5, 'neigh_op_lft_4')
// (22, 6, 'neigh_op_bnl_4')

reg n2781 = 0;
// (20, 4, 'neigh_op_tnr_5')
// (20, 5, 'neigh_op_rgt_5')
// (20, 6, 'neigh_op_bnr_5')
// (21, 4, 'neigh_op_top_5')
// (21, 5, 'lutff_5/out')
// (21, 6, 'neigh_op_bot_5')
// (22, 4, 'neigh_op_tnl_5')
// (22, 5, 'local_g1_5')
// (22, 5, 'lutff_3/in_3')
// (22, 5, 'lutff_4/in_0')
// (22, 5, 'neigh_op_lft_5')
// (22, 6, 'neigh_op_bnl_5')

reg n2782 = 0;
// (20, 4, 'neigh_op_tnr_6')
// (20, 5, 'neigh_op_rgt_6')
// (20, 6, 'neigh_op_bnr_6')
// (21, 4, 'neigh_op_top_6')
// (21, 5, 'local_g3_6')
// (21, 5, 'lutff_6/in_1')
// (21, 5, 'lutff_6/out')
// (21, 5, 'lutff_7/in_0')
// (21, 6, 'neigh_op_bot_6')
// (22, 4, 'neigh_op_tnl_6')
// (22, 5, 'neigh_op_lft_6')
// (22, 6, 'neigh_op_bnl_6')

wire n2783;
// (20, 4, 'neigh_op_tnr_7')
// (20, 5, 'neigh_op_rgt_7')
// (20, 6, 'neigh_op_bnr_7')
// (21, 4, 'neigh_op_top_7')
// (21, 5, 'lutff_7/out')
// (21, 6, 'neigh_op_bot_7')
// (22, 4, 'local_g3_7')
// (22, 4, 'lutff_2/in_0')
// (22, 4, 'neigh_op_tnl_7')
// (22, 5, 'neigh_op_lft_7')
// (22, 6, 'neigh_op_bnl_7')

wire n2784;
// (20, 5, 'lutff_1/cout')
// (20, 5, 'lutff_2/in_3')

wire n2785;
// (20, 6, 'lutff_1/cout')
// (20, 6, 'lutff_2/in_3')

wire n2786;
// (20, 6, 'lutff_2/cout')
// (20, 6, 'lutff_3/in_3')

wire n2787;
// (20, 6, 'lutff_3/cout')
// (20, 6, 'lutff_4/in_3')

wire n2788;
// (20, 6, 'lutff_4/cout')
// (20, 6, 'lutff_5/in_3')

wire n2789;
// (20, 6, 'lutff_5/cout')
// (20, 6, 'lutff_6/in_3')

reg n2790 = 0;
// (20, 6, 'neigh_op_tnr_1')
// (20, 7, 'local_g2_1')
// (20, 7, 'lutff_1/in_2')
// (20, 7, 'neigh_op_rgt_1')
// (20, 8, 'neigh_op_bnr_1')
// (21, 6, 'neigh_op_top_1')
// (21, 7, 'local_g1_1')
// (21, 7, 'lutff_1/in_1')
// (21, 7, 'lutff_1/out')
// (21, 8, 'neigh_op_bot_1')
// (22, 6, 'neigh_op_tnl_1')
// (22, 7, 'local_g1_1')
// (22, 7, 'lutff_4/in_0')
// (22, 7, 'neigh_op_lft_1')
// (22, 8, 'neigh_op_bnl_1')

wire n2791;
// (20, 6, 'neigh_op_tnr_2')
// (20, 7, 'neigh_op_rgt_2')
// (20, 8, 'neigh_op_bnr_2')
// (21, 6, 'neigh_op_top_2')
// (21, 7, 'lutff_2/out')
// (21, 8, 'neigh_op_bot_2')
// (22, 6, 'neigh_op_tnl_2')
// (22, 7, 'local_g1_2')
// (22, 7, 'lutff_2/in_1')
// (22, 7, 'neigh_op_lft_2')
// (22, 8, 'neigh_op_bnl_2')

wire n2792;
// (20, 6, 'neigh_op_tnr_4')
// (20, 7, 'neigh_op_rgt_4')
// (20, 8, 'neigh_op_bnr_4')
// (21, 6, 'neigh_op_top_4')
// (21, 7, 'lutff_4/out')
// (21, 7, 'sp4_h_r_8')
// (21, 8, 'neigh_op_bot_4')
// (22, 6, 'neigh_op_tnl_4')
// (22, 7, 'local_g0_5')
// (22, 7, 'lutff_6/in_3')
// (22, 7, 'neigh_op_lft_4')
// (22, 7, 'sp4_h_r_21')
// (22, 8, 'neigh_op_bnl_4')
// (23, 7, 'sp4_h_r_32')
// (24, 7, 'sp4_h_r_45')
// (25, 7, 'sp4_h_l_45')

wire n2793;
// (20, 6, 'neigh_op_tnr_6')
// (20, 7, 'neigh_op_rgt_6')
// (20, 8, 'neigh_op_bnr_6')
// (21, 6, 'neigh_op_top_6')
// (21, 7, 'lutff_6/out')
// (21, 8, 'neigh_op_bot_6')
// (22, 6, 'neigh_op_tnl_6')
// (22, 7, 'local_g0_6')
// (22, 7, 'lutff_3/in_1')
// (22, 7, 'neigh_op_lft_6')
// (22, 8, 'neigh_op_bnl_6')

reg n2794 = 0;
// (20, 7, 'local_g0_0')
// (20, 7, 'lutff_0/in_2')
// (20, 7, 'sp4_h_r_8')
// (21, 6, 'neigh_op_tnr_0')
// (21, 7, 'local_g2_0')
// (21, 7, 'local_g3_0')
// (21, 7, 'lutff_0/in_1')
// (21, 7, 'lutff_1/in_3')
// (21, 7, 'neigh_op_rgt_0')
// (21, 7, 'sp4_h_r_21')
// (21, 8, 'neigh_op_bnr_0')
// (22, 6, 'neigh_op_top_0')
// (22, 7, 'local_g0_0')
// (22, 7, 'lutff_0/in_0')
// (22, 7, 'lutff_0/out')
// (22, 7, 'lutff_4/in_2')
// (22, 7, 'sp4_h_r_32')
// (22, 8, 'neigh_op_bot_0')
// (23, 6, 'neigh_op_tnl_0')
// (23, 7, 'neigh_op_lft_0')
// (23, 7, 'sp4_h_r_45')
// (23, 8, 'neigh_op_bnl_0')
// (24, 7, 'sp4_h_l_45')

wire n2795;
// (20, 7, 'lutff_1/cout')
// (20, 7, 'lutff_2/in_3')

wire n2796;
// (20, 7, 'lutff_3/cout')
// (20, 7, 'lutff_4/in_3')

wire n2797;
// (20, 7, 'lutff_5/cout')
// (20, 7, 'lutff_6/in_3')

wire n2798;
// (20, 7, 'lutff_7/cout')
// (20, 8, 'carry_in')
// (20, 8, 'carry_in_mux')
// (20, 8, 'lutff_0/in_3')

wire n2799;
// (20, 7, 'neigh_op_tnr_0')
// (20, 8, 'neigh_op_rgt_0')
// (20, 9, 'neigh_op_bnr_0')
// (21, 7, 'neigh_op_top_0')
// (21, 8, 'local_g2_0')
// (21, 8, 'lutff_0/out')
// (21, 8, 'lutff_7/in_1')
// (21, 9, 'neigh_op_bot_0')
// (22, 7, 'neigh_op_tnl_0')
// (22, 8, 'neigh_op_lft_0')
// (22, 9, 'neigh_op_bnl_0')

wire n2800;
// (20, 7, 'neigh_op_tnr_2')
// (20, 8, 'neigh_op_rgt_2')
// (20, 9, 'neigh_op_bnr_2')
// (21, 7, 'neigh_op_top_2')
// (21, 8, 'local_g2_2')
// (21, 8, 'lutff_2/out')
// (21, 8, 'lutff_6/in_0')
// (21, 9, 'neigh_op_bot_2')
// (22, 7, 'neigh_op_tnl_2')
// (22, 8, 'neigh_op_lft_2')
// (22, 9, 'neigh_op_bnl_2')

reg n2801 = 0;
// (20, 7, 'neigh_op_tnr_4')
// (20, 8, 'neigh_op_rgt_4')
// (20, 9, 'neigh_op_bnr_4')
// (21, 7, 'neigh_op_top_4')
// (21, 8, 'local_g1_4')
// (21, 8, 'lutff_4/in_1')
// (21, 8, 'lutff_4/out')
// (21, 9, 'neigh_op_bot_4')
// (22, 7, 'neigh_op_tnl_4')
// (22, 8, 'local_g1_4')
// (22, 8, 'lutff_5/in_2')
// (22, 8, 'lutff_7/in_0')
// (22, 8, 'neigh_op_lft_4')
// (22, 9, 'neigh_op_bnl_4')

wire n2802;
// (20, 7, 'neigh_op_tnr_5')
// (20, 8, 'neigh_op_rgt_5')
// (20, 9, 'neigh_op_bnr_5')
// (21, 7, 'neigh_op_top_5')
// (21, 8, 'lutff_5/out')
// (21, 9, 'neigh_op_bot_5')
// (22, 7, 'neigh_op_tnl_5')
// (22, 8, 'local_g1_5')
// (22, 8, 'lutff_global/s_r')
// (22, 8, 'neigh_op_lft_5')
// (22, 9, 'neigh_op_bnl_5')

reg n2803 = 0;
// (20, 7, 'neigh_op_tnr_6')
// (20, 8, 'local_g3_6')
// (20, 8, 'lutff_3/in_2')
// (20, 8, 'neigh_op_rgt_6')
// (20, 9, 'neigh_op_bnr_6')
// (21, 7, 'neigh_op_top_6')
// (21, 8, 'local_g1_6')
// (21, 8, 'local_g2_6')
// (21, 8, 'lutff_3/in_1')
// (21, 8, 'lutff_6/in_3')
// (21, 8, 'lutff_6/out')
// (21, 9, 'neigh_op_bot_6')
// (22, 7, 'neigh_op_tnl_6')
// (22, 8, 'local_g0_6')
// (22, 8, 'lutff_5/in_1')
// (22, 8, 'lutff_7/in_1')
// (22, 8, 'neigh_op_lft_6')
// (22, 9, 'neigh_op_bnl_6')

reg n2804 = 0;
// (20, 7, 'neigh_op_tnr_7')
// (20, 8, 'local_g3_7')
// (20, 8, 'lutff_1/in_1')
// (20, 8, 'neigh_op_rgt_7')
// (20, 9, 'neigh_op_bnr_7')
// (21, 7, 'neigh_op_top_7')
// (21, 8, 'local_g2_7')
// (21, 8, 'lutff_1/in_2')
// (21, 8, 'lutff_7/in_2')
// (21, 8, 'lutff_7/out')
// (21, 9, 'neigh_op_bot_7')
// (22, 7, 'local_g3_7')
// (22, 7, 'lutff_7/in_3')
// (22, 7, 'neigh_op_tnl_7')
// (22, 8, 'neigh_op_lft_7')
// (22, 9, 'neigh_op_bnl_7')

wire n2805;
// (20, 8, 'lutff_1/cout')
// (20, 8, 'lutff_2/in_3')

wire n2806;
// (20, 8, 'lutff_3/cout')
// (20, 8, 'lutff_4/in_3')

reg n2807 = 0;
// (20, 9, 'neigh_op_tnr_2')
// (20, 10, 'neigh_op_rgt_2')
// (20, 11, 'neigh_op_bnr_2')
// (21, 9, 'neigh_op_top_2')
// (21, 10, 'lutff_2/out')
// (21, 10, 'sp4_r_v_b_37')
// (21, 11, 'neigh_op_bot_2')
// (21, 11, 'sp4_r_v_b_24')
// (21, 12, 'local_g2_5')
// (21, 12, 'lutff_5/in_2')
// (21, 12, 'sp4_r_v_b_13')
// (21, 13, 'sp4_r_v_b_0')
// (22, 9, 'neigh_op_tnl_2')
// (22, 9, 'sp4_v_t_37')
// (22, 10, 'neigh_op_lft_2')
// (22, 10, 'sp4_v_b_37')
// (22, 11, 'neigh_op_bnl_2')
// (22, 11, 'sp4_v_b_24')
// (22, 12, 'sp4_v_b_13')
// (22, 13, 'sp4_v_b_0')

reg n2808 = 0;
// (20, 9, 'neigh_op_tnr_5')
// (20, 10, 'neigh_op_rgt_5')
// (20, 11, 'neigh_op_bnr_5')
// (21, 9, 'neigh_op_top_5')
// (21, 10, 'lutff_5/out')
// (21, 10, 'sp4_r_v_b_43')
// (21, 11, 'neigh_op_bot_5')
// (21, 11, 'sp4_r_v_b_30')
// (21, 12, 'sp4_r_v_b_19')
// (21, 13, 'sp4_r_v_b_6')
// (22, 9, 'neigh_op_tnl_5')
// (22, 9, 'sp4_v_t_43')
// (22, 10, 'neigh_op_lft_5')
// (22, 10, 'sp4_v_b_43')
// (22, 11, 'neigh_op_bnl_5')
// (22, 11, 'sp4_v_b_30')
// (22, 12, 'sp4_v_b_19')
// (22, 13, 'local_g0_6')
// (22, 13, 'lutff_2/in_2')
// (22, 13, 'sp4_v_b_6')

reg n2809 = 0;
// (20, 9, 'sp4_r_v_b_47')
// (20, 10, 'sp4_r_v_b_34')
// (20, 11, 'sp4_r_v_b_23')
// (20, 12, 'local_g2_2')
// (20, 12, 'lutff_1/in_1')
// (20, 12, 'lutff_6/in_0')
// (20, 12, 'sp4_r_v_b_10')
// (21, 8, 'sp4_v_t_47')
// (21, 9, 'sp4_v_b_47')
// (21, 10, 'sp4_v_b_34')
// (21, 11, 'sp4_v_b_23')
// (21, 12, 'local_g0_2')
// (21, 12, 'lutff_0/in_0')
// (21, 12, 'lutff_1/in_3')
// (21, 12, 'lutff_2/in_0')
// (21, 12, 'lutff_6/in_2')
// (21, 12, 'lutff_7/in_3')
// (21, 12, 'sp4_h_r_10')
// (21, 12, 'sp4_v_b_10')
// (22, 11, 'neigh_op_tnr_1')
// (22, 12, 'local_g2_1')
// (22, 12, 'lutff_4/in_3')
// (22, 12, 'lutff_7/in_2')
// (22, 12, 'neigh_op_rgt_1')
// (22, 12, 'sp4_h_r_23')
// (22, 13, 'neigh_op_bnr_1')
// (23, 11, 'neigh_op_top_1')
// (23, 12, 'local_g2_1')
// (23, 12, 'lutff_1/in_2')
// (23, 12, 'lutff_1/out')
// (23, 12, 'sp4_h_r_34')
// (23, 13, 'neigh_op_bot_1')
// (24, 11, 'neigh_op_tnl_1')
// (24, 12, 'neigh_op_lft_1')
// (24, 12, 'sp4_h_r_47')
// (24, 13, 'neigh_op_bnl_1')
// (25, 12, 'sp4_h_l_47')

reg n2810 = 0;
// (20, 10, 'sp4_r_v_b_38')
// (20, 11, 'neigh_op_tnr_7')
// (20, 11, 'sp4_r_v_b_27')
// (20, 12, 'neigh_op_rgt_7')
// (20, 12, 'sp4_r_v_b_14')
// (20, 13, 'neigh_op_bnr_7')
// (20, 13, 'sp4_r_v_b_3')
// (21, 9, 'sp4_v_t_38')
// (21, 10, 'sp4_v_b_38')
// (21, 11, 'neigh_op_top_7')
// (21, 11, 'sp4_v_b_27')
// (21, 12, 'lutff_7/out')
// (21, 12, 'sp4_v_b_14')
// (21, 13, 'neigh_op_bot_7')
// (21, 13, 'sp4_h_r_9')
// (21, 13, 'sp4_v_b_3')
// (22, 11, 'neigh_op_tnl_7')
// (22, 12, 'neigh_op_lft_7')
// (22, 13, 'neigh_op_bnl_7')
// (22, 13, 'sp4_h_r_20')
// (23, 13, 'local_g2_1')
// (23, 13, 'lutff_6/in_3')
// (23, 13, 'sp4_h_r_33')
// (24, 13, 'sp4_h_r_44')
// (25, 13, 'sp4_h_l_44')

reg n2811 = 0;
// (20, 11, 'neigh_op_tnr_0')
// (20, 12, 'neigh_op_rgt_0')
// (20, 13, 'neigh_op_bnr_0')
// (21, 10, 'sp4_r_v_b_41')
// (21, 11, 'neigh_op_top_0')
// (21, 11, 'sp4_r_v_b_28')
// (21, 12, 'lutff_0/out')
// (21, 12, 'sp4_r_v_b_17')
// (21, 13, 'neigh_op_bot_0')
// (21, 13, 'sp4_r_v_b_4')
// (22, 9, 'sp4_v_t_41')
// (22, 10, 'sp4_v_b_41')
// (22, 11, 'neigh_op_tnl_0')
// (22, 11, 'sp4_v_b_28')
// (22, 12, 'neigh_op_lft_0')
// (22, 12, 'sp4_v_b_17')
// (22, 13, 'neigh_op_bnl_0')
// (22, 13, 'sp4_h_r_4')
// (22, 13, 'sp4_v_b_4')
// (23, 13, 'local_g0_1')
// (23, 13, 'lutff_2/in_1')
// (23, 13, 'sp4_h_r_17')
// (24, 13, 'sp4_h_r_28')
// (25, 13, 'sp4_h_r_41')

reg n2812 = 0;
// (20, 11, 'neigh_op_tnr_1')
// (20, 12, 'neigh_op_rgt_1')
// (20, 13, 'neigh_op_bnr_1')
// (21, 11, 'neigh_op_top_1')
// (21, 11, 'sp4_r_v_b_46')
// (21, 12, 'lutff_1/out')
// (21, 12, 'sp4_r_v_b_35')
// (21, 13, 'neigh_op_bot_1')
// (21, 13, 'sp4_r_v_b_22')
// (21, 14, 'local_g2_3')
// (21, 14, 'lutff_3/in_0')
// (21, 14, 'sp4_r_v_b_11')
// (22, 10, 'sp4_v_t_46')
// (22, 11, 'neigh_op_tnl_1')
// (22, 11, 'sp4_v_b_46')
// (22, 12, 'neigh_op_lft_1')
// (22, 12, 'sp4_v_b_35')
// (22, 13, 'neigh_op_bnl_1')
// (22, 13, 'sp4_v_b_22')
// (22, 14, 'sp4_v_b_11')

reg n2813 = 0;
// (20, 11, 'neigh_op_tnr_2')
// (20, 12, 'neigh_op_rgt_2')
// (20, 12, 'sp4_r_v_b_36')
// (20, 13, 'neigh_op_bnr_2')
// (20, 13, 'sp4_r_v_b_25')
// (20, 14, 'sp4_r_v_b_12')
// (20, 15, 'sp4_r_v_b_1')
// (21, 11, 'neigh_op_top_2')
// (21, 11, 'sp4_v_t_36')
// (21, 12, 'lutff_2/out')
// (21, 12, 'sp4_v_b_36')
// (21, 13, 'neigh_op_bot_2')
// (21, 13, 'sp4_v_b_25')
// (21, 14, 'local_g0_4')
// (21, 14, 'lutff_0/in_2')
// (21, 14, 'sp4_v_b_12')
// (21, 15, 'sp4_v_b_1')
// (22, 11, 'neigh_op_tnl_2')
// (22, 12, 'neigh_op_lft_2')
// (22, 13, 'neigh_op_bnl_2')

wire n2814;
// (20, 11, 'neigh_op_tnr_3')
// (20, 12, 'neigh_op_rgt_3')
// (20, 13, 'local_g0_3')
// (20, 13, 'lutff_0/in_3')
// (20, 13, 'lutff_4/in_1')
// (20, 13, 'lutff_5/in_2')
// (20, 13, 'neigh_op_bnr_3')
// (21, 11, 'neigh_op_top_3')
// (21, 12, 'local_g1_3')
// (21, 12, 'lutff_3/out')
// (21, 12, 'lutff_5/in_1')
// (21, 13, 'neigh_op_bot_3')
// (22, 11, 'neigh_op_tnl_3')
// (22, 12, 'local_g0_3')
// (22, 12, 'lutff_2/in_1')
// (22, 12, 'neigh_op_lft_3')
// (22, 13, 'local_g3_3')
// (22, 13, 'lutff_0/in_2')
// (22, 13, 'lutff_2/in_0')
// (22, 13, 'lutff_3/in_3')
// (22, 13, 'neigh_op_bnl_3')

reg n2815 = 0;
// (20, 11, 'neigh_op_tnr_4')
// (20, 12, 'neigh_op_rgt_4')
// (20, 13, 'neigh_op_bnr_4')
// (21, 11, 'neigh_op_top_4')
// (21, 11, 'sp4_r_v_b_36')
// (21, 12, 'lutff_4/out')
// (21, 12, 'sp4_r_v_b_25')
// (21, 13, 'neigh_op_bot_4')
// (21, 13, 'sp4_r_v_b_12')
// (21, 14, 'local_g1_1')
// (21, 14, 'lutff_7/in_1')
// (21, 14, 'sp4_r_v_b_1')
// (22, 10, 'sp4_v_t_36')
// (22, 11, 'neigh_op_tnl_4')
// (22, 11, 'sp4_v_b_36')
// (22, 12, 'neigh_op_lft_4')
// (22, 12, 'sp4_v_b_25')
// (22, 13, 'neigh_op_bnl_4')
// (22, 13, 'sp4_v_b_12')
// (22, 14, 'sp4_v_b_1')

reg n2816 = 0;
// (20, 11, 'neigh_op_tnr_5')
// (20, 12, 'neigh_op_rgt_5')
// (20, 12, 'sp4_r_v_b_42')
// (20, 13, 'neigh_op_bnr_5')
// (20, 13, 'sp4_r_v_b_31')
// (20, 14, 'sp4_r_v_b_18')
// (20, 15, 'sp4_r_v_b_7')
// (21, 11, 'neigh_op_top_5')
// (21, 11, 'sp4_v_t_42')
// (21, 12, 'lutff_5/out')
// (21, 12, 'sp4_v_b_42')
// (21, 13, 'neigh_op_bot_5')
// (21, 13, 'sp4_v_b_31')
// (21, 14, 'local_g0_2')
// (21, 14, 'lutff_2/in_0')
// (21, 14, 'sp4_v_b_18')
// (21, 15, 'sp4_v_b_7')
// (22, 11, 'neigh_op_tnl_5')
// (22, 12, 'neigh_op_lft_5')
// (22, 13, 'neigh_op_bnl_5')

wire n2817;
// (20, 11, 'neigh_op_tnr_6')
// (20, 12, 'neigh_op_rgt_6')
// (20, 13, 'local_g0_6')
// (20, 13, 'lutff_1/in_1')
// (20, 13, 'lutff_2/in_0')
// (20, 13, 'lutff_6/in_2')
// (20, 13, 'lutff_7/in_1')
// (20, 13, 'neigh_op_bnr_6')
// (21, 11, 'neigh_op_top_6')
// (21, 12, 'local_g0_6')
// (21, 12, 'lutff_3/in_1')
// (21, 12, 'lutff_6/out')
// (21, 13, 'neigh_op_bot_6')
// (22, 11, 'neigh_op_tnl_6')
// (22, 12, 'neigh_op_lft_6')
// (22, 13, 'neigh_op_bnl_6')

reg n2818 = 0;
// (20, 11, 'sp4_r_v_b_37')
// (20, 12, 'sp4_r_v_b_24')
// (20, 13, 'sp4_r_v_b_13')
// (20, 14, 'local_g1_1')
// (20, 14, 'lutff_7/in_3')
// (20, 14, 'sp4_h_r_1')
// (20, 14, 'sp4_r_v_b_0')
// (20, 15, 'local_g2_4')
// (20, 15, 'lutff_7/in_3')
// (20, 15, 'sp4_r_v_b_36')
// (20, 16, 'sp4_r_v_b_25')
// (20, 17, 'sp4_r_v_b_12')
// (20, 18, 'sp4_r_v_b_1')
// (21, 10, 'sp4_v_t_37')
// (21, 11, 'sp4_r_v_b_42')
// (21, 11, 'sp4_v_b_37')
// (21, 12, 'sp4_r_v_b_31')
// (21, 12, 'sp4_v_b_24')
// (21, 13, 'local_g0_5')
// (21, 13, 'lutff_0/in_1')
// (21, 13, 'lutff_6/in_1')
// (21, 13, 'sp4_r_v_b_18')
// (21, 13, 'sp4_v_b_13')
// (21, 14, 'local_g1_4')
// (21, 14, 'lutff_1/in_0')
// (21, 14, 'sp4_h_r_12')
// (21, 14, 'sp4_h_r_7')
// (21, 14, 'sp4_r_v_b_7')
// (21, 14, 'sp4_v_b_0')
// (21, 14, 'sp4_v_t_36')
// (21, 15, 'local_g2_7')
// (21, 15, 'lutff_0/in_3')
// (21, 15, 'lutff_5/in_0')
// (21, 15, 'sp4_r_v_b_39')
// (21, 15, 'sp4_v_b_36')
// (21, 16, 'sp4_r_v_b_26')
// (21, 16, 'sp4_v_b_25')
// (21, 17, 'sp4_r_v_b_15')
// (21, 17, 'sp4_v_b_12')
// (21, 18, 'sp4_r_v_b_2')
// (21, 18, 'sp4_v_b_1')
// (22, 10, 'sp4_v_t_42')
// (22, 11, 'sp4_v_b_42')
// (22, 12, 'sp4_v_b_31')
// (22, 13, 'local_g1_2')
// (22, 13, 'lutff_7/in_0')
// (22, 13, 'sp4_v_b_18')
// (22, 14, 'sp4_h_r_18')
// (22, 14, 'sp4_h_r_2')
// (22, 14, 'sp4_h_r_25')
// (22, 14, 'sp4_v_b_7')
// (22, 14, 'sp4_v_t_39')
// (22, 15, 'sp4_v_b_39')
// (22, 16, 'sp4_v_b_26')
// (22, 17, 'sp4_v_b_15')
// (22, 18, 'sp4_v_b_2')
// (23, 13, 'neigh_op_tnr_5')
// (23, 14, 'neigh_op_rgt_5')
// (23, 14, 'sp4_h_r_15')
// (23, 14, 'sp4_h_r_31')
// (23, 14, 'sp4_h_r_36')
// (23, 15, 'neigh_op_bnr_5')
// (24, 13, 'neigh_op_top_5')
// (24, 14, 'local_g1_5')
// (24, 14, 'lutff_5/in_3')
// (24, 14, 'lutff_5/out')
// (24, 14, 'sp4_h_l_36')
// (24, 14, 'sp4_h_r_10')
// (24, 14, 'sp4_h_r_26')
// (24, 14, 'sp4_h_r_42')
// (24, 15, 'neigh_op_bot_5')
// (25, 13, 'neigh_op_tnl_5')
// (25, 14, 'neigh_op_lft_5')
// (25, 14, 'sp4_h_l_42')
// (25, 14, 'sp4_h_r_23')
// (25, 14, 'sp4_h_r_39')
// (25, 15, 'neigh_op_bnl_5')

wire n2819;
// (20, 11, 'sp4_r_v_b_43')
// (20, 12, 'sp4_r_v_b_30')
// (20, 13, 'sp4_r_v_b_19')
// (20, 14, 'sp4_r_v_b_6')
// (21, 10, 'sp4_v_t_43')
// (21, 11, 'sp4_v_b_43')
// (21, 12, 'sp4_v_b_30')
// (21, 13, 'local_g1_3')
// (21, 13, 'lutff_global/cen')
// (21, 13, 'sp4_v_b_19')
// (21, 14, 'sp4_h_r_6')
// (21, 14, 'sp4_v_b_6')
// (22, 13, 'neigh_op_tnr_7')
// (22, 14, 'neigh_op_rgt_7')
// (22, 14, 'sp4_h_r_19')
// (22, 14, 'sp4_h_r_3')
// (22, 15, 'neigh_op_bnr_7')
// (23, 13, 'neigh_op_top_7')
// (23, 14, 'local_g2_7')
// (23, 14, 'lutff_1/in_2')
// (23, 14, 'lutff_7/out')
// (23, 14, 'sp4_h_r_14')
// (23, 14, 'sp4_h_r_30')
// (23, 15, 'neigh_op_bot_7')
// (24, 13, 'neigh_op_tnl_7')
// (24, 14, 'local_g3_3')
// (24, 14, 'lutff_global/cen')
// (24, 14, 'neigh_op_lft_7')
// (24, 14, 'sp4_h_r_27')
// (24, 14, 'sp4_h_r_43')
// (24, 15, 'neigh_op_bnl_7')
// (25, 14, 'sp4_h_l_43')
// (25, 14, 'sp4_h_r_38')

reg n2820 = 0;
// (20, 12, 'neigh_op_tnr_2')
// (20, 13, 'neigh_op_rgt_2')
// (20, 13, 'sp4_r_v_b_36')
// (20, 14, 'local_g0_2')
// (20, 14, 'lutff_1/in_1')
// (20, 14, 'neigh_op_bnr_2')
// (20, 14, 'sp4_r_v_b_25')
// (20, 15, 'sp4_r_v_b_12')
// (20, 16, 'sp4_r_v_b_1')
// (21, 12, 'neigh_op_top_2')
// (21, 12, 'sp4_v_t_36')
// (21, 13, 'local_g1_2')
// (21, 13, 'lutff_2/in_1')
// (21, 13, 'lutff_2/out')
// (21, 13, 'lutff_7/in_2')
// (21, 13, 'sp4_v_b_36')
// (21, 14, 'neigh_op_bot_2')
// (21, 14, 'sp4_v_b_25')
// (21, 15, 'local_g1_4')
// (21, 15, 'lutff_0/in_1')
// (21, 15, 'lutff_4/in_3')
// (21, 15, 'sp4_v_b_12')
// (21, 16, 'sp4_v_b_1')
// (22, 12, 'neigh_op_tnl_2')
// (22, 13, 'neigh_op_lft_2')
// (22, 14, 'neigh_op_bnl_2')

reg n2821 = 0;
// (20, 12, 'neigh_op_tnr_3')
// (20, 13, 'neigh_op_rgt_3')
// (20, 13, 'sp4_r_v_b_38')
// (20, 14, 'local_g0_3')
// (20, 14, 'lutff_2/in_1')
// (20, 14, 'neigh_op_bnr_3')
// (20, 14, 'sp4_r_v_b_27')
// (20, 15, 'sp4_r_v_b_14')
// (20, 16, 'sp4_r_v_b_3')
// (21, 12, 'neigh_op_top_3')
// (21, 12, 'sp4_v_t_38')
// (21, 13, 'local_g0_3')
// (21, 13, 'lutff_3/in_0')
// (21, 13, 'lutff_3/out')
// (21, 13, 'sp4_v_b_38')
// (21, 14, 'neigh_op_bot_3')
// (21, 14, 'sp4_v_b_27')
// (21, 15, 'local_g0_6')
// (21, 15, 'lutff_0/in_0')
// (21, 15, 'lutff_4/in_0')
// (21, 15, 'sp4_v_b_14')
// (21, 16, 'sp4_v_b_3')
// (22, 12, 'neigh_op_tnl_3')
// (22, 13, 'neigh_op_lft_3')
// (22, 14, 'neigh_op_bnl_3')

wire n2822;
// (20, 12, 'neigh_op_tnr_4')
// (20, 13, 'neigh_op_rgt_4')
// (20, 14, 'local_g1_4')
// (20, 14, 'lutff_7/in_2')
// (20, 14, 'neigh_op_bnr_4')
// (21, 12, 'neigh_op_top_4')
// (21, 13, 'lutff_4/out')
// (21, 14, 'neigh_op_bot_4')
// (22, 12, 'neigh_op_tnl_4')
// (22, 13, 'neigh_op_lft_4')
// (22, 14, 'neigh_op_bnl_4')

wire n2823;
// (20, 12, 'neigh_op_tnr_5')
// (20, 13, 'neigh_op_rgt_5')
// (20, 14, 'neigh_op_bnr_5')
// (21, 12, 'neigh_op_top_5')
// (21, 13, 'local_g1_5')
// (21, 13, 'lutff_5/out')
// (21, 13, 'lutff_global/s_r')
// (21, 14, 'neigh_op_bot_5')
// (22, 12, 'neigh_op_tnl_5')
// (22, 13, 'neigh_op_lft_5')
// (22, 14, 'neigh_op_bnl_5')

reg n2824 = 0;
// (20, 12, 'neigh_op_tnr_6')
// (20, 13, 'neigh_op_rgt_6')
// (20, 13, 'sp4_r_v_b_44')
// (20, 14, 'local_g1_6')
// (20, 14, 'lutff_0/in_1')
// (20, 14, 'lutff_7/in_0')
// (20, 14, 'neigh_op_bnr_6')
// (20, 14, 'sp4_r_v_b_33')
// (20, 15, 'sp4_r_v_b_20')
// (20, 16, 'sp4_r_v_b_9')
// (21, 12, 'neigh_op_top_6')
// (21, 12, 'sp4_v_t_44')
// (21, 13, 'local_g1_6')
// (21, 13, 'lutff_1/in_2')
// (21, 13, 'lutff_6/in_3')
// (21, 13, 'lutff_6/out')
// (21, 13, 'lutff_7/in_0')
// (21, 13, 'sp4_v_b_44')
// (21, 14, 'local_g0_6')
// (21, 14, 'lutff_6/in_2')
// (21, 14, 'neigh_op_bot_6')
// (21, 14, 'sp4_v_b_33')
// (21, 15, 'local_g0_4')
// (21, 15, 'lutff_0/in_2')
// (21, 15, 'lutff_4/in_2')
// (21, 15, 'sp4_v_b_20')
// (21, 16, 'sp4_v_b_9')
// (22, 12, 'neigh_op_tnl_6')
// (22, 13, 'neigh_op_lft_6')
// (22, 14, 'neigh_op_bnl_6')

wire n2825;
// (20, 12, 'neigh_op_tnr_7')
// (20, 13, 'neigh_op_rgt_7')
// (20, 14, 'neigh_op_bnr_7')
// (21, 12, 'neigh_op_top_7')
// (21, 13, 'local_g3_7')
// (21, 13, 'lutff_4/in_2')
// (21, 13, 'lutff_7/out')
// (21, 14, 'local_g1_7')
// (21, 14, 'lutff_1/in_1')
// (21, 14, 'lutff_5/in_1')
// (21, 14, 'neigh_op_bot_7')
// (22, 12, 'neigh_op_tnl_7')
// (22, 13, 'local_g1_7')
// (22, 13, 'lutff_7/in_1')
// (22, 13, 'neigh_op_lft_7')
// (22, 14, 'neigh_op_bnl_7')

wire n2826;
// (20, 12, 'sp4_h_r_10')
// (21, 11, 'neigh_op_tnr_1')
// (21, 12, 'neigh_op_rgt_1')
// (21, 12, 'sp4_h_r_23')
// (21, 13, 'neigh_op_bnr_1')
// (22, 11, 'neigh_op_top_1')
// (22, 11, 'sp4_r_v_b_46')
// (22, 12, 'lutff_1/out')
// (22, 12, 'sp4_h_r_34')
// (22, 12, 'sp4_r_v_b_35')
// (22, 13, 'neigh_op_bot_1')
// (22, 13, 'sp4_r_v_b_22')
// (22, 14, 'sp4_r_v_b_11')
// (23, 9, 'sp4_r_v_b_43')
// (23, 10, 'sp4_r_v_b_30')
// (23, 10, 'sp4_v_t_46')
// (23, 11, 'local_g3_3')
// (23, 11, 'lutff_global/cen')
// (23, 11, 'neigh_op_tnl_1')
// (23, 11, 'sp4_r_v_b_19')
// (23, 11, 'sp4_v_b_46')
// (23, 12, 'local_g3_3')
// (23, 12, 'lutff_global/cen')
// (23, 12, 'neigh_op_lft_1')
// (23, 12, 'sp4_h_r_47')
// (23, 12, 'sp4_r_v_b_6')
// (23, 12, 'sp4_v_b_35')
// (23, 13, 'neigh_op_bnl_1')
// (23, 13, 'sp4_v_b_22')
// (23, 14, 'sp4_v_b_11')
// (24, 8, 'sp4_v_t_43')
// (24, 9, 'sp4_v_b_43')
// (24, 10, 'sp4_v_b_30')
// (24, 11, 'sp4_v_b_19')
// (24, 12, 'sp4_h_l_47')
// (24, 12, 'sp4_h_r_6')
// (24, 12, 'sp4_v_b_6')
// (25, 12, 'sp4_h_r_19')

wire n2827;
// (20, 12, 'sp4_r_v_b_37')
// (20, 13, 'sp4_r_v_b_24')
// (20, 14, 'neigh_op_tnr_0')
// (20, 14, 'sp4_r_v_b_13')
// (20, 15, 'local_g3_0')
// (20, 15, 'lutff_7/in_0')
// (20, 15, 'neigh_op_rgt_0')
// (20, 15, 'sp4_h_r_5')
// (20, 15, 'sp4_r_v_b_0')
// (20, 16, 'neigh_op_bnr_0')
// (21, 11, 'sp4_v_t_37')
// (21, 12, 'sp4_v_b_37')
// (21, 13, 'local_g2_0')
// (21, 13, 'lutff_5/in_3')
// (21, 13, 'sp4_v_b_24')
// (21, 14, 'neigh_op_top_0')
// (21, 14, 'sp4_v_b_13')
// (21, 15, 'lutff_0/out')
// (21, 15, 'sp4_h_r_0')
// (21, 15, 'sp4_h_r_16')
// (21, 15, 'sp4_v_b_0')
// (21, 16, 'neigh_op_bot_0')
// (22, 14, 'neigh_op_tnl_0')
// (22, 15, 'neigh_op_lft_0')
// (22, 15, 'sp4_h_r_13')
// (22, 15, 'sp4_h_r_29')
// (22, 16, 'neigh_op_bnl_0')
// (23, 12, 'sp4_r_v_b_40')
// (23, 13, 'sp4_r_v_b_29')
// (23, 14, 'local_g3_0')
// (23, 14, 'lutff_1/in_0')
// (23, 14, 'sp4_r_v_b_16')
// (23, 15, 'sp4_h_r_24')
// (23, 15, 'sp4_h_r_40')
// (23, 15, 'sp4_r_v_b_5')
// (24, 11, 'sp4_v_t_40')
// (24, 12, 'sp4_r_v_b_37')
// (24, 12, 'sp4_v_b_40')
// (24, 13, 'sp4_r_v_b_24')
// (24, 13, 'sp4_v_b_29')
// (24, 14, 'local_g2_5')
// (24, 14, 'lutff_5/in_2')
// (24, 14, 'sp4_r_v_b_13')
// (24, 14, 'sp4_v_b_16')
// (24, 15, 'sp4_h_l_40')
// (24, 15, 'sp4_h_r_37')
// (24, 15, 'sp4_r_v_b_0')
// (24, 15, 'sp4_v_b_5')
// (25, 11, 'sp4_v_t_37')
// (25, 12, 'sp4_v_b_37')
// (25, 13, 'sp4_v_b_24')
// (25, 14, 'sp4_v_b_13')
// (25, 15, 'sp4_h_l_37')
// (25, 15, 'sp4_v_b_0')

wire n2828;
// (20, 12, 'sp4_r_v_b_47')
// (20, 13, 'sp4_r_v_b_34')
// (20, 14, 'sp4_r_v_b_23')
// (20, 15, 'neigh_op_tnr_5')
// (20, 15, 'sp4_r_v_b_10')
// (20, 16, 'neigh_op_rgt_5')
// (20, 16, 'sp4_r_v_b_42')
// (20, 17, 'neigh_op_bnr_5')
// (20, 17, 'sp4_r_v_b_31')
// (20, 18, 'sp4_r_v_b_18')
// (20, 19, 'sp4_r_v_b_7')
// (21, 11, 'sp4_v_t_47')
// (21, 12, 'sp4_v_b_47')
// (21, 13, 'sp4_v_b_34')
// (21, 14, 'sp4_v_b_23')
// (21, 15, 'local_g0_2')
// (21, 15, 'lutff_global/cen')
// (21, 15, 'neigh_op_top_5')
// (21, 15, 'sp4_v_b_10')
// (21, 15, 'sp4_v_t_42')
// (21, 16, 'lutff_5/out')
// (21, 16, 'sp4_v_b_42')
// (21, 17, 'neigh_op_bot_5')
// (21, 17, 'sp4_v_b_31')
// (21, 18, 'sp4_v_b_18')
// (21, 19, 'sp4_v_b_7')
// (22, 15, 'neigh_op_tnl_5')
// (22, 16, 'neigh_op_lft_5')
// (22, 17, 'neigh_op_bnl_5')

reg n2829 = 0;
// (20, 13, 'neigh_op_tnr_0')
// (20, 14, 'neigh_op_rgt_0')
// (20, 15, 'neigh_op_bnr_0')
// (21, 13, 'neigh_op_top_0')
// (21, 14, 'local_g2_0')
// (21, 14, 'lutff_0/out')
// (21, 14, 'lutff_1/in_3')
// (21, 15, 'neigh_op_bot_0')
// (22, 13, 'neigh_op_tnl_0')
// (22, 14, 'neigh_op_lft_0')
// (22, 15, 'neigh_op_bnl_0')

wire n2830;
// (20, 13, 'neigh_op_tnr_1')
// (20, 14, 'neigh_op_rgt_1')
// (20, 15, 'neigh_op_bnr_1')
// (21, 13, 'neigh_op_top_1')
// (21, 14, 'local_g3_1')
// (21, 14, 'lutff_1/out')
// (21, 14, 'lutff_6/in_0')
// (21, 15, 'neigh_op_bot_1')
// (22, 13, 'neigh_op_tnl_1')
// (22, 14, 'neigh_op_lft_1')
// (22, 15, 'neigh_op_bnl_1')

reg n2831 = 0;
// (20, 13, 'neigh_op_tnr_2')
// (20, 14, 'neigh_op_rgt_2')
// (20, 15, 'neigh_op_bnr_2')
// (21, 13, 'neigh_op_top_2')
// (21, 14, 'local_g1_2')
// (21, 14, 'lutff_2/out')
// (21, 14, 'lutff_5/in_2')
// (21, 15, 'neigh_op_bot_2')
// (22, 13, 'neigh_op_tnl_2')
// (22, 14, 'neigh_op_lft_2')
// (22, 15, 'neigh_op_bnl_2')

reg n2832 = 0;
// (20, 13, 'neigh_op_tnr_3')
// (20, 14, 'neigh_op_rgt_3')
// (20, 15, 'neigh_op_bnr_3')
// (21, 13, 'neigh_op_top_3')
// (21, 14, 'local_g0_3')
// (21, 14, 'lutff_1/in_2')
// (21, 14, 'lutff_3/out')
// (21, 15, 'neigh_op_bot_3')
// (22, 13, 'neigh_op_tnl_3')
// (22, 14, 'neigh_op_lft_3')
// (22, 15, 'neigh_op_bnl_3')

reg n2833 = 0;
// (20, 13, 'neigh_op_tnr_4')
// (20, 14, 'neigh_op_rgt_4')
// (20, 15, 'neigh_op_bnr_4')
// (21, 13, 'local_g0_4')
// (21, 13, 'lutff_4/in_0')
// (21, 13, 'neigh_op_top_4')
// (21, 14, 'lutff_4/out')
// (21, 15, 'neigh_op_bot_4')
// (22, 13, 'neigh_op_tnl_4')
// (22, 14, 'neigh_op_lft_4')
// (22, 15, 'neigh_op_bnl_4')

wire n2834;
// (20, 13, 'neigh_op_tnr_5')
// (20, 14, 'local_g3_5')
// (20, 14, 'lutff_7/in_1')
// (20, 14, 'neigh_op_rgt_5')
// (20, 15, 'neigh_op_bnr_5')
// (21, 13, 'neigh_op_top_5')
// (21, 14, 'lutff_5/out')
// (21, 15, 'neigh_op_bot_5')
// (22, 13, 'neigh_op_tnl_5')
// (22, 14, 'neigh_op_lft_5')
// (22, 15, 'neigh_op_bnl_5')

wire n2835;
// (20, 13, 'neigh_op_tnr_6')
// (20, 14, 'local_g3_6')
// (20, 14, 'lutff_3/in_2')
// (20, 14, 'neigh_op_rgt_6')
// (20, 15, 'neigh_op_bnr_6')
// (21, 13, 'neigh_op_top_6')
// (21, 14, 'lutff_6/out')
// (21, 15, 'neigh_op_bot_6')
// (22, 13, 'neigh_op_tnl_6')
// (22, 14, 'neigh_op_lft_6')
// (22, 15, 'neigh_op_bnl_6')

reg n2836 = 0;
// (20, 13, 'neigh_op_tnr_7')
// (20, 14, 'neigh_op_rgt_7')
// (20, 15, 'neigh_op_bnr_7')
// (21, 13, 'neigh_op_top_7')
// (21, 14, 'local_g3_7')
// (21, 14, 'lutff_5/in_3')
// (21, 14, 'lutff_7/out')
// (21, 15, 'neigh_op_bot_7')
// (22, 13, 'neigh_op_tnl_7')
// (22, 14, 'neigh_op_lft_7')
// (22, 15, 'neigh_op_bnl_7')

wire n2837;
// (20, 14, 'lutff_1/cout')
// (20, 14, 'lutff_2/in_3')

wire n2838;
// (20, 14, 'lutff_2/cout')
// (20, 14, 'lutff_3/in_3')

reg n2839 = 0;
// (20, 14, 'neigh_op_tnr_3')
// (20, 15, 'neigh_op_rgt_3')
// (20, 16, 'neigh_op_bnr_3')
// (21, 14, 'neigh_op_top_3')
// (21, 15, 'lutff_3/out')
// (21, 16, 'local_g0_3')
// (21, 16, 'lutff_3/in_0')
// (21, 16, 'neigh_op_bot_3')
// (22, 14, 'neigh_op_tnl_3')
// (22, 15, 'neigh_op_lft_3')
// (22, 16, 'neigh_op_bnl_3')

wire n2840;
// (20, 14, 'neigh_op_tnr_4')
// (20, 15, 'local_g3_4')
// (20, 15, 'lutff_7/in_2')
// (20, 15, 'neigh_op_rgt_4')
// (20, 16, 'neigh_op_bnr_4')
// (21, 14, 'neigh_op_top_4')
// (21, 15, 'local_g3_4')
// (21, 15, 'lutff_4/out')
// (21, 15, 'lutff_5/in_2')
// (21, 16, 'neigh_op_bot_4')
// (22, 14, 'neigh_op_tnl_4')
// (22, 15, 'neigh_op_lft_4')
// (22, 16, 'neigh_op_bnl_4')

wire n2841;
// (20, 14, 'neigh_op_tnr_5')
// (20, 15, 'neigh_op_rgt_5')
// (20, 15, 'sp4_r_v_b_42')
// (20, 16, 'neigh_op_bnr_5')
// (20, 16, 'sp4_r_v_b_31')
// (20, 17, 'sp4_r_v_b_18')
// (20, 18, 'sp4_r_v_b_7')
// (21, 12, 'sp4_r_v_b_46')
// (21, 13, 'local_g0_0')
// (21, 13, 'lutff_5/in_1')
// (21, 13, 'sp4_r_v_b_35')
// (21, 14, 'neigh_op_top_5')
// (21, 14, 'sp4_h_r_0')
// (21, 14, 'sp4_r_v_b_22')
// (21, 14, 'sp4_r_v_b_38')
// (21, 14, 'sp4_v_t_42')
// (21, 15, 'lutff_5/out')
// (21, 15, 'sp4_h_r_10')
// (21, 15, 'sp4_r_v_b_11')
// (21, 15, 'sp4_r_v_b_27')
// (21, 15, 'sp4_v_b_42')
// (21, 16, 'neigh_op_bot_5')
// (21, 16, 'sp4_r_v_b_14')
// (21, 16, 'sp4_v_b_31')
// (21, 17, 'sp4_r_v_b_3')
// (21, 17, 'sp4_v_b_18')
// (21, 18, 'sp4_v_b_7')
// (22, 11, 'sp4_v_t_46')
// (22, 12, 'sp4_v_b_46')
// (22, 13, 'sp4_h_r_3')
// (22, 13, 'sp4_v_b_35')
// (22, 13, 'sp4_v_t_38')
// (22, 14, 'neigh_op_tnl_5')
// (22, 14, 'sp4_h_r_13')
// (22, 14, 'sp4_v_b_22')
// (22, 14, 'sp4_v_b_38')
// (22, 15, 'neigh_op_lft_5')
// (22, 15, 'sp4_h_r_23')
// (22, 15, 'sp4_v_b_11')
// (22, 15, 'sp4_v_b_27')
// (22, 16, 'neigh_op_bnl_5')
// (22, 16, 'sp4_v_b_14')
// (22, 17, 'sp4_v_b_3')
// (23, 13, 'local_g1_6')
// (23, 13, 'lutff_1/in_0')
// (23, 13, 'lutff_7/in_0')
// (23, 13, 'sp4_h_r_14')
// (23, 14, 'sp4_h_r_24')
// (23, 15, 'local_g3_2')
// (23, 15, 'lutff_0/in_1')
// (23, 15, 'sp4_h_r_34')
// (24, 13, 'sp4_h_r_27')
// (24, 14, 'local_g3_5')
// (24, 14, 'lutff_global/s_r')
// (24, 14, 'sp4_h_r_37')
// (24, 15, 'sp4_h_r_47')
// (25, 13, 'sp4_h_r_38')
// (25, 14, 'sp4_h_l_37')
// (25, 15, 'sp4_h_l_47')

wire n2842;
// (20, 14, 'sp4_h_r_6')
// (21, 14, 'local_g1_3')
// (21, 14, 'lutff_global/cen')
// (21, 14, 'sp4_h_r_19')
// (22, 12, 'neigh_op_tnr_1')
// (22, 13, 'neigh_op_rgt_1')
// (22, 13, 'sp4_h_r_7')
// (22, 14, 'neigh_op_bnr_1')
// (22, 14, 'sp4_h_r_30')
// (23, 11, 'sp4_r_v_b_43')
// (23, 12, 'neigh_op_top_1')
// (23, 12, 'sp4_r_v_b_30')
// (23, 13, 'local_g0_2')
// (23, 13, 'lutff_1/out')
// (23, 13, 'lutff_global/cen')
// (23, 13, 'sp4_h_r_18')
// (23, 13, 'sp4_r_v_b_19')
// (23, 14, 'neigh_op_bot_1')
// (23, 14, 'sp4_h_r_43')
// (23, 14, 'sp4_r_v_b_6')
// (24, 10, 'sp4_v_t_43')
// (24, 11, 'sp4_v_b_43')
// (24, 12, 'neigh_op_tnl_1')
// (24, 12, 'sp4_v_b_30')
// (24, 13, 'neigh_op_lft_1')
// (24, 13, 'sp4_h_r_31')
// (24, 13, 'sp4_v_b_19')
// (24, 14, 'neigh_op_bnl_1')
// (24, 14, 'sp4_h_l_43')
// (24, 14, 'sp4_v_b_6')
// (25, 13, 'sp4_h_r_42')

wire n2843;
// (20, 15, 'neigh_op_tnr_0')
// (20, 16, 'neigh_op_rgt_0')
// (20, 17, 'local_g1_0')
// (20, 17, 'lutff_0/in_1')
// (20, 17, 'neigh_op_bnr_0')
// (21, 15, 'neigh_op_top_0')
// (21, 16, 'lutff_0/out')
// (21, 17, 'neigh_op_bot_0')
// (22, 15, 'neigh_op_tnl_0')
// (22, 16, 'neigh_op_lft_0')
// (22, 17, 'neigh_op_bnl_0')

wire n2844;
// (20, 15, 'neigh_op_tnr_1')
// (20, 16, 'neigh_op_rgt_1')
// (20, 17, 'neigh_op_bnr_1')
// (21, 15, 'neigh_op_top_1')
// (21, 16, 'local_g1_1')
// (21, 16, 'lutff_0/in_2')
// (21, 16, 'lutff_1/out')
// (21, 17, 'neigh_op_bot_1')
// (22, 15, 'neigh_op_tnl_1')
// (22, 16, 'neigh_op_lft_1')
// (22, 17, 'neigh_op_bnl_1')

wire n2845;
// (20, 15, 'neigh_op_tnr_3')
// (20, 16, 'neigh_op_rgt_3')
// (20, 17, 'neigh_op_bnr_3')
// (21, 15, 'neigh_op_top_3')
// (21, 16, 'local_g2_3')
// (21, 16, 'lutff_0/in_3')
// (21, 16, 'lutff_3/out')
// (21, 17, 'neigh_op_bot_3')
// (22, 15, 'neigh_op_tnl_3')
// (22, 16, 'neigh_op_lft_3')
// (22, 17, 'neigh_op_bnl_3')

wire n2846;
// (20, 15, 'neigh_op_tnr_4')
// (20, 16, 'neigh_op_rgt_4')
// (20, 17, 'neigh_op_bnr_4')
// (21, 15, 'neigh_op_top_4')
// (21, 16, 'local_g3_4')
// (21, 16, 'lutff_3/in_2')
// (21, 16, 'lutff_4/out')
// (21, 17, 'neigh_op_bot_4')
// (22, 15, 'neigh_op_tnl_4')
// (22, 16, 'neigh_op_lft_4')
// (22, 17, 'neigh_op_bnl_4')

reg n2847 = 0;
// (20, 15, 'neigh_op_tnr_7')
// (20, 16, 'neigh_op_rgt_7')
// (20, 17, 'neigh_op_bnr_7')
// (21, 15, 'neigh_op_top_7')
// (21, 16, 'local_g2_7')
// (21, 16, 'lutff_4/in_1')
// (21, 16, 'lutff_7/out')
// (21, 17, 'neigh_op_bot_7')
// (22, 15, 'neigh_op_tnl_7')
// (22, 16, 'neigh_op_lft_7')
// (22, 17, 'neigh_op_bnl_7')

wire n2848;
// (20, 15, 'sp4_r_v_b_41')
// (20, 16, 'sp4_r_v_b_28')
// (20, 17, 'sp4_r_v_b_17')
// (20, 18, 'sp4_r_v_b_4')
// (20, 19, 'sp4_r_v_b_36')
// (20, 20, 'neigh_op_tnr_6')
// (20, 20, 'sp4_r_v_b_25')
// (20, 21, 'neigh_op_rgt_6')
// (20, 21, 'sp4_r_v_b_12')
// (20, 22, 'local_g0_6')
// (20, 22, 'lutff_4/in_2')
// (20, 22, 'neigh_op_bnr_6')
// (20, 22, 'sp4_r_v_b_1')
// (21, 14, 'sp4_v_t_41')
// (21, 15, 'sp4_v_b_41')
// (21, 16, 'sp4_v_b_28')
// (21, 17, 'local_g1_1')
// (21, 17, 'lutff_1/in_3')
// (21, 17, 'lutff_6/in_2')
// (21, 17, 'sp4_v_b_17')
// (21, 18, 'sp4_v_b_4')
// (21, 18, 'sp4_v_t_36')
// (21, 19, 'sp4_r_v_b_37')
// (21, 19, 'sp4_v_b_36')
// (21, 20, 'neigh_op_top_6')
// (21, 20, 'sp4_r_v_b_24')
// (21, 20, 'sp4_v_b_25')
// (21, 21, 'local_g3_6')
// (21, 21, 'lutff_3/in_2')
// (21, 21, 'lutff_6/out')
// (21, 21, 'sp4_r_v_b_13')
// (21, 21, 'sp4_v_b_12')
// (21, 22, 'neigh_op_bot_6')
// (21, 22, 'sp4_r_v_b_0')
// (21, 22, 'sp4_v_b_1')
// (22, 18, 'local_g0_0')
// (22, 18, 'lutff_3/in_1')
// (22, 18, 'sp4_h_r_0')
// (22, 18, 'sp4_v_t_37')
// (22, 19, 'sp4_v_b_37')
// (22, 20, 'local_g2_6')
// (22, 20, 'lutff_3/in_1')
// (22, 20, 'neigh_op_tnl_6')
// (22, 20, 'sp4_v_b_24')
// (22, 21, 'local_g1_6')
// (22, 21, 'lutff_7/in_0')
// (22, 21, 'neigh_op_lft_6')
// (22, 21, 'sp4_v_b_13')
// (22, 22, 'local_g3_6')
// (22, 22, 'lutff_7/in_0')
// (22, 22, 'neigh_op_bnl_6')
// (22, 22, 'sp4_v_b_0')
// (23, 18, 'sp4_h_r_13')
// (24, 18, 'sp4_h_r_24')
// (25, 18, 'sp4_h_r_37')

wire n2849;
// (20, 16, 'neigh_op_tnr_3')
// (20, 17, 'neigh_op_rgt_3')
// (20, 18, 'local_g1_3')
// (20, 18, 'lutff_6/in_0')
// (20, 18, 'neigh_op_bnr_3')
// (21, 16, 'neigh_op_top_3')
// (21, 17, 'lutff_3/out')
// (21, 18, 'neigh_op_bot_3')
// (22, 16, 'neigh_op_tnl_3')
// (22, 17, 'neigh_op_lft_3')
// (22, 18, 'neigh_op_bnl_3')

wire n2850;
// (20, 16, 'neigh_op_tnr_4')
// (20, 17, 'neigh_op_rgt_4')
// (20, 18, 'neigh_op_bnr_4')
// (21, 16, 'neigh_op_top_4')
// (21, 17, 'local_g1_4')
// (21, 17, 'lutff_3/in_2')
// (21, 17, 'lutff_4/out')
// (21, 18, 'neigh_op_bot_4')
// (22, 16, 'neigh_op_tnl_4')
// (22, 17, 'neigh_op_lft_4')
// (22, 18, 'neigh_op_bnl_4')

wire n2851;
// (20, 16, 'neigh_op_tnr_5')
// (20, 17, 'neigh_op_rgt_5')
// (20, 18, 'neigh_op_bnr_5')
// (21, 16, 'neigh_op_top_5')
// (21, 17, 'local_g2_5')
// (21, 17, 'lutff_3/in_0')
// (21, 17, 'lutff_5/out')
// (21, 18, 'neigh_op_bot_5')
// (22, 16, 'neigh_op_tnl_5')
// (22, 17, 'neigh_op_lft_5')
// (22, 18, 'neigh_op_bnl_5')

wire n2852;
// (20, 16, 'neigh_op_tnr_6')
// (20, 17, 'neigh_op_rgt_6')
// (20, 17, 'sp4_r_v_b_44')
// (20, 18, 'neigh_op_bnr_6')
// (20, 18, 'sp4_r_v_b_33')
// (20, 19, 'sp4_r_v_b_20')
// (20, 20, 'sp4_r_v_b_9')
// (21, 16, 'local_g0_2')
// (21, 16, 'lutff_global/cen')
// (21, 16, 'neigh_op_top_6')
// (21, 16, 'sp4_h_r_2')
// (21, 16, 'sp4_v_t_44')
// (21, 17, 'lutff_6/out')
// (21, 17, 'sp4_v_b_44')
// (21, 18, 'neigh_op_bot_6')
// (21, 18, 'sp4_v_b_33')
// (21, 19, 'sp4_v_b_20')
// (21, 20, 'sp4_v_b_9')
// (22, 16, 'neigh_op_tnl_6')
// (22, 16, 'sp4_h_r_15')
// (22, 17, 'neigh_op_lft_6')
// (22, 18, 'neigh_op_bnl_6')
// (23, 16, 'sp4_h_r_26')
// (24, 16, 'sp4_h_r_39')
// (25, 16, 'sp4_h_l_39')

reg n2853 = 0;
// (20, 16, 'neigh_op_tnr_7')
// (20, 17, 'neigh_op_rgt_7')
// (20, 18, 'neigh_op_bnr_7')
// (21, 16, 'neigh_op_top_7')
// (21, 17, 'local_g3_7')
// (21, 17, 'lutff_4/in_0')
// (21, 17, 'lutff_7/out')
// (21, 18, 'neigh_op_bot_7')
// (22, 16, 'neigh_op_tnl_7')
// (22, 17, 'neigh_op_lft_7')
// (22, 18, 'neigh_op_bnl_7')

reg n2854 = 0;
// (20, 16, 'sp4_h_r_9')
// (21, 16, 'local_g0_4')
// (21, 16, 'lutff_3/in_1')
// (21, 16, 'sp4_h_r_20')
// (22, 15, 'neigh_op_tnr_6')
// (22, 16, 'neigh_op_rgt_6')
// (22, 16, 'sp4_h_r_33')
// (22, 17, 'neigh_op_bnr_6')
// (23, 15, 'neigh_op_top_6')
// (23, 16, 'lutff_6/out')
// (23, 16, 'sp4_h_r_44')
// (23, 17, 'neigh_op_bot_6')
// (24, 15, 'neigh_op_tnl_6')
// (24, 16, 'neigh_op_lft_6')
// (24, 16, 'sp4_h_l_44')
// (24, 17, 'neigh_op_bnl_6')

wire n2855;
// (20, 16, 'sp4_r_v_b_43')
// (20, 17, 'local_g1_6')
// (20, 17, 'lutff_7/in_2')
// (20, 17, 'sp4_r_v_b_30')
// (20, 18, 'neigh_op_tnr_3')
// (20, 18, 'sp4_r_v_b_19')
// (20, 19, 'neigh_op_rgt_3')
// (20, 19, 'sp4_r_v_b_6')
// (20, 20, 'local_g1_3')
// (20, 20, 'lutff_0/in_2')
// (20, 20, 'neigh_op_bnr_3')
// (21, 15, 'sp4_v_t_43')
// (21, 16, 'sp4_r_v_b_42')
// (21, 16, 'sp4_v_b_43')
// (21, 17, 'sp4_r_v_b_31')
// (21, 17, 'sp4_v_b_30')
// (21, 18, 'neigh_op_top_3')
// (21, 18, 'sp4_r_v_b_18')
// (21, 18, 'sp4_v_b_19')
// (21, 19, 'local_g3_3')
// (21, 19, 'lutff_3/out')
// (21, 19, 'lutff_7/in_1')
// (21, 19, 'sp4_r_v_b_7')
// (21, 19, 'sp4_v_b_6')
// (21, 20, 'local_g0_3')
// (21, 20, 'lutff_5/in_2')
// (21, 20, 'neigh_op_bot_3')
// (22, 15, 'sp4_v_t_42')
// (22, 16, 'sp4_v_b_42')
// (22, 17, 'local_g2_7')
// (22, 17, 'lutff_1/in_2')
// (22, 17, 'lutff_6/in_1')
// (22, 17, 'sp4_v_b_31')
// (22, 18, 'local_g2_3')
// (22, 18, 'lutff_0/in_3')
// (22, 18, 'neigh_op_tnl_3')
// (22, 18, 'sp4_v_b_18')
// (22, 19, 'neigh_op_lft_3')
// (22, 19, 'sp4_v_b_7')
// (22, 20, 'local_g2_3')
// (22, 20, 'lutff_4/in_3')
// (22, 20, 'neigh_op_bnl_3')

wire n2856;
// (20, 17, 'local_g1_3')
// (20, 17, 'lutff_5/in_1')
// (20, 17, 'sp4_h_r_11')
// (21, 17, 'sp4_h_r_22')
// (22, 16, 'neigh_op_tnr_7')
// (22, 17, 'neigh_op_rgt_7')
// (22, 17, 'sp4_h_r_35')
// (22, 18, 'neigh_op_bnr_7')
// (23, 16, 'neigh_op_top_7')
// (23, 17, 'lutff_7/out')
// (23, 17, 'sp4_h_r_46')
// (23, 18, 'neigh_op_bot_7')
// (24, 16, 'neigh_op_tnl_7')
// (24, 17, 'neigh_op_lft_7')
// (24, 17, 'sp4_h_l_46')
// (24, 18, 'neigh_op_bnl_7')

reg n2857 = 0;
// (20, 17, 'neigh_op_tnr_0')
// (20, 18, 'neigh_op_rgt_0')
// (20, 19, 'neigh_op_bnr_0')
// (21, 17, 'local_g1_0')
// (21, 17, 'lutff_5/in_2')
// (21, 17, 'neigh_op_top_0')
// (21, 18, 'lutff_0/out')
// (21, 19, 'neigh_op_bot_0')
// (22, 17, 'neigh_op_tnl_0')
// (22, 18, 'neigh_op_lft_0')
// (22, 19, 'neigh_op_bnl_0')

wire n2858;
// (20, 17, 'neigh_op_tnr_3')
// (20, 18, 'local_g3_3')
// (20, 18, 'lutff_1/in_3')
// (20, 18, 'neigh_op_rgt_3')
// (20, 19, 'neigh_op_bnr_3')
// (21, 17, 'neigh_op_top_3')
// (21, 18, 'lutff_3/out')
// (21, 19, 'neigh_op_bot_3')
// (22, 17, 'neigh_op_tnl_3')
// (22, 18, 'neigh_op_lft_3')
// (22, 19, 'neigh_op_bnl_3')

wire n2859;
// (20, 17, 'sp4_h_r_10')
// (21, 16, 'neigh_op_tnr_1')
// (21, 17, 'neigh_op_rgt_1')
// (21, 17, 'sp4_h_r_23')
// (21, 18, 'neigh_op_bnr_1')
// (22, 16, 'neigh_op_top_1')
// (22, 17, 'lutff_1/out')
// (22, 17, 'sp4_h_r_34')
// (22, 18, 'neigh_op_bot_1')
// (23, 14, 'sp4_r_v_b_43')
// (23, 15, 'sp4_r_v_b_30')
// (23, 16, 'local_g3_3')
// (23, 16, 'lutff_global/cen')
// (23, 16, 'neigh_op_tnl_1')
// (23, 16, 'sp4_r_v_b_19')
// (23, 17, 'neigh_op_lft_1')
// (23, 17, 'sp4_h_r_47')
// (23, 17, 'sp4_r_v_b_6')
// (23, 18, 'neigh_op_bnl_1')
// (24, 13, 'sp4_v_t_43')
// (24, 14, 'sp4_v_b_43')
// (24, 15, 'sp4_v_b_30')
// (24, 16, 'sp4_v_b_19')
// (24, 17, 'sp4_h_l_47')
// (24, 17, 'sp4_h_r_6')
// (24, 17, 'sp4_v_b_6')
// (25, 17, 'sp4_h_r_19')

reg n2860 = 0;
// (20, 18, 'neigh_op_tnr_4')
// (20, 19, 'neigh_op_rgt_4')
// (20, 20, 'neigh_op_bnr_4')
// (21, 18, 'neigh_op_top_4')
// (21, 19, 'lutff_4/out')
// (21, 20, 'local_g1_4')
// (21, 20, 'lutff_2/in_1')
// (21, 20, 'neigh_op_bot_4')
// (22, 18, 'neigh_op_tnl_4')
// (22, 19, 'neigh_op_lft_4')
// (22, 20, 'neigh_op_bnl_4')

wire n2861;
// (20, 18, 'neigh_op_tnr_7')
// (20, 19, 'neigh_op_rgt_7')
// (20, 19, 'sp4_h_r_3')
// (20, 19, 'sp4_h_r_6')
// (20, 20, 'neigh_op_bnr_7')
// (21, 18, 'neigh_op_top_7')
// (21, 19, 'local_g1_3')
// (21, 19, 'lutff_7/out')
// (21, 19, 'lutff_global/cen')
// (21, 19, 'sp4_h_r_14')
// (21, 19, 'sp4_h_r_19')
// (21, 20, 'neigh_op_bot_7')
// (22, 18, 'neigh_op_tnl_7')
// (22, 19, 'neigh_op_lft_7')
// (22, 19, 'sp4_h_r_27')
// (22, 19, 'sp4_h_r_30')
// (22, 20, 'neigh_op_bnl_7')
// (23, 19, 'sp4_h_r_38')
// (23, 19, 'sp4_h_r_43')
// (24, 19, 'sp4_h_l_38')
// (24, 19, 'sp4_h_l_43')
// (24, 19, 'sp4_h_r_3')
// (25, 19, 'sp4_h_r_14')

wire n2862;
// (20, 18, 'sp4_h_r_8')
// (21, 17, 'neigh_op_tnr_0')
// (21, 18, 'neigh_op_rgt_0')
// (21, 18, 'sp4_h_r_21')
// (21, 19, 'neigh_op_bnr_0')
// (22, 17, 'neigh_op_top_0')
// (22, 18, 'lutff_0/out')
// (22, 18, 'sp4_h_r_32')
// (22, 19, 'neigh_op_bot_0')
// (23, 17, 'neigh_op_tnl_0')
// (23, 18, 'neigh_op_lft_0')
// (23, 18, 'sp4_h_r_45')
// (23, 19, 'neigh_op_bnl_0')
// (24, 18, 'local_g1_3')
// (24, 18, 'lutff_global/cen')
// (24, 18, 'sp4_h_l_45')
// (24, 18, 'sp4_h_r_11')
// (25, 18, 'sp4_h_r_22')

wire n2863;
// (20, 19, 'neigh_op_tnr_2')
// (20, 20, 'local_g3_2')
// (20, 20, 'lutff_3/in_2')
// (20, 20, 'neigh_op_rgt_2')
// (20, 21, 'neigh_op_bnr_2')
// (21, 19, 'neigh_op_top_2')
// (21, 20, 'lutff_2/out')
// (21, 21, 'neigh_op_bot_2')
// (22, 19, 'neigh_op_tnl_2')
// (22, 20, 'neigh_op_lft_2')
// (22, 21, 'neigh_op_bnl_2')

wire n2864;
// (20, 19, 'neigh_op_tnr_4')
// (20, 20, 'neigh_op_rgt_4')
// (20, 21, 'neigh_op_bnr_4')
// (21, 19, 'neigh_op_top_4')
// (21, 20, 'local_g3_4')
// (21, 20, 'lutff_4/out')
// (21, 20, 'lutff_7/in_2')
// (21, 21, 'neigh_op_bot_4')
// (22, 19, 'neigh_op_tnl_4')
// (22, 20, 'neigh_op_lft_4')
// (22, 21, 'neigh_op_bnl_4')

wire n2865;
// (20, 19, 'neigh_op_tnr_5')
// (20, 20, 'neigh_op_rgt_5')
// (20, 21, 'neigh_op_bnr_5')
// (21, 19, 'neigh_op_top_5')
// (21, 20, 'local_g0_2')
// (21, 20, 'lutff_5/out')
// (21, 20, 'lutff_global/cen')
// (21, 20, 'sp4_h_r_10')
// (21, 21, 'neigh_op_bot_5')
// (22, 19, 'neigh_op_tnl_5')
// (22, 20, 'neigh_op_lft_5')
// (22, 20, 'sp4_h_r_23')
// (22, 21, 'neigh_op_bnl_5')
// (23, 20, 'sp4_h_r_34')
// (24, 20, 'sp4_h_r_47')
// (25, 20, 'sp4_h_l_47')

reg n2866 = 0;
// (20, 19, 'neigh_op_tnr_6')
// (20, 20, 'neigh_op_rgt_6')
// (20, 21, 'neigh_op_bnr_6')
// (21, 19, 'neigh_op_top_6')
// (21, 20, 'local_g2_6')
// (21, 20, 'lutff_4/in_2')
// (21, 20, 'lutff_6/out')
// (21, 21, 'neigh_op_bot_6')
// (22, 19, 'neigh_op_tnl_6')
// (22, 20, 'neigh_op_lft_6')
// (22, 21, 'neigh_op_bnl_6')

wire n2867;
// (20, 19, 'neigh_op_tnr_7')
// (20, 20, 'local_g2_7')
// (20, 20, 'lutff_1/in_2')
// (20, 20, 'neigh_op_rgt_7')
// (20, 21, 'neigh_op_bnr_7')
// (21, 19, 'neigh_op_top_7')
// (21, 20, 'lutff_7/out')
// (21, 21, 'neigh_op_bot_7')
// (22, 19, 'neigh_op_tnl_7')
// (22, 20, 'neigh_op_lft_7')
// (22, 21, 'neigh_op_bnl_7')

wire n2868;
// (20, 19, 'sp4_h_r_8')
// (21, 18, 'neigh_op_tnr_0')
// (21, 19, 'neigh_op_rgt_0')
// (21, 19, 'sp4_h_r_21')
// (21, 20, 'neigh_op_bnr_0')
// (22, 18, 'neigh_op_top_0')
// (22, 19, 'lutff_0/out')
// (22, 19, 'sp4_h_r_32')
// (22, 20, 'neigh_op_bot_0')
// (23, 18, 'neigh_op_tnl_0')
// (23, 19, 'neigh_op_lft_0')
// (23, 19, 'sp4_h_r_45')
// (23, 20, 'neigh_op_bnl_0')
// (24, 19, 'local_g1_3')
// (24, 19, 'lutff_global/cen')
// (24, 19, 'sp4_h_l_45')
// (24, 19, 'sp4_h_r_11')
// (25, 19, 'sp4_h_r_22')

wire n2869;
// (20, 20, 'local_g3_5')
// (20, 20, 'lutff_1/in_3')
// (20, 20, 'neigh_op_tnr_5')
// (20, 21, 'neigh_op_rgt_5')
// (20, 22, 'neigh_op_bnr_5')
// (21, 20, 'neigh_op_top_5')
// (21, 21, 'lutff_5/out')
// (21, 22, 'neigh_op_bot_5')
// (22, 20, 'neigh_op_tnl_5')
// (22, 21, 'neigh_op_lft_5')
// (22, 22, 'neigh_op_bnl_5')

reg n2870 = 0;
// (20, 20, 'neigh_op_tnr_0')
// (20, 21, 'neigh_op_rgt_0')
// (20, 22, 'neigh_op_bnr_0')
// (21, 20, 'neigh_op_top_0')
// (21, 21, 'local_g3_0')
// (21, 21, 'lutff_0/out')
// (21, 21, 'lutff_4/in_1')
// (21, 22, 'neigh_op_bot_0')
// (22, 20, 'neigh_op_tnl_0')
// (22, 21, 'neigh_op_lft_0')
// (22, 22, 'neigh_op_bnl_0')

wire n2871;
// (20, 20, 'neigh_op_tnr_1')
// (20, 21, 'neigh_op_rgt_1')
// (20, 22, 'neigh_op_bnr_1')
// (21, 20, 'neigh_op_top_1')
// (21, 21, 'local_g3_1')
// (21, 21, 'lutff_1/out')
// (21, 21, 'lutff_5/in_1')
// (21, 22, 'neigh_op_bot_1')
// (22, 20, 'neigh_op_tnl_1')
// (22, 21, 'neigh_op_lft_1')
// (22, 22, 'neigh_op_bnl_1')

wire n2872;
// (20, 20, 'neigh_op_tnr_2')
// (20, 21, 'neigh_op_rgt_2')
// (20, 22, 'neigh_op_bnr_2')
// (21, 20, 'neigh_op_top_2')
// (21, 21, 'local_g3_2')
// (21, 21, 'lutff_2/out')
// (21, 21, 'lutff_5/in_2')
// (21, 22, 'neigh_op_bot_2')
// (22, 20, 'neigh_op_tnl_2')
// (22, 21, 'neigh_op_lft_2')
// (22, 22, 'neigh_op_bnl_2')

wire n2873;
// (20, 20, 'neigh_op_tnr_3')
// (20, 21, 'neigh_op_rgt_3')
// (20, 22, 'neigh_op_bnr_3')
// (21, 20, 'neigh_op_top_3')
// (21, 21, 'local_g1_3')
// (21, 21, 'lutff_3/out')
// (21, 21, 'lutff_global/cen')
// (21, 22, 'neigh_op_bot_3')
// (22, 20, 'neigh_op_tnl_3')
// (22, 21, 'neigh_op_lft_3')
// (22, 22, 'neigh_op_bnl_3')

wire n2874;
// (20, 20, 'neigh_op_tnr_4')
// (20, 21, 'neigh_op_rgt_4')
// (20, 22, 'neigh_op_bnr_4')
// (21, 20, 'local_g0_4')
// (21, 20, 'lutff_2/in_0')
// (21, 20, 'neigh_op_top_4')
// (21, 21, 'lutff_4/out')
// (21, 22, 'neigh_op_bot_4')
// (22, 20, 'neigh_op_tnl_4')
// (22, 21, 'neigh_op_lft_4')
// (22, 22, 'neigh_op_bnl_4')

wire n2875;
// (20, 20, 'neigh_op_tnr_7')
// (20, 21, 'neigh_op_rgt_7')
// (20, 22, 'neigh_op_bnr_7')
// (21, 20, 'neigh_op_top_7')
// (21, 21, 'local_g2_7')
// (21, 21, 'lutff_2/in_3')
// (21, 21, 'lutff_7/out')
// (21, 22, 'neigh_op_bot_7')
// (22, 20, 'neigh_op_tnl_7')
// (22, 21, 'neigh_op_lft_7')
// (22, 22, 'neigh_op_bnl_7')

wire n2876;
// (20, 20, 'sp4_h_r_4')
// (21, 19, 'neigh_op_tnr_6')
// (21, 20, 'neigh_op_rgt_6')
// (21, 20, 'sp4_h_r_17')
// (21, 21, 'neigh_op_bnr_6')
// (22, 19, 'neigh_op_top_6')
// (22, 20, 'lutff_6/out')
// (22, 20, 'sp4_h_r_28')
// (22, 21, 'neigh_op_bot_6')
// (23, 17, 'sp4_r_v_b_47')
// (23, 18, 'sp4_r_v_b_34')
// (23, 19, 'neigh_op_tnl_6')
// (23, 19, 'sp4_r_v_b_23')
// (23, 20, 'neigh_op_lft_6')
// (23, 20, 'sp4_h_r_41')
// (23, 20, 'sp4_r_v_b_10')
// (23, 21, 'neigh_op_bnl_6')
// (24, 16, 'sp4_v_t_47')
// (24, 17, 'sp4_v_b_47')
// (24, 18, 'sp4_v_b_34')
// (24, 19, 'sp4_v_b_23')
// (24, 20, 'local_g0_2')
// (24, 20, 'lutff_global/cen')
// (24, 20, 'sp4_h_l_41')
// (24, 20, 'sp4_v_b_10')

wire n2877;
// (20, 20, 'sp4_h_r_6')
// (21, 20, 'local_g1_3')
// (21, 20, 'lutff_7/in_1')
// (21, 20, 'sp4_h_r_19')
// (22, 18, 'neigh_op_tnr_1')
// (22, 19, 'neigh_op_rgt_1')
// (22, 20, 'neigh_op_bnr_1')
// (22, 20, 'sp4_h_r_30')
// (23, 17, 'sp4_r_v_b_43')
// (23, 18, 'neigh_op_top_1')
// (23, 18, 'sp4_r_v_b_30')
// (23, 19, 'lutff_1/out')
// (23, 19, 'sp4_r_v_b_19')
// (23, 20, 'neigh_op_bot_1')
// (23, 20, 'sp4_h_r_43')
// (23, 20, 'sp4_r_v_b_6')
// (24, 16, 'sp4_v_t_43')
// (24, 17, 'sp4_v_b_43')
// (24, 18, 'neigh_op_tnl_1')
// (24, 18, 'sp4_v_b_30')
// (24, 19, 'neigh_op_lft_1')
// (24, 19, 'sp4_v_b_19')
// (24, 20, 'neigh_op_bnl_1')
// (24, 20, 'sp4_h_l_43')
// (24, 20, 'sp4_v_b_6')

reg n2878 = 0;
// (20, 20, 'sp4_r_v_b_39')
// (20, 21, 'sp4_r_v_b_26')
// (20, 22, 'neigh_op_tnr_1')
// (20, 22, 'sp4_r_v_b_15')
// (20, 23, 'neigh_op_rgt_1')
// (20, 23, 'sp4_r_v_b_2')
// (20, 24, 'neigh_op_bnr_1')
// (21, 19, 'sp4_v_t_39')
// (21, 20, 'sp4_v_b_39')
// (21, 21, 'local_g2_2')
// (21, 21, 'lutff_7/in_1')
// (21, 21, 'sp4_v_b_26')
// (21, 22, 'neigh_op_top_1')
// (21, 22, 'sp4_v_b_15')
// (21, 23, 'lutff_1/out')
// (21, 23, 'sp4_v_b_2')
// (21, 24, 'neigh_op_bot_1')
// (22, 22, 'neigh_op_tnl_1')
// (22, 23, 'neigh_op_lft_1')
// (22, 24, 'neigh_op_bnl_1')

wire n2879;
// (20, 20, 'sp4_r_v_b_45')
// (20, 21, 'sp4_r_v_b_32')
// (20, 22, 'neigh_op_tnr_4')
// (20, 22, 'sp4_r_v_b_21')
// (20, 23, 'neigh_op_rgt_4')
// (20, 23, 'sp4_r_v_b_8')
// (20, 24, 'neigh_op_bnr_4')
// (21, 19, 'sp4_v_t_45')
// (21, 20, 'sp4_v_b_45')
// (21, 21, 'sp4_v_b_32')
// (21, 22, 'neigh_op_top_4')
// (21, 22, 'sp4_v_b_21')
// (21, 23, 'local_g0_2')
// (21, 23, 'lutff_4/out')
// (21, 23, 'lutff_global/cen')
// (21, 23, 'sp4_h_r_2')
// (21, 23, 'sp4_v_b_8')
// (21, 24, 'neigh_op_bot_4')
// (22, 22, 'neigh_op_tnl_4')
// (22, 23, 'neigh_op_lft_4')
// (22, 23, 'sp4_h_r_15')
// (22, 24, 'neigh_op_bnl_4')
// (23, 23, 'sp4_h_r_26')
// (24, 23, 'sp4_h_r_39')
// (25, 23, 'sp4_h_l_39')

reg n2880 = 0;
// (20, 21, 'neigh_op_tnr_3')
// (20, 22, 'neigh_op_rgt_3')
// (20, 23, 'neigh_op_bnr_3')
// (21, 21, 'local_g0_3')
// (21, 21, 'lutff_1/in_2')
// (21, 21, 'neigh_op_top_3')
// (21, 22, 'lutff_3/out')
// (21, 23, 'neigh_op_bot_3')
// (22, 21, 'neigh_op_tnl_3')
// (22, 22, 'neigh_op_lft_3')
// (22, 23, 'neigh_op_bnl_3')

wire n2881;
// (20, 21, 'neigh_op_tnr_5')
// (20, 22, 'neigh_op_rgt_5')
// (20, 23, 'neigh_op_bnr_5')
// (21, 21, 'neigh_op_top_5')
// (21, 22, 'local_g0_2')
// (21, 22, 'lutff_5/out')
// (21, 22, 'lutff_global/cen')
// (21, 22, 'sp4_h_r_10')
// (21, 23, 'neigh_op_bot_5')
// (22, 21, 'neigh_op_tnl_5')
// (22, 22, 'neigh_op_lft_5')
// (22, 22, 'sp4_h_r_23')
// (22, 23, 'neigh_op_bnl_5')
// (23, 22, 'sp4_h_r_34')
// (24, 22, 'sp4_h_r_47')
// (25, 22, 'sp4_h_l_47')

wire n2882;
// (20, 21, 'sp4_h_r_10')
// (20, 21, 'sp4_h_r_6')
// (21, 20, 'neigh_op_tnr_7')
// (21, 21, 'neigh_op_rgt_7')
// (21, 21, 'sp4_h_r_19')
// (21, 21, 'sp4_h_r_23')
// (21, 22, 'neigh_op_bnr_7')
// (22, 20, 'neigh_op_top_7')
// (22, 21, 'local_g2_2')
// (22, 21, 'lutff_7/out')
// (22, 21, 'lutff_global/cen')
// (22, 21, 'sp4_h_r_30')
// (22, 21, 'sp4_h_r_34')
// (22, 22, 'neigh_op_bot_7')
// (23, 20, 'neigh_op_tnl_7')
// (23, 21, 'neigh_op_lft_7')
// (23, 21, 'sp4_h_r_43')
// (23, 21, 'sp4_h_r_47')
// (23, 22, 'neigh_op_bnl_7')
// (24, 21, 'sp4_h_l_43')
// (24, 21, 'sp4_h_l_47')
// (24, 21, 'sp4_h_r_2')
// (25, 21, 'sp4_h_r_15')

reg n2883 = 0;
// (20, 22, 'local_g1_0')
// (20, 22, 'lutff_7/in_0')
// (20, 22, 'sp4_h_r_0')
// (21, 21, 'neigh_op_tnr_4')
// (21, 22, 'neigh_op_rgt_4')
// (21, 22, 'sp4_h_r_13')
// (21, 23, 'neigh_op_bnr_4')
// (22, 21, 'neigh_op_top_4')
// (22, 22, 'lutff_4/out')
// (22, 22, 'sp4_h_r_24')
// (22, 23, 'neigh_op_bot_4')
// (23, 21, 'neigh_op_tnl_4')
// (23, 22, 'neigh_op_lft_4')
// (23, 22, 'sp4_h_r_37')
// (23, 23, 'neigh_op_bnl_4')
// (24, 22, 'sp4_h_l_37')

wire n2884;
// (20, 22, 'neigh_op_tnr_7')
// (20, 22, 'sp4_r_v_b_43')
// (20, 23, 'neigh_op_rgt_7')
// (20, 23, 'sp4_r_v_b_30')
// (20, 24, 'neigh_op_bnr_7')
// (20, 24, 'sp4_r_v_b_19')
// (20, 25, 'sp4_r_v_b_6')
// (21, 21, 'sp4_v_t_43')
// (21, 22, 'neigh_op_top_7')
// (21, 22, 'sp4_v_b_43')
// (21, 23, 'lutff_7/out')
// (21, 23, 'sp4_v_b_30')
// (21, 24, 'local_g1_3')
// (21, 24, 'lutff_global/cen')
// (21, 24, 'neigh_op_bot_7')
// (21, 24, 'sp4_v_b_19')
// (21, 25, 'sp4_v_b_6')
// (22, 22, 'neigh_op_tnl_7')
// (22, 23, 'neigh_op_lft_7')
// (22, 24, 'neigh_op_bnl_7')

reg n2885 = 0;
// (20, 22, 'sp4_r_v_b_36')
// (20, 23, 'neigh_op_tnr_6')
// (20, 23, 'sp4_r_v_b_25')
// (20, 24, 'neigh_op_rgt_6')
// (20, 24, 'sp4_r_v_b_12')
// (20, 25, 'neigh_op_bnr_6')
// (20, 25, 'sp4_r_v_b_1')
// (21, 21, 'local_g0_1')
// (21, 21, 'lutff_1/in_0')
// (21, 21, 'sp4_h_r_1')
// (21, 21, 'sp4_v_t_36')
// (21, 22, 'sp4_v_b_36')
// (21, 23, 'neigh_op_top_6')
// (21, 23, 'sp4_v_b_25')
// (21, 24, 'lutff_6/out')
// (21, 24, 'sp4_v_b_12')
// (21, 25, 'neigh_op_bot_6')
// (21, 25, 'sp4_v_b_1')
// (22, 21, 'sp4_h_r_12')
// (22, 23, 'neigh_op_tnl_6')
// (22, 24, 'neigh_op_lft_6')
// (22, 25, 'neigh_op_bnl_6')
// (23, 21, 'sp4_h_r_25')
// (24, 21, 'sp4_h_r_36')
// (25, 21, 'sp4_h_l_36')

wire n2886;
// (21, 1, 'neigh_op_tnr_0')
// (21, 2, 'neigh_op_rgt_0')
// (21, 3, 'neigh_op_bnr_0')
// (22, 1, 'neigh_op_top_0')
// (22, 2, 'local_g0_0')
// (22, 2, 'local_g3_0')
// (22, 2, 'lutff_0/out')
// (22, 2, 'lutff_4/in_2')
// (22, 2, 'lutff_5/in_2')
// (22, 3, 'neigh_op_bot_0')
// (23, 1, 'neigh_op_tnl_0')
// (23, 2, 'neigh_op_lft_0')
// (23, 3, 'neigh_op_bnl_0')

reg n2887 = 0;
// (21, 1, 'neigh_op_tnr_1')
// (21, 2, 'neigh_op_rgt_1')
// (21, 3, 'neigh_op_bnr_1')
// (22, 1, 'neigh_op_top_1')
// (22, 2, 'local_g1_1')
// (22, 2, 'lutff_1/out')
// (22, 2, 'lutff_7/in_3')
// (22, 3, 'neigh_op_bot_1')
// (23, 1, 'neigh_op_tnl_1')
// (23, 2, 'neigh_op_lft_1')
// (23, 3, 'local_g3_1')
// (23, 3, 'lutff_4/in_2')
// (23, 3, 'neigh_op_bnl_1')

wire n2888;
// (21, 1, 'neigh_op_tnr_2')
// (21, 2, 'neigh_op_rgt_2')
// (21, 3, 'neigh_op_bnr_2')
// (22, 1, 'neigh_op_top_2')
// (22, 1, 'sp4_r_v_b_16')
// (22, 2, 'local_g0_2')
// (22, 2, 'local_g1_2')
// (22, 2, 'lutff_2/out')
// (22, 2, 'lutff_4/in_3')
// (22, 2, 'lutff_5/in_3')
// (22, 2, 'sp4_r_v_b_37')
// (22, 2, 'sp4_r_v_b_5')
// (22, 3, 'neigh_op_bot_2')
// (22, 3, 'sp4_r_v_b_24')
// (22, 3, 'sp4_r_v_b_45')
// (22, 4, 'sp4_r_v_b_13')
// (22, 4, 'sp4_r_v_b_32')
// (22, 5, 'sp4_r_v_b_0')
// (22, 5, 'sp4_r_v_b_21')
// (22, 6, 'sp4_r_v_b_8')
// (23, 0, 'span4_vert_16')
// (23, 1, 'neigh_op_tnl_2')
// (23, 1, 'sp4_v_b_16')
// (23, 1, 'sp4_v_t_37')
// (23, 2, 'local_g3_5')
// (23, 2, 'lutff_global/s_r')
// (23, 2, 'neigh_op_lft_2')
// (23, 2, 'sp4_v_b_37')
// (23, 2, 'sp4_v_b_5')
// (23, 2, 'sp4_v_t_45')
// (23, 3, 'local_g3_5')
// (23, 3, 'lutff_global/s_r')
// (23, 3, 'neigh_op_bnl_2')
// (23, 3, 'sp4_v_b_24')
// (23, 3, 'sp4_v_b_45')
// (23, 4, 'sp4_v_b_13')
// (23, 4, 'sp4_v_b_32')
// (23, 5, 'sp4_v_b_0')
// (23, 5, 'sp4_v_b_21')
// (23, 6, 'sp4_v_b_8')

wire n2889;
// (21, 1, 'neigh_op_tnr_3')
// (21, 2, 'local_g3_3')
// (21, 2, 'lutff_0/in_0')
// (21, 2, 'lutff_3/in_1')
// (21, 2, 'lutff_4/in_2')
// (21, 2, 'neigh_op_rgt_3')
// (21, 3, 'neigh_op_bnr_3')
// (22, 1, 'neigh_op_top_3')
// (22, 2, 'local_g2_3')
// (22, 2, 'lutff_1/in_2')
// (22, 2, 'lutff_2/in_1')
// (22, 2, 'lutff_3/out')
// (22, 2, 'lutff_6/in_3')
// (22, 3, 'local_g1_3')
// (22, 3, 'lutff_2/in_2')
// (22, 3, 'lutff_4/in_2')
// (22, 3, 'lutff_6/in_2')
// (22, 3, 'neigh_op_bot_3')
// (23, 1, 'neigh_op_tnl_3')
// (23, 2, 'neigh_op_lft_3')
// (23, 3, 'neigh_op_bnl_3')

reg n2890 = 0;
// (21, 1, 'neigh_op_tnr_4')
// (21, 2, 'neigh_op_rgt_4')
// (21, 3, 'neigh_op_bnr_4')
// (22, 1, 'neigh_op_top_4')
// (22, 2, 'local_g0_4')
// (22, 2, 'local_g1_4')
// (22, 2, 'lutff_3/in_3')
// (22, 2, 'lutff_4/in_1')
// (22, 2, 'lutff_4/out')
// (22, 3, 'neigh_op_bot_4')
// (23, 1, 'neigh_op_tnl_4')
// (23, 2, 'local_g1_4')
// (23, 2, 'lutff_1/in_2')
// (23, 2, 'neigh_op_lft_4')
// (23, 3, 'neigh_op_bnl_4')

reg n2891 = 0;
// (21, 1, 'neigh_op_tnr_5')
// (21, 2, 'neigh_op_rgt_5')
// (21, 3, 'neigh_op_bnr_5')
// (22, 1, 'neigh_op_top_5')
// (22, 2, 'local_g0_5')
// (22, 2, 'lutff_3/in_2')
// (22, 2, 'lutff_5/in_0')
// (22, 2, 'lutff_5/out')
// (22, 3, 'neigh_op_bot_5')
// (23, 1, 'neigh_op_tnl_5')
// (23, 2, 'local_g1_5')
// (23, 2, 'lutff_6/in_2')
// (23, 2, 'neigh_op_lft_5')
// (23, 3, 'neigh_op_bnl_5')

reg n2892 = 0;
// (21, 1, 'neigh_op_tnr_6')
// (21, 2, 'neigh_op_rgt_6')
// (21, 3, 'neigh_op_bnr_6')
// (22, 1, 'neigh_op_top_6')
// (22, 2, 'local_g1_6')
// (22, 2, 'lutff_6/out')
// (22, 2, 'lutff_7/in_2')
// (22, 3, 'neigh_op_bot_6')
// (23, 1, 'neigh_op_tnl_6')
// (23, 2, 'local_g0_6')
// (23, 2, 'lutff_7/in_1')
// (23, 2, 'neigh_op_lft_6')
// (23, 3, 'neigh_op_bnl_6')

wire n2893;
// (21, 1, 'neigh_op_tnr_7')
// (21, 2, 'neigh_op_rgt_7')
// (21, 3, 'neigh_op_bnr_7')
// (22, 1, 'neigh_op_top_7')
// (22, 2, 'local_g1_7')
// (22, 2, 'lutff_3/in_1')
// (22, 2, 'lutff_7/out')
// (22, 3, 'neigh_op_bot_7')
// (23, 1, 'neigh_op_tnl_7')
// (23, 2, 'neigh_op_lft_7')
// (23, 3, 'neigh_op_bnl_7')

reg n2894 = 0;
// (21, 1, 'sp4_r_v_b_32')
// (21, 2, 'sp4_r_v_b_21')
// (21, 3, 'local_g2_0')
// (21, 3, 'lutff_1/in_1')
// (21, 3, 'sp4_r_v_b_8')
// (22, 0, 'span4_vert_32')
// (22, 1, 'sp4_v_b_32')
// (22, 2, 'sp4_v_b_21')
// (22, 3, 'local_g0_0')
// (22, 3, 'lutff_7/in_1')
// (22, 3, 'sp4_h_r_8')
// (22, 3, 'sp4_v_b_8')
// (23, 2, 'neigh_op_tnr_0')
// (23, 3, 'neigh_op_rgt_0')
// (23, 3, 'sp4_h_r_21')
// (23, 4, 'neigh_op_bnr_0')
// (24, 2, 'neigh_op_top_0')
// (24, 3, 'local_g0_0')
// (24, 3, 'lutff_0/in_0')
// (24, 3, 'lutff_0/out')
// (24, 3, 'sp4_h_r_32')
// (24, 4, 'neigh_op_bot_0')
// (25, 2, 'neigh_op_tnl_0')
// (25, 3, 'neigh_op_lft_0')
// (25, 3, 'sp4_h_r_45')
// (25, 4, 'neigh_op_bnl_0')

wire n2895;
// (21, 2, 'neigh_op_tnr_0')
// (21, 3, 'neigh_op_rgt_0')
// (21, 4, 'neigh_op_bnr_0')
// (22, 2, 'local_g1_0')
// (22, 2, 'lutff_3/in_0')
// (22, 2, 'neigh_op_top_0')
// (22, 3, 'lutff_0/out')
// (22, 4, 'neigh_op_bot_0')
// (23, 2, 'neigh_op_tnl_0')
// (23, 3, 'neigh_op_lft_0')
// (23, 4, 'neigh_op_bnl_0')

reg n2896 = 0;
// (21, 2, 'neigh_op_tnr_2')
// (21, 3, 'neigh_op_rgt_2')
// (21, 4, 'neigh_op_bnr_2')
// (22, 2, 'neigh_op_top_2')
// (22, 3, 'local_g2_2')
// (22, 3, 'lutff_0/in_2')
// (22, 3, 'lutff_2/in_0')
// (22, 3, 'lutff_2/out')
// (22, 4, 'neigh_op_bot_2')
// (23, 2, 'neigh_op_tnl_2')
// (23, 3, 'local_g1_2')
// (23, 3, 'lutff_1/in_2')
// (23, 3, 'neigh_op_lft_2')
// (23, 4, 'neigh_op_bnl_2')

reg n2897 = 0;
// (21, 2, 'neigh_op_tnr_4')
// (21, 3, 'neigh_op_rgt_4')
// (21, 4, 'neigh_op_bnr_4')
// (22, 2, 'neigh_op_top_4')
// (22, 3, 'local_g2_4')
// (22, 3, 'local_g3_4')
// (22, 3, 'lutff_0/in_0')
// (22, 3, 'lutff_4/in_1')
// (22, 3, 'lutff_4/out')
// (22, 4, 'neigh_op_bot_4')
// (23, 2, 'neigh_op_tnl_4')
// (23, 3, 'local_g1_4')
// (23, 3, 'lutff_3/in_2')
// (23, 3, 'neigh_op_lft_4')
// (23, 4, 'neigh_op_bnl_4')

wire n2898;
// (21, 2, 'neigh_op_tnr_5')
// (21, 3, 'neigh_op_rgt_5')
// (21, 4, 'neigh_op_bnr_5')
// (22, 2, 'neigh_op_top_5')
// (22, 3, 'lutff_5/out')
// (22, 4, 'local_g0_5')
// (22, 4, 'lutff_2/in_1')
// (22, 4, 'neigh_op_bot_5')
// (23, 2, 'neigh_op_tnl_5')
// (23, 3, 'neigh_op_lft_5')
// (23, 4, 'neigh_op_bnl_5')

reg n2899 = 0;
// (21, 2, 'neigh_op_tnr_6')
// (21, 3, 'neigh_op_rgt_6')
// (21, 4, 'neigh_op_bnr_6')
// (22, 2, 'neigh_op_top_6')
// (22, 3, 'local_g3_6')
// (22, 3, 'lutff_0/in_3')
// (22, 3, 'lutff_6/in_3')
// (22, 3, 'lutff_6/out')
// (22, 4, 'neigh_op_bot_6')
// (23, 2, 'local_g2_6')
// (23, 2, 'lutff_4/in_2')
// (23, 2, 'neigh_op_tnl_6')
// (23, 3, 'neigh_op_lft_6')
// (23, 4, 'neigh_op_bnl_6')

wire n2900;
// (21, 2, 'neigh_op_tnr_7')
// (21, 3, 'neigh_op_rgt_7')
// (21, 4, 'neigh_op_bnr_7')
// (22, 2, 'neigh_op_top_7')
// (22, 3, 'lutff_7/out')
// (22, 4, 'local_g1_7')
// (22, 4, 'lutff_2/in_2')
// (22, 4, 'neigh_op_bot_7')
// (23, 2, 'neigh_op_tnl_7')
// (23, 3, 'neigh_op_lft_7')
// (23, 4, 'neigh_op_bnl_7')

reg n2901 = 0;
// (21, 3, 'local_g0_5')
// (21, 3, 'lutff_0/in_1')
// (21, 3, 'sp4_h_r_5')
// (22, 3, 'local_g1_0')
// (22, 3, 'lutff_5/in_0')
// (22, 3, 'sp4_h_r_16')
// (23, 2, 'neigh_op_tnr_4')
// (23, 3, 'neigh_op_rgt_4')
// (23, 3, 'sp4_h_r_29')
// (23, 4, 'neigh_op_bnr_4')
// (24, 2, 'neigh_op_top_4')
// (24, 3, 'local_g1_4')
// (24, 3, 'lutff_0/in_1')
// (24, 3, 'lutff_4/in_3')
// (24, 3, 'lutff_4/out')
// (24, 3, 'sp4_h_r_40')
// (24, 4, 'neigh_op_bot_4')
// (25, 2, 'neigh_op_tnl_4')
// (25, 3, 'neigh_op_lft_4')
// (25, 3, 'sp4_h_l_40')
// (25, 4, 'neigh_op_bnl_4')

wire n2902;
// (21, 3, 'local_g3_3')
// (21, 3, 'lutff_global/cen')
// (21, 3, 'neigh_op_tnr_3')
// (21, 4, 'local_g3_3')
// (21, 4, 'lutff_global/cen')
// (21, 4, 'neigh_op_rgt_3')
// (21, 5, 'local_g1_3')
// (21, 5, 'lutff_global/cen')
// (21, 5, 'neigh_op_bnr_3')
// (22, 3, 'neigh_op_top_3')
// (22, 4, 'lutff_3/out')
// (22, 4, 'sp4_r_v_b_39')
// (22, 5, 'neigh_op_bot_3')
// (22, 5, 'sp4_r_v_b_26')
// (22, 6, 'sp4_r_v_b_15')
// (22, 7, 'sp4_r_v_b_2')
// (23, 3, 'neigh_op_tnl_3')
// (23, 3, 'sp4_h_r_7')
// (23, 3, 'sp4_v_t_39')
// (23, 4, 'neigh_op_lft_3')
// (23, 4, 'sp4_v_b_39')
// (23, 5, 'neigh_op_bnl_3')
// (23, 5, 'sp4_v_b_26')
// (23, 6, 'sp4_v_b_15')
// (23, 7, 'sp4_v_b_2')
// (24, 3, 'local_g0_2')
// (24, 3, 'lutff_global/cen')
// (24, 3, 'sp4_h_r_18')
// (25, 3, 'sp4_h_r_31')

wire n2903;
// (21, 3, 'lutff_1/cout')
// (21, 3, 'lutff_2/in_3')

wire n2904;
// (21, 3, 'lutff_2/cout')
// (21, 3, 'lutff_3/in_3')

wire n2905;
// (21, 3, 'lutff_3/cout')
// (21, 3, 'lutff_4/in_3')

wire n2906;
// (21, 3, 'lutff_4/cout')
// (21, 3, 'lutff_5/in_3')

wire n2907;
// (21, 3, 'lutff_5/cout')
// (21, 3, 'lutff_6/in_3')

wire n2908;
// (21, 3, 'lutff_6/cout')
// (21, 3, 'lutff_7/in_3')

wire n2909;
// (21, 3, 'lutff_7/cout')
// (21, 4, 'carry_in')
// (21, 4, 'carry_in_mux')
// (21, 4, 'lutff_0/in_3')

wire n2910;
// (21, 3, 'neigh_op_tnr_1')
// (21, 4, 'neigh_op_rgt_1')
// (21, 5, 'neigh_op_bnr_1')
// (22, 3, 'neigh_op_top_1')
// (22, 4, 'lutff_1/out')
// (22, 5, 'local_g1_1')
// (22, 5, 'lutff_3/in_1')
// (22, 5, 'neigh_op_bot_1')
// (23, 3, 'neigh_op_tnl_1')
// (23, 4, 'neigh_op_lft_1')
// (23, 5, 'neigh_op_bnl_1')

wire n2911;
// (21, 3, 'neigh_op_tnr_2')
// (21, 4, 'neigh_op_rgt_2')
// (21, 5, 'neigh_op_bnr_2')
// (22, 3, 'neigh_op_top_2')
// (22, 4, 'lutff_2/out')
// (22, 5, 'local_g0_2')
// (22, 5, 'lutff_7/in_1')
// (22, 5, 'neigh_op_bot_2')
// (23, 3, 'neigh_op_tnl_2')
// (23, 4, 'neigh_op_lft_2')
// (23, 5, 'neigh_op_bnl_2')

wire n2912;
// (21, 3, 'neigh_op_tnr_4')
// (21, 4, 'local_g3_4')
// (21, 4, 'lutff_3/in_2')
// (21, 4, 'neigh_op_rgt_4')
// (21, 5, 'neigh_op_bnr_4')
// (22, 3, 'neigh_op_top_4')
// (22, 4, 'lutff_4/out')
// (22, 5, 'neigh_op_bot_4')
// (23, 3, 'neigh_op_tnl_4')
// (23, 4, 'neigh_op_lft_4')
// (23, 5, 'neigh_op_bnl_4')

wire n2913;
// (21, 3, 'neigh_op_tnr_5')
// (21, 4, 'neigh_op_rgt_5')
// (21, 5, 'neigh_op_bnr_5')
// (22, 3, 'neigh_op_top_5')
// (22, 4, 'local_g2_5')
// (22, 4, 'lutff_2/in_3')
// (22, 4, 'lutff_5/out')
// (22, 5, 'neigh_op_bot_5')
// (23, 3, 'neigh_op_tnl_5')
// (23, 4, 'neigh_op_lft_5')
// (23, 5, 'neigh_op_bnl_5')

wire n2914;
// (21, 3, 'neigh_op_tnr_6')
// (21, 4, 'local_g2_6')
// (21, 4, 'lutff_2/in_2')
// (21, 4, 'neigh_op_rgt_6')
// (21, 5, 'neigh_op_bnr_6')
// (22, 3, 'neigh_op_top_6')
// (22, 4, 'lutff_6/out')
// (22, 5, 'neigh_op_bot_6')
// (23, 3, 'neigh_op_tnl_6')
// (23, 4, 'neigh_op_lft_6')
// (23, 5, 'neigh_op_bnl_6')

wire n2915;
// (21, 3, 'neigh_op_tnr_7')
// (21, 4, 'local_g2_7')
// (21, 4, 'lutff_1/in_2')
// (21, 4, 'neigh_op_rgt_7')
// (21, 5, 'neigh_op_bnr_7')
// (22, 3, 'neigh_op_top_7')
// (22, 4, 'lutff_7/out')
// (22, 5, 'neigh_op_bot_7')
// (23, 3, 'neigh_op_tnl_7')
// (23, 4, 'neigh_op_lft_7')
// (23, 5, 'neigh_op_bnl_7')

wire n2916;
// (21, 3, 'sp4_r_v_b_36')
// (21, 4, 'neigh_op_tnr_6')
// (21, 4, 'sp4_r_v_b_25')
// (21, 5, 'neigh_op_rgt_6')
// (21, 5, 'sp4_r_v_b_12')
// (21, 6, 'neigh_op_bnr_6')
// (21, 6, 'sp4_r_v_b_1')
// (22, 2, 'sp4_v_t_36')
// (22, 3, 'sp4_v_b_36')
// (22, 4, 'neigh_op_top_6')
// (22, 4, 'sp4_v_b_25')
// (22, 5, 'lutff_6/out')
// (22, 5, 'sp4_v_b_12')
// (22, 6, 'local_g1_6')
// (22, 6, 'lutff_5/in_0')
// (22, 6, 'neigh_op_bot_6')
// (22, 6, 'sp4_h_r_1')
// (22, 6, 'sp4_v_b_1')
// (23, 4, 'neigh_op_tnl_6')
// (23, 5, 'neigh_op_lft_6')
// (23, 6, 'local_g0_4')
// (23, 6, 'lutff_global/s_r')
// (23, 6, 'neigh_op_bnl_6')
// (23, 6, 'sp4_h_r_12')
// (24, 6, 'sp4_h_r_25')
// (25, 6, 'sp4_h_r_36')

wire n2917;
// (21, 4, 'lutff_0/cout')
// (21, 4, 'lutff_1/in_3')

wire n2918;
// (21, 4, 'lutff_1/cout')
// (21, 4, 'lutff_2/in_3')

wire n2919;
// (21, 4, 'lutff_2/cout')
// (21, 4, 'lutff_3/in_3')

wire n2920;
// (21, 4, 'lutff_3/cout')
// (21, 4, 'lutff_4/in_3')

wire n2921;
// (21, 4, 'lutff_4/cout')
// (21, 4, 'lutff_5/in_3')

wire n2922;
// (21, 4, 'lutff_5/cout')
// (21, 4, 'lutff_6/in_3')

wire n2923;
// (21, 4, 'lutff_6/cout')
// (21, 4, 'lutff_7/in_3')

wire n2924;
// (21, 4, 'lutff_7/cout')
// (21, 5, 'carry_in')
// (21, 5, 'carry_in_mux')
// (21, 5, 'lutff_0/in_3')

wire n2925;
// (21, 4, 'neigh_op_tnr_0')
// (21, 5, 'neigh_op_rgt_0')
// (21, 6, 'neigh_op_bnr_0')
// (22, 4, 'neigh_op_top_0')
// (22, 5, 'local_g2_0')
// (22, 5, 'lutff_0/out')
// (22, 5, 'lutff_7/in_3')
// (22, 6, 'neigh_op_bot_0')
// (23, 4, 'neigh_op_tnl_0')
// (23, 5, 'neigh_op_lft_0')
// (23, 6, 'neigh_op_bnl_0')

wire n2926;
// (21, 4, 'neigh_op_tnr_1')
// (21, 5, 'local_g2_1')
// (21, 5, 'lutff_2/in_1')
// (21, 5, 'neigh_op_rgt_1')
// (21, 6, 'neigh_op_bnr_1')
// (22, 4, 'neigh_op_top_1')
// (22, 5, 'lutff_1/out')
// (22, 6, 'neigh_op_bot_1')
// (23, 4, 'neigh_op_tnl_1')
// (23, 5, 'neigh_op_lft_1')
// (23, 6, 'neigh_op_bnl_1')

wire n2927;
// (21, 4, 'neigh_op_tnr_2')
// (21, 5, 'neigh_op_rgt_2')
// (21, 6, 'neigh_op_bnr_2')
// (22, 4, 'neigh_op_top_2')
// (22, 5, 'local_g2_2')
// (22, 5, 'lutff_2/out')
// (22, 5, 'lutff_6/in_0')
// (22, 5, 'sp4_r_v_b_37')
// (22, 6, 'neigh_op_bot_2')
// (22, 6, 'sp4_r_v_b_24')
// (22, 7, 'sp4_r_v_b_13')
// (22, 8, 'sp4_r_v_b_0')
// (23, 4, 'neigh_op_tnl_2')
// (23, 4, 'sp4_v_t_37')
// (23, 5, 'local_g3_5')
// (23, 5, 'lutff_global/s_r')
// (23, 5, 'neigh_op_lft_2')
// (23, 5, 'sp4_v_b_37')
// (23, 6, 'neigh_op_bnl_2')
// (23, 6, 'sp4_v_b_24')
// (23, 7, 'sp4_v_b_13')
// (23, 8, 'sp4_v_b_0')

wire n2928;
// (21, 4, 'neigh_op_tnr_3')
// (21, 5, 'neigh_op_rgt_3')
// (21, 6, 'neigh_op_bnr_3')
// (22, 4, 'neigh_op_top_3')
// (22, 5, 'local_g3_3')
// (22, 5, 'lutff_0/in_2')
// (22, 5, 'lutff_3/out')
// (22, 6, 'neigh_op_bot_3')
// (23, 4, 'neigh_op_tnl_3')
// (23, 5, 'neigh_op_lft_3')
// (23, 6, 'neigh_op_bnl_3')

wire n2929;
// (21, 4, 'neigh_op_tnr_4')
// (21, 5, 'local_g2_4')
// (21, 5, 'lutff_5/in_1')
// (21, 5, 'neigh_op_rgt_4')
// (21, 6, 'neigh_op_bnr_4')
// (22, 4, 'neigh_op_top_4')
// (22, 5, 'lutff_4/out')
// (22, 6, 'neigh_op_bot_4')
// (23, 4, 'neigh_op_tnl_4')
// (23, 5, 'neigh_op_lft_4')
// (23, 6, 'neigh_op_bnl_4')

wire n2930;
// (21, 5, 'lutff_0/cout')
// (21, 5, 'lutff_1/in_3')

wire n2931;
// (21, 5, 'lutff_1/cout')
// (21, 5, 'lutff_2/in_3')

wire n2932;
// (21, 5, 'lutff_2/cout')
// (21, 5, 'lutff_3/in_3')

wire n2933;
// (21, 5, 'lutff_3/cout')
// (21, 5, 'lutff_4/in_3')

wire n2934;
// (21, 5, 'lutff_4/cout')
// (21, 5, 'lutff_5/in_3')

wire n2935;
// (21, 5, 'lutff_5/cout')
// (21, 5, 'lutff_6/in_3')

wire n2936;
// (21, 5, 'sp4_r_v_b_47')
// (21, 6, 'sp4_r_v_b_34')
// (21, 7, 'neigh_op_tnr_5')
// (21, 7, 'sp4_r_v_b_23')
// (21, 8, 'neigh_op_rgt_5')
// (21, 8, 'sp4_r_v_b_10')
// (21, 9, 'neigh_op_bnr_5')
// (22, 4, 'sp4_v_t_47')
// (22, 5, 'sp4_r_v_b_46')
// (22, 5, 'sp4_v_b_47')
// (22, 6, 'local_g2_2')
// (22, 6, 'lutff_5/in_1')
// (22, 6, 'sp4_r_v_b_35')
// (22, 6, 'sp4_v_b_34')
// (22, 7, 'local_g1_5')
// (22, 7, 'lutff_5/in_1')
// (22, 7, 'neigh_op_top_5')
// (22, 7, 'sp4_r_v_b_22')
// (22, 7, 'sp4_v_b_23')
// (22, 8, 'lutff_5/out')
// (22, 8, 'sp4_r_v_b_11')
// (22, 8, 'sp4_v_b_10')
// (22, 9, 'neigh_op_bot_5')
// (23, 4, 'sp4_v_t_46')
// (23, 5, 'sp4_v_b_46')
// (23, 6, 'local_g3_3')
// (23, 6, 'lutff_2/in_0')
// (23, 6, 'sp4_v_b_35')
// (23, 7, 'neigh_op_tnl_5')
// (23, 7, 'sp4_v_b_22')
// (23, 8, 'neigh_op_lft_5')
// (23, 8, 'sp4_v_b_11')
// (23, 9, 'neigh_op_bnl_5')

wire n2937;
// (21, 6, 'neigh_op_tnr_4')
// (21, 7, 'neigh_op_rgt_4')
// (21, 8, 'neigh_op_bnr_4')
// (22, 6, 'neigh_op_top_4')
// (22, 7, 'lutff_4/out')
// (22, 8, 'local_g0_4')
// (22, 8, 'lutff_5/in_3')
// (22, 8, 'lutff_7/in_3')
// (22, 8, 'neigh_op_bot_4')
// (23, 6, 'neigh_op_tnl_4')
// (23, 7, 'neigh_op_lft_4')
// (23, 8, 'neigh_op_bnl_4')

wire n2938;
// (21, 6, 'neigh_op_tnr_5')
// (21, 7, 'neigh_op_rgt_5')
// (21, 8, 'neigh_op_bnr_5')
// (22, 6, 'neigh_op_top_5')
// (22, 7, 'local_g3_5')
// (22, 7, 'lutff_1/in_3')
// (22, 7, 'lutff_5/out')
// (22, 8, 'neigh_op_bot_5')
// (23, 6, 'neigh_op_tnl_5')
// (23, 7, 'neigh_op_lft_5')
// (23, 8, 'neigh_op_bnl_5')

wire n2939;
// (21, 6, 'neigh_op_tnr_7')
// (21, 7, 'neigh_op_rgt_7')
// (21, 8, 'neigh_op_bnr_7')
// (22, 6, 'neigh_op_top_7')
// (22, 7, 'local_g0_7')
// (22, 7, 'lutff_4/in_1')
// (22, 7, 'lutff_7/out')
// (22, 8, 'neigh_op_bot_7')
// (23, 6, 'neigh_op_tnl_7')
// (23, 7, 'neigh_op_lft_7')
// (23, 8, 'neigh_op_bnl_7')

wire n2940;
// (21, 7, 'local_g3_4')
// (21, 7, 'lutff_1/in_0')
// (21, 7, 'neigh_op_tnr_4')
// (21, 8, 'local_g2_4')
// (21, 8, 'lutff_4/in_2')
// (21, 8, 'lutff_6/in_2')
// (21, 8, 'lutff_7/in_3')
// (21, 8, 'neigh_op_rgt_4')
// (21, 9, 'neigh_op_bnr_4')
// (22, 7, 'local_g0_4')
// (22, 7, 'lutff_1/in_1')
// (22, 7, 'lutff_2/in_2')
// (22, 7, 'lutff_3/in_3')
// (22, 7, 'lutff_6/in_0')
// (22, 7, 'neigh_op_top_4')
// (22, 8, 'lutff_4/out')
// (22, 9, 'neigh_op_bot_4')
// (23, 7, 'neigh_op_tnl_4')
// (23, 8, 'neigh_op_lft_4')
// (23, 9, 'neigh_op_bnl_4')

wire n2941;
// (21, 7, 'lutff_1/cout')
// (21, 7, 'lutff_2/in_3')

wire n2942;
// (21, 7, 'lutff_3/cout')
// (21, 7, 'lutff_4/in_3')

wire n2943;
// (21, 7, 'lutff_5/cout')
// (21, 7, 'lutff_6/in_3')

wire n2944;
// (21, 7, 'lutff_7/cout')
// (21, 8, 'carry_in')
// (21, 8, 'carry_in_mux')
// (21, 8, 'lutff_0/in_3')

wire n2945;
// (21, 7, 'neigh_op_tnr_1')
// (21, 8, 'neigh_op_rgt_1')
// (21, 9, 'neigh_op_bnr_1')
// (22, 7, 'neigh_op_top_1')
// (22, 8, 'lutff_1/out')
// (22, 9, 'neigh_op_bot_1')
// (23, 7, 'neigh_op_tnl_1')
// (23, 8, 'local_g1_1')
// (23, 8, 'lutff_2/in_0')
// (23, 8, 'neigh_op_lft_1')
// (23, 9, 'neigh_op_bnl_1')

reg n2946 = 0;
// (21, 7, 'neigh_op_tnr_3')
// (21, 8, 'neigh_op_rgt_3')
// (21, 9, 'neigh_op_bnr_3')
// (22, 7, 'neigh_op_top_3')
// (22, 8, 'local_g2_3')
// (22, 8, 'lutff_1/in_0')
// (22, 8, 'lutff_3/out')
// (22, 8, 'lutff_6/in_3')
// (22, 9, 'neigh_op_bot_3')
// (23, 7, 'neigh_op_tnl_3')
// (23, 8, 'neigh_op_lft_3')
// (23, 9, 'neigh_op_bnl_3')

wire n2947;
// (21, 7, 'neigh_op_tnr_7')
// (21, 8, 'neigh_op_rgt_7')
// (21, 9, 'neigh_op_bnr_7')
// (22, 7, 'neigh_op_top_7')
// (22, 8, 'local_g2_7')
// (22, 8, 'lutff_3/in_2')
// (22, 8, 'lutff_4/in_1')
// (22, 8, 'lutff_7/out')
// (22, 9, 'neigh_op_bot_7')
// (23, 7, 'neigh_op_tnl_7')
// (23, 8, 'local_g0_7')
// (23, 8, 'lutff_2/in_1')
// (23, 8, 'neigh_op_lft_7')
// (23, 9, 'neigh_op_bnl_7')

wire n2948;
// (21, 8, 'lutff_1/cout')
// (21, 8, 'lutff_2/in_3')

wire n2949;
// (21, 8, 'lutff_3/cout')
// (21, 8, 'lutff_4/in_3')

reg n2950 = 0;
// (21, 8, 'neigh_op_tnr_3')
// (21, 9, 'neigh_op_rgt_3')
// (21, 9, 'sp4_r_v_b_38')
// (21, 10, 'neigh_op_bnr_3')
// (21, 10, 'sp4_r_v_b_27')
// (21, 11, 'sp4_r_v_b_14')
// (21, 12, 'sp4_r_v_b_3')
// (22, 8, 'neigh_op_top_3')
// (22, 8, 'sp4_v_t_38')
// (22, 9, 'lutff_3/out')
// (22, 9, 'sp4_v_b_38')
// (22, 10, 'local_g0_3')
// (22, 10, 'local_g1_3')
// (22, 10, 'lutff_3/in_0')
// (22, 10, 'lutff_5/in_3')
// (22, 10, 'neigh_op_bot_3')
// (22, 10, 'sp4_v_b_27')
// (22, 11, 'local_g1_6')
// (22, 11, 'lutff_3/in_0')
// (22, 11, 'lutff_4/in_1')
// (22, 11, 'sp4_v_b_14')
// (22, 12, 'sp4_v_b_3')
// (23, 8, 'neigh_op_tnl_3')
// (23, 9, 'neigh_op_lft_3')
// (23, 10, 'neigh_op_bnl_3')

reg n2951 = 0;
// (21, 8, 'neigh_op_tnr_4')
// (21, 9, 'neigh_op_rgt_4')
// (21, 10, 'neigh_op_bnr_4')
// (22, 8, 'neigh_op_top_4')
// (22, 9, 'lutff_4/out')
// (22, 10, 'local_g1_4')
// (22, 10, 'lutff_3/in_2')
// (22, 10, 'lutff_4/in_1')
// (22, 10, 'lutff_5/in_2')
// (22, 10, 'neigh_op_bot_4')
// (23, 8, 'neigh_op_tnl_4')
// (23, 9, 'neigh_op_lft_4')
// (23, 10, 'neigh_op_bnl_4')

reg n2952 = 0;
// (21, 8, 'neigh_op_tnr_6')
// (21, 9, 'neigh_op_rgt_6')
// (21, 10, 'neigh_op_bnr_6')
// (22, 8, 'neigh_op_top_6')
// (22, 8, 'sp4_r_v_b_40')
// (22, 9, 'lutff_6/out')
// (22, 9, 'sp4_r_v_b_29')
// (22, 10, 'local_g0_6')
// (22, 10, 'lutff_3/in_3')
// (22, 10, 'lutff_5/in_1')
// (22, 10, 'neigh_op_bot_6')
// (22, 10, 'sp4_r_v_b_16')
// (22, 11, 'local_g1_5')
// (22, 11, 'lutff_3/in_1')
// (22, 11, 'lutff_4/in_0')
// (22, 11, 'sp4_r_v_b_5')
// (23, 7, 'sp4_v_t_40')
// (23, 8, 'neigh_op_tnl_6')
// (23, 8, 'sp4_v_b_40')
// (23, 9, 'neigh_op_lft_6')
// (23, 9, 'sp4_v_b_29')
// (23, 10, 'neigh_op_bnl_6')
// (23, 10, 'sp4_v_b_16')
// (23, 11, 'sp4_v_b_5')

reg n2953 = 0;
// (21, 8, 'neigh_op_tnr_7')
// (21, 9, 'neigh_op_rgt_7')
// (21, 10, 'neigh_op_bnr_7')
// (22, 8, 'neigh_op_top_7')
// (22, 9, 'lutff_7/out')
// (22, 10, 'local_g0_7')
// (22, 10, 'lutff_4/in_3')
// (22, 10, 'lutff_5/in_0')
// (22, 10, 'neigh_op_bot_7')
// (23, 8, 'neigh_op_tnl_7')
// (23, 9, 'neigh_op_lft_7')
// (23, 10, 'neigh_op_bnl_7')

wire n2954;
// (21, 9, 'neigh_op_tnr_4')
// (21, 10, 'neigh_op_rgt_4')
// (21, 11, 'neigh_op_bnr_4')
// (22, 9, 'neigh_op_top_4')
// (22, 10, 'lutff_4/out')
// (22, 11, 'local_g0_4')
// (22, 11, 'lutff_3/in_3')
// (22, 11, 'lutff_4/in_2')
// (22, 11, 'neigh_op_bot_4')
// (23, 9, 'neigh_op_tnl_4')
// (23, 10, 'neigh_op_lft_4')
// (23, 11, 'neigh_op_bnl_4')

wire n2955;
// (21, 10, 'neigh_op_tnr_2')
// (21, 11, 'neigh_op_rgt_2')
// (21, 12, 'neigh_op_bnr_2')
// (22, 10, 'neigh_op_top_2')
// (22, 11, 'local_g0_2')
// (22, 11, 'lutff_2/out')
// (22, 11, 'lutff_global/cen')
// (22, 12, 'neigh_op_bot_2')
// (23, 10, 'neigh_op_tnl_2')
// (23, 11, 'neigh_op_lft_2')
// (23, 12, 'neigh_op_bnl_2')

reg n2956 = 0;
// (21, 11, 'neigh_op_tnr_0')
// (21, 12, 'local_g2_0')
// (21, 12, 'lutff_0/in_2')
// (21, 12, 'neigh_op_rgt_0')
// (21, 13, 'neigh_op_bnr_0')
// (22, 11, 'neigh_op_top_0')
// (22, 12, 'lutff_0/out')
// (22, 13, 'neigh_op_bot_0')
// (23, 11, 'neigh_op_tnl_0')
// (23, 12, 'neigh_op_lft_0')
// (23, 13, 'neigh_op_bnl_0')

wire n2957;
// (21, 11, 'neigh_op_tnr_2')
// (21, 12, 'neigh_op_rgt_2')
// (21, 13, 'neigh_op_bnr_2')
// (22, 10, 'sp4_r_v_b_45')
// (22, 11, 'neigh_op_top_2')
// (22, 11, 'sp4_r_v_b_32')
// (22, 12, 'lutff_2/out')
// (22, 12, 'sp4_r_v_b_21')
// (22, 13, 'neigh_op_bot_2')
// (22, 13, 'sp4_r_v_b_8')
// (23, 9, 'sp4_v_t_45')
// (23, 10, 'sp4_v_b_45')
// (23, 11, 'neigh_op_tnl_2')
// (23, 11, 'sp4_v_b_32')
// (23, 12, 'local_g1_5')
// (23, 12, 'lutff_global/s_r')
// (23, 12, 'neigh_op_lft_2')
// (23, 12, 'sp4_v_b_21')
// (23, 13, 'neigh_op_bnl_2')
// (23, 13, 'sp4_v_b_8')

reg n2958 = 0;
// (21, 12, 'neigh_op_tnr_0')
// (21, 13, 'neigh_op_rgt_0')
// (21, 14, 'local_g0_0')
// (21, 14, 'lutff_3/in_1')
// (21, 14, 'neigh_op_bnr_0')
// (22, 12, 'neigh_op_top_0')
// (22, 13, 'lutff_0/out')
// (22, 14, 'neigh_op_bot_0')
// (23, 12, 'neigh_op_tnl_0')
// (23, 13, 'neigh_op_lft_0')
// (23, 14, 'neigh_op_bnl_0')

reg n2959 = 0;
// (21, 12, 'neigh_op_tnr_2')
// (21, 13, 'neigh_op_rgt_2')
// (21, 14, 'neigh_op_bnr_2')
// (22, 12, 'neigh_op_top_2')
// (22, 13, 'lutff_2/out')
// (22, 14, 'neigh_op_bot_2')
// (23, 12, 'neigh_op_tnl_2')
// (23, 13, 'local_g1_2')
// (23, 13, 'lutff_0/in_1')
// (23, 13, 'neigh_op_lft_2')
// (23, 14, 'neigh_op_bnl_2')

reg n2960 = 0;
// (21, 12, 'neigh_op_tnr_3')
// (21, 13, 'neigh_op_rgt_3')
// (21, 14, 'neigh_op_bnr_3')
// (22, 12, 'neigh_op_top_3')
// (22, 13, 'lutff_3/out')
// (22, 14, 'neigh_op_bot_3')
// (23, 12, 'neigh_op_tnl_3')
// (23, 13, 'local_g1_3')
// (23, 13, 'lutff_2/in_2')
// (23, 13, 'neigh_op_lft_3')
// (23, 14, 'neigh_op_bnl_3')

wire n2961;
// (21, 12, 'neigh_op_tnr_7')
// (21, 13, 'neigh_op_rgt_7')
// (21, 14, 'local_g0_7')
// (21, 14, 'lutff_6/in_3')
// (21, 14, 'neigh_op_bnr_7')
// (22, 12, 'neigh_op_top_7')
// (22, 13, 'lutff_7/out')
// (22, 14, 'neigh_op_bot_7')
// (23, 12, 'neigh_op_tnl_7')
// (23, 13, 'neigh_op_lft_7')
// (23, 14, 'neigh_op_bnl_7')

reg n2962 = 0;
// (21, 13, 'local_g1_4')
// (21, 13, 'lutff_4/in_1')
// (21, 13, 'sp4_h_r_4')
// (22, 12, 'neigh_op_tnr_6')
// (22, 13, 'neigh_op_rgt_6')
// (22, 13, 'sp4_h_r_17')
// (22, 14, 'neigh_op_bnr_6')
// (23, 12, 'neigh_op_top_6')
// (23, 13, 'lutff_6/out')
// (23, 13, 'sp4_h_r_28')
// (23, 14, 'neigh_op_bot_6')
// (24, 12, 'neigh_op_tnl_6')
// (24, 13, 'neigh_op_lft_6')
// (24, 13, 'sp4_h_r_41')
// (24, 14, 'neigh_op_bnl_6')
// (25, 13, 'sp4_h_l_41')

wire n2963;
// (21, 13, 'lutff_1/cout')
// (21, 13, 'lutff_2/in_3')

wire n2964;
// (21, 13, 'lutff_2/cout')
// (21, 13, 'lutff_3/in_3')

wire n2965;
// (21, 13, 'neigh_op_tnr_1')
// (21, 14, 'neigh_op_rgt_1')
// (21, 15, 'neigh_op_bnr_1')
// (22, 13, 'neigh_op_top_1')
// (22, 14, 'lutff_1/out')
// (22, 15, 'neigh_op_bot_1')
// (23, 13, 'neigh_op_tnl_1')
// (23, 14, 'local_g1_1')
// (23, 14, 'lutff_0/in_2')
// (23, 14, 'neigh_op_lft_1')
// (23, 15, 'neigh_op_bnl_1')

reg n2966 = 0;
// (21, 13, 'neigh_op_tnr_2')
// (21, 14, 'neigh_op_rgt_2')
// (21, 15, 'neigh_op_bnr_2')
// (22, 13, 'neigh_op_top_2')
// (22, 14, 'local_g0_2')
// (22, 14, 'lutff_2/in_2')
// (22, 14, 'lutff_2/out')
// (22, 15, 'local_g0_2')
// (22, 15, 'lutff_5/in_1')
// (22, 15, 'neigh_op_bot_2')
// (23, 13, 'neigh_op_tnl_2')
// (23, 14, 'neigh_op_lft_2')
// (23, 15, 'neigh_op_bnl_2')

wire n2967;
// (21, 13, 'neigh_op_tnr_3')
// (21, 14, 'neigh_op_rgt_3')
// (21, 15, 'neigh_op_bnr_3')
// (22, 13, 'neigh_op_top_3')
// (22, 14, 'lutff_3/out')
// (22, 15, 'neigh_op_bot_3')
// (23, 13, 'neigh_op_tnl_3')
// (23, 14, 'local_g1_3')
// (23, 14, 'lutff_5/in_1')
// (23, 14, 'neigh_op_lft_3')
// (23, 15, 'neigh_op_bnl_3')

wire n2968;
// (21, 13, 'neigh_op_tnr_4')
// (21, 14, 'neigh_op_rgt_4')
// (21, 15, 'neigh_op_bnr_4')
// (22, 13, 'neigh_op_top_4')
// (22, 14, 'lutff_4/out')
// (22, 15, 'neigh_op_bot_4')
// (23, 13, 'neigh_op_tnl_4')
// (23, 14, 'local_g0_4')
// (23, 14, 'lutff_2/in_0')
// (23, 14, 'neigh_op_lft_4')
// (23, 15, 'neigh_op_bnl_4')

reg n2969 = 0;
// (21, 13, 'neigh_op_tnr_6')
// (21, 14, 'neigh_op_rgt_6')
// (21, 15, 'neigh_op_bnr_6')
// (22, 13, 'neigh_op_top_6')
// (22, 14, 'local_g3_6')
// (22, 14, 'lutff_6/in_1')
// (22, 14, 'lutff_6/out')
// (22, 15, 'local_g0_6')
// (22, 15, 'lutff_7/in_1')
// (22, 15, 'neigh_op_bot_6')
// (23, 13, 'neigh_op_tnl_6')
// (23, 14, 'neigh_op_lft_6')
// (23, 15, 'neigh_op_bnl_6')

wire n2970;
// (21, 13, 'neigh_op_tnr_7')
// (21, 14, 'neigh_op_rgt_7')
// (21, 15, 'neigh_op_bnr_7')
// (22, 13, 'neigh_op_top_7')
// (22, 14, 'lutff_7/out')
// (22, 15, 'neigh_op_bot_7')
// (23, 13, 'neigh_op_tnl_7')
// (23, 14, 'local_g0_7')
// (23, 14, 'lutff_6/in_3')
// (23, 14, 'neigh_op_lft_7')
// (23, 15, 'neigh_op_bnl_7')

wire n2971;
// (21, 13, 'sp4_r_v_b_45')
// (21, 14, 'sp4_r_v_b_32')
// (21, 15, 'neigh_op_tnr_4')
// (21, 15, 'sp4_r_v_b_21')
// (21, 16, 'neigh_op_rgt_4')
// (21, 16, 'sp4_r_v_b_8')
// (21, 17, 'neigh_op_bnr_4')
// (22, 12, 'sp4_v_t_45')
// (22, 13, 'sp4_v_b_45')
// (22, 14, 'sp4_v_b_32')
// (22, 15, 'neigh_op_top_4')
// (22, 15, 'sp4_v_b_21')
// (22, 16, 'local_g0_2')
// (22, 16, 'lutff_4/out')
// (22, 16, 'lutff_global/cen')
// (22, 16, 'sp4_h_r_2')
// (22, 16, 'sp4_v_b_8')
// (22, 17, 'neigh_op_bot_4')
// (23, 15, 'neigh_op_tnl_4')
// (23, 16, 'neigh_op_lft_4')
// (23, 16, 'sp4_h_r_15')
// (23, 17, 'neigh_op_bnl_4')
// (24, 16, 'sp4_h_r_26')
// (25, 16, 'sp4_h_r_39')

wire n2972;
// (21, 14, 'neigh_op_tnr_1')
// (21, 15, 'neigh_op_rgt_1')
// (21, 16, 'neigh_op_bnr_1')
// (22, 14, 'neigh_op_top_1')
// (22, 15, 'lutff_1/out')
// (22, 16, 'neigh_op_bot_1')
// (23, 14, 'local_g2_1')
// (23, 14, 'lutff_4/in_3')
// (23, 14, 'neigh_op_tnl_1')
// (23, 15, 'neigh_op_lft_1')
// (23, 16, 'neigh_op_bnl_1')

reg n2973 = 0;
// (21, 14, 'neigh_op_tnr_3')
// (21, 15, 'neigh_op_rgt_3')
// (21, 16, 'neigh_op_bnr_3')
// (22, 14, 'neigh_op_top_3')
// (22, 15, 'local_g1_3')
// (22, 15, 'lutff_3/in_1')
// (22, 15, 'lutff_3/out')
// (22, 15, 'lutff_7/in_3')
// (22, 16, 'neigh_op_bot_3')
// (23, 14, 'neigh_op_tnl_3')
// (23, 15, 'neigh_op_lft_3')
// (23, 16, 'neigh_op_bnl_3')

reg n2974 = 0;
// (21, 14, 'neigh_op_tnr_4')
// (21, 15, 'neigh_op_rgt_4')
// (21, 16, 'neigh_op_bnr_4')
// (22, 14, 'neigh_op_top_4')
// (22, 15, 'local_g3_4')
// (22, 15, 'lutff_4/in_1')
// (22, 15, 'lutff_4/out')
// (22, 15, 'lutff_7/in_0')
// (22, 16, 'neigh_op_bot_4')
// (23, 14, 'neigh_op_tnl_4')
// (23, 15, 'neigh_op_lft_4')
// (23, 16, 'neigh_op_bnl_4')

wire n2975;
// (21, 14, 'neigh_op_tnr_5')
// (21, 15, 'neigh_op_rgt_5')
// (21, 16, 'neigh_op_bnr_5')
// (22, 14, 'neigh_op_top_5')
// (22, 15, 'lutff_5/out')
// (22, 16, 'neigh_op_bot_5')
// (23, 14, 'neigh_op_tnl_5')
// (23, 15, 'local_g0_5')
// (23, 15, 'lutff_2/in_3')
// (23, 15, 'neigh_op_lft_5')
// (23, 16, 'neigh_op_bnl_5')

reg n2976 = 0;
// (21, 14, 'neigh_op_tnr_6')
// (21, 15, 'neigh_op_rgt_6')
// (21, 16, 'neigh_op_bnr_6')
// (22, 14, 'local_g0_6')
// (22, 14, 'lutff_0/in_2')
// (22, 14, 'lutff_1/in_3')
// (22, 14, 'neigh_op_top_6')
// (22, 15, 'local_g2_6')
// (22, 15, 'lutff_5/in_3')
// (22, 15, 'lutff_6/in_0')
// (22, 15, 'lutff_6/out')
// (22, 16, 'neigh_op_bot_6')
// (23, 14, 'neigh_op_tnl_6')
// (23, 15, 'neigh_op_lft_6')
// (23, 16, 'neigh_op_bnl_6')

wire n2977;
// (21, 14, 'neigh_op_tnr_7')
// (21, 15, 'neigh_op_rgt_7')
// (21, 16, 'neigh_op_bnr_7')
// (22, 14, 'neigh_op_top_7')
// (22, 15, 'lutff_7/out')
// (22, 16, 'neigh_op_bot_7')
// (23, 14, 'neigh_op_tnl_7')
// (23, 15, 'local_g0_7')
// (23, 15, 'lutff_2/in_1')
// (23, 15, 'neigh_op_lft_7')
// (23, 16, 'neigh_op_bnl_7')

wire n2978;
// (21, 15, 'neigh_op_tnr_2')
// (21, 16, 'local_g3_2')
// (21, 16, 'lutff_0/in_1')
// (21, 16, 'neigh_op_rgt_2')
// (21, 17, 'neigh_op_bnr_2')
// (22, 15, 'neigh_op_top_2')
// (22, 16, 'lutff_2/out')
// (22, 17, 'neigh_op_bot_2')
// (23, 15, 'neigh_op_tnl_2')
// (23, 16, 'neigh_op_lft_2')
// (23, 17, 'neigh_op_bnl_2')

reg n2979 = 0;
// (21, 15, 'neigh_op_tnr_3')
// (21, 16, 'neigh_op_rgt_3')
// (21, 17, 'local_g0_3')
// (21, 17, 'lutff_5/in_0')
// (21, 17, 'neigh_op_bnr_3')
// (22, 15, 'neigh_op_top_3')
// (22, 16, 'lutff_3/out')
// (22, 17, 'neigh_op_bot_3')
// (23, 15, 'neigh_op_tnl_3')
// (23, 16, 'neigh_op_lft_3')
// (23, 17, 'neigh_op_bnl_3')

wire n2980;
// (21, 15, 'neigh_op_tnr_5')
// (21, 16, 'neigh_op_rgt_5')
// (21, 17, 'neigh_op_bnr_5')
// (22, 15, 'neigh_op_top_5')
// (22, 16, 'lutff_5/out')
// (22, 16, 'sp4_h_r_10')
// (22, 17, 'neigh_op_bot_5')
// (23, 15, 'neigh_op_tnl_5')
// (23, 16, 'neigh_op_lft_5')
// (23, 16, 'sp4_h_r_23')
// (23, 17, 'neigh_op_bnl_5')
// (24, 16, 'local_g2_2')
// (24, 16, 'lutff_global/cen')
// (24, 16, 'sp4_h_r_34')
// (25, 16, 'sp4_h_r_47')

wire n2981;
// (21, 15, 'neigh_op_tnr_6')
// (21, 16, 'neigh_op_rgt_6')
// (21, 16, 'sp4_r_v_b_44')
// (21, 17, 'neigh_op_bnr_6')
// (21, 17, 'sp4_r_v_b_33')
// (21, 18, 'sp4_r_v_b_20')
// (21, 19, 'sp4_r_v_b_9')
// (22, 15, 'neigh_op_top_6')
// (22, 15, 'sp4_h_r_2')
// (22, 15, 'sp4_v_t_44')
// (22, 16, 'lutff_6/out')
// (22, 16, 'sp4_v_b_44')
// (22, 17, 'neigh_op_bot_6')
// (22, 17, 'sp4_v_b_33')
// (22, 18, 'sp4_v_b_20')
// (22, 19, 'sp4_v_b_9')
// (23, 15, 'neigh_op_tnl_6')
// (23, 15, 'sp4_h_r_15')
// (23, 16, 'neigh_op_lft_6')
// (23, 17, 'neigh_op_bnl_6')
// (24, 15, 'local_g2_2')
// (24, 15, 'lutff_global/cen')
// (24, 15, 'sp4_h_r_26')
// (25, 15, 'sp4_h_r_39')

wire n2982;
// (21, 15, 'neigh_op_tnr_7')
// (21, 16, 'neigh_op_rgt_7')
// (21, 17, 'neigh_op_bnr_7')
// (22, 14, 'sp4_r_v_b_39')
// (22, 15, 'neigh_op_top_7')
// (22, 15, 'sp4_r_v_b_26')
// (22, 16, 'lutff_7/out')
// (22, 16, 'sp4_r_v_b_15')
// (22, 17, 'neigh_op_bot_7')
// (22, 17, 'sp4_r_v_b_2')
// (23, 13, 'sp4_v_t_39')
// (23, 14, 'sp4_v_b_39')
// (23, 15, 'local_g2_2')
// (23, 15, 'lutff_global/cen')
// (23, 15, 'neigh_op_tnl_7')
// (23, 15, 'sp4_v_b_26')
// (23, 16, 'neigh_op_lft_7')
// (23, 16, 'sp4_v_b_15')
// (23, 17, 'neigh_op_bnl_7')
// (23, 17, 'sp4_v_b_2')

reg n2983 = 0;
// (21, 16, 'local_g0_6')
// (21, 16, 'lutff_1/in_3')
// (21, 16, 'sp4_h_r_6')
// (22, 16, 'sp4_h_r_19')
// (23, 14, 'neigh_op_tnr_1')
// (23, 15, 'neigh_op_rgt_1')
// (23, 16, 'neigh_op_bnr_1')
// (23, 16, 'sp4_h_r_30')
// (24, 13, 'sp4_r_v_b_43')
// (24, 14, 'neigh_op_top_1')
// (24, 14, 'sp4_r_v_b_30')
// (24, 15, 'lutff_1/out')
// (24, 15, 'sp4_r_v_b_19')
// (24, 16, 'neigh_op_bot_1')
// (24, 16, 'sp4_h_r_43')
// (24, 16, 'sp4_r_v_b_6')
// (25, 12, 'sp4_v_t_43')
// (25, 13, 'sp4_v_b_43')
// (25, 14, 'neigh_op_tnl_1')
// (25, 14, 'sp4_v_b_30')
// (25, 15, 'neigh_op_lft_1')
// (25, 15, 'sp4_v_b_19')
// (25, 16, 'neigh_op_bnl_1')
// (25, 16, 'sp4_h_l_43')
// (25, 16, 'sp4_v_b_6')

reg n2984 = 0;
// (21, 16, 'neigh_op_tnr_2')
// (21, 17, 'local_g3_2')
// (21, 17, 'lutff_4/in_3')
// (21, 17, 'neigh_op_rgt_2')
// (21, 18, 'neigh_op_bnr_2')
// (22, 16, 'neigh_op_top_2')
// (22, 17, 'lutff_2/out')
// (22, 18, 'neigh_op_bot_2')
// (23, 16, 'neigh_op_tnl_2')
// (23, 17, 'neigh_op_lft_2')
// (23, 18, 'neigh_op_bnl_2')

wire n2985;
// (21, 16, 'neigh_op_tnr_4')
// (21, 17, 'neigh_op_rgt_4')
// (21, 18, 'neigh_op_bnr_4')
// (22, 14, 'sp4_r_v_b_44')
// (22, 15, 'sp4_r_v_b_33')
// (22, 16, 'neigh_op_top_4')
// (22, 16, 'sp4_r_v_b_20')
// (22, 17, 'lutff_4/out')
// (22, 17, 'sp4_r_v_b_9')
// (22, 18, 'neigh_op_bot_4')
// (23, 13, 'sp4_v_t_44')
// (23, 14, 'sp4_v_b_44')
// (23, 15, 'sp4_v_b_33')
// (23, 16, 'neigh_op_tnl_4')
// (23, 16, 'sp4_v_b_20')
// (23, 17, 'local_g1_3')
// (23, 17, 'lutff_global/cen')
// (23, 17, 'neigh_op_lft_4')
// (23, 17, 'sp4_h_r_3')
// (23, 17, 'sp4_v_b_9')
// (23, 18, 'neigh_op_bnl_4')
// (24, 17, 'sp4_h_r_14')
// (25, 17, 'sp4_h_r_27')

wire n2986;
// (21, 16, 'sp4_r_v_b_47')
// (21, 17, 'sp4_r_v_b_34')
// (21, 18, 'local_g3_5')
// (21, 18, 'lutff_6/in_2')
// (21, 18, 'neigh_op_tnr_5')
// (21, 18, 'sp4_r_v_b_23')
// (21, 19, 'neigh_op_rgt_5')
// (21, 19, 'sp4_r_v_b_10')
// (21, 20, 'neigh_op_bnr_5')
// (21, 20, 'sp4_r_v_b_41')
// (21, 21, 'sp4_r_v_b_28')
// (21, 22, 'sp4_r_v_b_17')
// (21, 23, 'local_g1_4')
// (21, 23, 'lutff_4/in_1')
// (21, 23, 'sp4_r_v_b_4')
// (22, 15, 'sp4_v_t_47')
// (22, 16, 'local_g2_7')
// (22, 16, 'lutff_6/in_1')
// (22, 16, 'sp4_v_b_47')
// (22, 17, 'local_g3_2')
// (22, 17, 'lutff_3/in_2')
// (22, 17, 'lutff_4/in_1')
// (22, 17, 'sp4_v_b_34')
// (22, 18, 'neigh_op_top_5')
// (22, 18, 'sp4_v_b_23')
// (22, 19, 'local_g0_5')
// (22, 19, 'lutff_0/in_3')
// (22, 19, 'lutff_5/out')
// (22, 19, 'sp4_h_r_10')
// (22, 19, 'sp4_v_b_10')
// (22, 19, 'sp4_v_t_41')
// (22, 20, 'neigh_op_bot_5')
// (22, 20, 'sp4_v_b_41')
// (22, 21, 'sp4_v_b_28')
// (22, 22, 'sp4_v_b_17')
// (22, 23, 'local_g1_4')
// (22, 23, 'lutff_1/in_2')
// (22, 23, 'sp4_v_b_4')
// (23, 18, 'neigh_op_tnl_5')
// (23, 19, 'neigh_op_lft_5')
// (23, 19, 'sp4_h_r_23')
// (23, 20, 'neigh_op_bnl_5')
// (24, 19, 'sp4_h_r_34')
// (25, 19, 'sp4_h_r_47')

wire n2987;
// (21, 17, 'neigh_op_tnr_1')
// (21, 18, 'neigh_op_rgt_1')
// (21, 19, 'neigh_op_bnr_1')
// (22, 15, 'sp4_r_v_b_38')
// (22, 16, 'sp4_r_v_b_27')
// (22, 17, 'neigh_op_top_1')
// (22, 17, 'sp4_r_v_b_14')
// (22, 18, 'lutff_1/out')
// (22, 18, 'sp4_r_v_b_3')
// (22, 19, 'neigh_op_bot_1')
// (23, 14, 'sp4_v_t_38')
// (23, 15, 'sp4_v_b_38')
// (23, 16, 'sp4_v_b_27')
// (23, 17, 'neigh_op_tnl_1')
// (23, 17, 'sp4_v_b_14')
// (23, 18, 'local_g1_3')
// (23, 18, 'lutff_global/cen')
// (23, 18, 'neigh_op_lft_1')
// (23, 18, 'sp4_v_b_3')
// (23, 19, 'neigh_op_bnl_1')

wire n2988;
// (21, 17, 'neigh_op_tnr_2')
// (21, 18, 'local_g2_2')
// (21, 18, 'lutff_3/in_1')
// (21, 18, 'neigh_op_rgt_2')
// (21, 19, 'neigh_op_bnr_2')
// (22, 17, 'neigh_op_top_2')
// (22, 18, 'lutff_2/out')
// (22, 19, 'neigh_op_bot_2')
// (23, 17, 'neigh_op_tnl_2')
// (23, 18, 'neigh_op_lft_2')
// (23, 19, 'neigh_op_bnl_2')

wire n2989;
// (21, 17, 'neigh_op_tnr_3')
// (21, 18, 'neigh_op_rgt_3')
// (21, 19, 'neigh_op_bnr_3')
// (22, 17, 'neigh_op_top_3')
// (22, 18, 'local_g3_3')
// (22, 18, 'lutff_3/out')
// (22, 18, 'lutff_global/cen')
// (22, 19, 'neigh_op_bot_3')
// (23, 17, 'neigh_op_tnl_3')
// (23, 18, 'neigh_op_lft_3')
// (23, 19, 'neigh_op_bnl_3')

reg n2990 = 0;
// (21, 17, 'neigh_op_tnr_6')
// (21, 18, 'neigh_op_rgt_6')
// (21, 19, 'neigh_op_bnr_6')
// (22, 17, 'neigh_op_top_6')
// (22, 18, 'local_g2_6')
// (22, 18, 'lutff_6/out')
// (22, 18, 'lutff_7/in_3')
// (22, 19, 'neigh_op_bot_6')
// (23, 17, 'neigh_op_tnl_6')
// (23, 18, 'neigh_op_lft_6')
// (23, 19, 'neigh_op_bnl_6')

wire n2991;
// (21, 17, 'neigh_op_tnr_7')
// (21, 18, 'local_g2_7')
// (21, 18, 'lutff_3/in_2')
// (21, 18, 'neigh_op_rgt_7')
// (21, 19, 'neigh_op_bnr_7')
// (22, 17, 'neigh_op_top_7')
// (22, 18, 'lutff_7/out')
// (22, 19, 'neigh_op_bot_7')
// (23, 17, 'neigh_op_tnl_7')
// (23, 18, 'neigh_op_lft_7')
// (23, 19, 'neigh_op_bnl_7')

wire n2992;
// (21, 17, 'sp4_r_v_b_38')
// (21, 18, 'neigh_op_tnr_7')
// (21, 18, 'sp4_r_v_b_27')
// (21, 19, 'neigh_op_rgt_7')
// (21, 19, 'sp4_r_v_b_14')
// (21, 20, 'neigh_op_bnr_7')
// (21, 20, 'sp4_r_v_b_3')
// (22, 16, 'local_g0_0')
// (22, 16, 'lutff_4/in_0')
// (22, 16, 'lutff_5/in_1')
// (22, 16, 'lutff_7/in_1')
// (22, 16, 'sp4_h_r_8')
// (22, 16, 'sp4_v_t_38')
// (22, 17, 'sp4_v_b_38')
// (22, 18, 'local_g0_7')
// (22, 18, 'lutff_1/in_0')
// (22, 18, 'neigh_op_top_7')
// (22, 18, 'sp4_v_b_27')
// (22, 19, 'local_g2_7')
// (22, 19, 'lutff_4/in_1')
// (22, 19, 'lutff_6/in_1')
// (22, 19, 'lutff_7/out')
// (22, 19, 'sp4_v_b_14')
// (22, 20, 'local_g1_7')
// (22, 20, 'lutff_6/in_2')
// (22, 20, 'lutff_7/in_1')
// (22, 20, 'neigh_op_bot_7')
// (22, 20, 'sp4_v_b_3')
// (23, 16, 'sp4_h_r_21')
// (23, 18, 'neigh_op_tnl_7')
// (23, 19, 'neigh_op_lft_7')
// (23, 20, 'neigh_op_bnl_7')
// (24, 16, 'sp4_h_r_32')
// (25, 16, 'sp4_h_r_45')

wire n2993;
// (21, 18, 'neigh_op_tnr_4')
// (21, 19, 'neigh_op_rgt_4')
// (21, 20, 'neigh_op_bnr_4')
// (22, 16, 'sp4_r_v_b_44')
// (22, 17, 'sp4_r_v_b_33')
// (22, 18, 'neigh_op_top_4')
// (22, 18, 'sp4_r_v_b_20')
// (22, 19, 'lutff_4/out')
// (22, 19, 'sp4_r_v_b_9')
// (22, 20, 'neigh_op_bot_4')
// (23, 15, 'sp4_v_t_44')
// (23, 16, 'sp4_v_b_44')
// (23, 17, 'sp4_v_b_33')
// (23, 18, 'neigh_op_tnl_4')
// (23, 18, 'sp4_v_b_20')
// (23, 19, 'local_g1_3')
// (23, 19, 'lutff_global/cen')
// (23, 19, 'neigh_op_lft_4')
// (23, 19, 'sp4_h_r_3')
// (23, 19, 'sp4_v_b_9')
// (23, 20, 'neigh_op_bnl_4')
// (24, 19, 'sp4_h_r_14')
// (25, 19, 'sp4_h_r_27')

reg n2994 = 0;
// (21, 18, 'sp4_h_r_3')
// (22, 18, 'local_g1_6')
// (22, 18, 'lutff_2/in_1')
// (22, 18, 'sp4_h_r_14')
// (23, 17, 'neigh_op_tnr_3')
// (23, 18, 'neigh_op_rgt_3')
// (23, 18, 'sp4_h_r_27')
// (23, 19, 'neigh_op_bnr_3')
// (24, 17, 'neigh_op_top_3')
// (24, 18, 'lutff_3/out')
// (24, 18, 'sp4_h_r_38')
// (24, 19, 'neigh_op_bot_3')
// (25, 17, 'neigh_op_tnl_3')
// (25, 18, 'neigh_op_lft_3')
// (25, 18, 'sp4_h_l_38')
// (25, 19, 'neigh_op_bnl_3')

wire n2995;
// (21, 18, 'sp4_r_v_b_38')
// (21, 19, 'neigh_op_tnr_7')
// (21, 19, 'sp4_r_v_b_27')
// (21, 20, 'neigh_op_rgt_7')
// (21, 20, 'sp4_r_v_b_14')
// (21, 21, 'neigh_op_bnr_7')
// (21, 21, 'sp4_r_v_b_3')
// (22, 17, 'sp4_v_t_38')
// (22, 18, 'sp4_v_b_38')
// (22, 19, 'neigh_op_top_7')
// (22, 19, 'sp4_v_b_27')
// (22, 20, 'lutff_7/out')
// (22, 20, 'sp4_v_b_14')
// (22, 21, 'neigh_op_bot_7')
// (22, 21, 'sp4_h_r_3')
// (22, 21, 'sp4_v_b_3')
// (23, 19, 'neigh_op_tnl_7')
// (23, 20, 'neigh_op_lft_7')
// (23, 21, 'neigh_op_bnl_7')
// (23, 21, 'sp4_h_r_14')
// (24, 21, 'local_g3_3')
// (24, 21, 'lutff_global/cen')
// (24, 21, 'sp4_h_r_27')
// (25, 21, 'sp4_h_r_38')

reg n2996 = 0;
// (21, 19, 'neigh_op_tnr_1')
// (21, 20, 'local_g3_1')
// (21, 20, 'lutff_4/in_0')
// (21, 20, 'neigh_op_rgt_1')
// (21, 21, 'neigh_op_bnr_1')
// (22, 19, 'neigh_op_top_1')
// (22, 20, 'lutff_1/out')
// (22, 21, 'neigh_op_bot_1')
// (23, 19, 'neigh_op_tnl_1')
// (23, 20, 'neigh_op_lft_1')
// (23, 21, 'neigh_op_bnl_1')

wire n2997;
// (21, 19, 'neigh_op_tnr_2')
// (21, 20, 'neigh_op_rgt_2')
// (21, 21, 'neigh_op_bnr_2')
// (22, 19, 'neigh_op_top_2')
// (22, 20, 'lutff_2/out')
// (22, 21, 'neigh_op_bot_2')
// (23, 19, 'neigh_op_tnl_2')
// (23, 20, 'local_g0_2')
// (23, 20, 'lutff_global/cen')
// (23, 20, 'neigh_op_lft_2')
// (23, 21, 'neigh_op_bnl_2')

wire n2998;
// (21, 19, 'neigh_op_tnr_3')
// (21, 20, 'neigh_op_rgt_3')
// (21, 21, 'neigh_op_bnr_3')
// (22, 19, 'neigh_op_top_3')
// (22, 20, 'local_g1_3')
// (22, 20, 'lutff_3/out')
// (22, 20, 'lutff_global/cen')
// (22, 21, 'neigh_op_bot_3')
// (23, 19, 'neigh_op_tnl_3')
// (23, 20, 'neigh_op_lft_3')
// (23, 21, 'neigh_op_bnl_3')

reg n2999 = 0;
// (21, 20, 'local_g1_1')
// (21, 20, 'lutff_2/in_2')
// (21, 20, 'sp4_h_r_1')
// (22, 20, 'sp4_h_r_12')
// (23, 19, 'neigh_op_tnr_2')
// (23, 20, 'neigh_op_rgt_2')
// (23, 20, 'sp4_h_r_25')
// (23, 21, 'neigh_op_bnr_2')
// (24, 19, 'neigh_op_top_2')
// (24, 20, 'lutff_2/out')
// (24, 20, 'sp4_h_r_36')
// (24, 21, 'neigh_op_bot_2')
// (25, 19, 'neigh_op_tnl_2')
// (25, 20, 'neigh_op_lft_2')
// (25, 20, 'sp4_h_l_36')
// (25, 21, 'neigh_op_bnl_2')

reg n3000 = 0;
// (21, 20, 'neigh_op_tnr_3')
// (21, 21, 'local_g2_3')
// (21, 21, 'lutff_7/in_2')
// (21, 21, 'neigh_op_rgt_3')
// (21, 22, 'neigh_op_bnr_3')
// (22, 20, 'neigh_op_top_3')
// (22, 21, 'lutff_3/out')
// (22, 22, 'neigh_op_bot_3')
// (23, 20, 'neigh_op_tnl_3')
// (23, 21, 'neigh_op_lft_3')
// (23, 22, 'neigh_op_bnl_3')

wire n3001;
// (21, 20, 'neigh_op_tnr_4')
// (21, 21, 'local_g3_4')
// (21, 21, 'lutff_5/in_0')
// (21, 21, 'neigh_op_rgt_4')
// (21, 22, 'neigh_op_bnr_4')
// (22, 20, 'neigh_op_top_4')
// (22, 21, 'lutff_4/out')
// (22, 22, 'neigh_op_bot_4')
// (23, 20, 'neigh_op_tnl_4')
// (23, 21, 'neigh_op_lft_4')
// (23, 22, 'neigh_op_bnl_4')

reg n3002 = 0;
// (21, 21, 'local_g2_4')
// (21, 21, 'lutff_4/in_2')
// (21, 21, 'sp4_r_v_b_36')
// (21, 22, 'neigh_op_tnr_6')
// (21, 22, 'sp4_r_v_b_25')
// (21, 23, 'neigh_op_rgt_6')
// (21, 23, 'sp4_r_v_b_12')
// (21, 24, 'neigh_op_bnr_6')
// (21, 24, 'sp4_r_v_b_1')
// (22, 20, 'sp4_v_t_36')
// (22, 21, 'sp4_v_b_36')
// (22, 22, 'neigh_op_top_6')
// (22, 22, 'sp4_v_b_25')
// (22, 23, 'lutff_6/out')
// (22, 23, 'sp4_v_b_12')
// (22, 24, 'neigh_op_bot_6')
// (22, 24, 'sp4_v_b_1')
// (23, 22, 'neigh_op_tnl_6')
// (23, 23, 'neigh_op_lft_6')
// (23, 24, 'neigh_op_bnl_6')

wire n3003;
// (21, 21, 'neigh_op_tnr_3')
// (21, 22, 'neigh_op_rgt_3')
// (21, 23, 'neigh_op_bnr_3')
// (22, 21, 'neigh_op_top_3')
// (22, 22, 'lutff_3/out')
// (22, 23, 'neigh_op_bot_3')
// (23, 21, 'neigh_op_tnl_3')
// (23, 22, 'local_g1_3')
// (23, 22, 'lutff_global/cen')
// (23, 22, 'neigh_op_lft_3')
// (23, 23, 'neigh_op_bnl_3')

wire n3004;
// (21, 22, 'neigh_op_tnr_1')
// (21, 23, 'neigh_op_rgt_1')
// (21, 24, 'neigh_op_bnr_1')
// (22, 22, 'neigh_op_top_1')
// (22, 23, 'local_g0_2')
// (22, 23, 'lutff_1/out')
// (22, 23, 'lutff_global/cen')
// (22, 23, 'sp4_h_r_2')
// (22, 24, 'neigh_op_bot_1')
// (23, 22, 'neigh_op_tnl_1')
// (23, 23, 'neigh_op_lft_1')
// (23, 23, 'sp4_h_r_15')
// (23, 24, 'neigh_op_bnl_1')
// (24, 23, 'sp4_h_r_26')
// (25, 23, 'sp4_h_r_39')

reg n3005 = 0;
// (22, 1, 'neigh_op_tnr_2')
// (22, 2, 'neigh_op_rgt_2')
// (22, 3, 'local_g1_2')
// (22, 3, 'lutff_0/in_1')
// (22, 3, 'neigh_op_bnr_2')
// (23, 1, 'neigh_op_top_2')
// (23, 2, 'local_g1_2')
// (23, 2, 'lutff_2/in_1')
// (23, 2, 'lutff_2/out')
// (23, 3, 'neigh_op_bot_2')
// (24, 1, 'neigh_op_tnl_2')
// (24, 2, 'neigh_op_lft_2')
// (24, 3, 'neigh_op_bnl_2')

wire n3006;
// (22, 1, 'neigh_op_tnr_3')
// (22, 2, 'neigh_op_rgt_3')
// (22, 3, 'local_g0_3')
// (22, 3, 'lutff_6/in_1')
// (22, 3, 'neigh_op_bnr_3')
// (23, 1, 'neigh_op_top_3')
// (23, 2, 'lutff_3/out')
// (23, 3, 'neigh_op_bot_3')
// (24, 1, 'neigh_op_tnl_3')
// (24, 2, 'neigh_op_lft_3')
// (24, 3, 'neigh_op_bnl_3')

wire n3007;
// (22, 1, 'neigh_op_tnr_5')
// (22, 2, 'local_g3_5')
// (22, 2, 'lutff_5/in_1')
// (22, 2, 'neigh_op_rgt_5')
// (22, 3, 'neigh_op_bnr_5')
// (23, 1, 'neigh_op_top_5')
// (23, 2, 'lutff_5/out')
// (23, 3, 'neigh_op_bot_5')
// (24, 1, 'neigh_op_tnl_5')
// (24, 2, 'neigh_op_lft_5')
// (24, 3, 'neigh_op_bnl_5')

wire n3008;
// (22, 1, 'neigh_op_tnr_7')
// (22, 2, 'local_g2_7')
// (22, 2, 'lutff_6/in_1')
// (22, 2, 'neigh_op_rgt_7')
// (22, 3, 'neigh_op_bnr_7')
// (23, 1, 'neigh_op_top_7')
// (23, 2, 'lutff_7/out')
// (23, 3, 'neigh_op_bot_7')
// (24, 1, 'neigh_op_tnl_7')
// (24, 2, 'neigh_op_lft_7')
// (24, 3, 'neigh_op_bnl_7')

wire n3009;
// (22, 2, 'local_g2_4')
// (22, 2, 'lutff_1/in_1')
// (22, 2, 'neigh_op_tnr_4')
// (22, 3, 'neigh_op_rgt_4')
// (22, 4, 'neigh_op_bnr_4')
// (23, 2, 'neigh_op_top_4')
// (23, 3, 'lutff_4/out')
// (23, 4, 'neigh_op_bot_4')
// (24, 2, 'neigh_op_tnl_4')
// (24, 3, 'neigh_op_lft_4')
// (24, 4, 'neigh_op_bnl_4')

reg n3010 = 0;
// (22, 2, 'local_g2_5')
// (22, 2, 'lutff_7/in_0')
// (22, 2, 'neigh_op_tnr_5')
// (22, 3, 'neigh_op_rgt_5')
// (22, 4, 'neigh_op_bnr_5')
// (23, 2, 'neigh_op_top_5')
// (23, 3, 'local_g1_5')
// (23, 3, 'lutff_5/in_1')
// (23, 3, 'lutff_5/out')
// (23, 4, 'neigh_op_bot_5')
// (24, 2, 'neigh_op_tnl_5')
// (24, 3, 'neigh_op_lft_5')
// (24, 4, 'neigh_op_bnl_5')

reg n3011 = 0;
// (22, 2, 'local_g3_7')
// (22, 2, 'lutff_4/in_0')
// (22, 2, 'lutff_7/in_1')
// (22, 2, 'neigh_op_tnr_7')
// (22, 3, 'neigh_op_rgt_7')
// (22, 4, 'neigh_op_bnr_7')
// (23, 2, 'local_g0_7')
// (23, 2, 'lutff_0/in_1')
// (23, 2, 'neigh_op_top_7')
// (23, 3, 'local_g0_7')
// (23, 3, 'lutff_7/in_2')
// (23, 3, 'lutff_7/out')
// (23, 4, 'neigh_op_bot_7')
// (24, 2, 'neigh_op_tnl_7')
// (24, 3, 'neigh_op_lft_7')
// (24, 4, 'neigh_op_bnl_7')

wire n3012;
// (22, 2, 'neigh_op_tnr_0')
// (22, 3, 'local_g3_0')
// (22, 3, 'lutff_2/in_3')
// (22, 3, 'neigh_op_rgt_0')
// (22, 4, 'neigh_op_bnr_0')
// (23, 2, 'neigh_op_top_0')
// (23, 3, 'lutff_0/out')
// (23, 4, 'neigh_op_bot_0')
// (24, 2, 'neigh_op_tnl_0')
// (24, 3, 'neigh_op_lft_0')
// (24, 4, 'neigh_op_bnl_0')

wire n3013;
// (22, 2, 'neigh_op_tnr_2')
// (22, 3, 'local_g3_2')
// (22, 3, 'lutff_4/in_3')
// (22, 3, 'neigh_op_rgt_2')
// (22, 4, 'neigh_op_bnr_2')
// (23, 2, 'neigh_op_top_2')
// (23, 3, 'lutff_2/out')
// (23, 4, 'neigh_op_bot_2')
// (24, 2, 'neigh_op_tnl_2')
// (24, 3, 'neigh_op_lft_2')
// (24, 4, 'neigh_op_bnl_2')

reg n3014 = 0;
// (22, 7, 'local_g3_2')
// (22, 7, 'lutff_5/in_0')
// (22, 7, 'neigh_op_tnr_2')
// (22, 8, 'local_g2_2')
// (22, 8, 'lutff_1/in_3')
// (22, 8, 'lutff_2/in_0')
// (22, 8, 'lutff_4/in_2')
// (22, 8, 'neigh_op_rgt_2')
// (22, 9, 'neigh_op_bnr_2')
// (23, 7, 'local_g1_2')
// (23, 7, 'lutff_2/in_1')
// (23, 7, 'neigh_op_top_2')
// (23, 8, 'lutff_2/out')
// (23, 9, 'neigh_op_bot_2')
// (24, 7, 'neigh_op_tnl_2')
// (24, 8, 'neigh_op_lft_2')
// (24, 9, 'neigh_op_bnl_2')

reg n3015 = 0;
// (22, 7, 'neigh_op_tnr_1')
// (22, 8, 'local_g3_1')
// (22, 8, 'lutff_0/in_2')
// (22, 8, 'neigh_op_rgt_1')
// (22, 9, 'neigh_op_bnr_1')
// (23, 7, 'neigh_op_top_1')
// (23, 8, 'local_g2_1')
// (23, 8, 'lutff_1/out')
// (23, 8, 'lutff_2/in_3')
// (23, 9, 'neigh_op_bot_1')
// (24, 7, 'neigh_op_tnl_1')
// (24, 8, 'neigh_op_lft_1')
// (24, 9, 'neigh_op_bnl_1')

reg n3016 = 0;
// (22, 12, 'neigh_op_tnr_0')
// (22, 13, 'local_g3_0')
// (22, 13, 'lutff_7/in_2')
// (22, 13, 'neigh_op_rgt_0')
// (22, 14, 'neigh_op_bnr_0')
// (23, 12, 'neigh_op_top_0')
// (23, 13, 'lutff_0/out')
// (23, 14, 'neigh_op_bot_0')
// (24, 12, 'neigh_op_tnl_0')
// (24, 13, 'neigh_op_lft_0')
// (24, 14, 'neigh_op_bnl_0')

reg n3017 = 0;
// (22, 12, 'neigh_op_tnr_2')
// (22, 13, 'local_g2_2')
// (22, 13, 'lutff_7/in_3')
// (22, 13, 'neigh_op_rgt_2')
// (22, 14, 'neigh_op_bnr_2')
// (23, 12, 'neigh_op_top_2')
// (23, 13, 'lutff_2/out')
// (23, 14, 'neigh_op_bot_2')
// (24, 12, 'neigh_op_tnl_2')
// (24, 13, 'neigh_op_lft_2')
// (24, 14, 'neigh_op_bnl_2')

wire n3018;
// (22, 12, 'neigh_op_tnr_7')
// (22, 13, 'local_g3_7')
// (22, 13, 'lutff_4/in_0')
// (22, 13, 'neigh_op_rgt_7')
// (22, 14, 'neigh_op_bnr_7')
// (23, 12, 'neigh_op_top_7')
// (23, 13, 'lutff_7/out')
// (23, 14, 'local_g1_7')
// (23, 14, 'lutff_0/in_0')
// (23, 14, 'lutff_5/in_3')
// (23, 14, 'lutff_7/in_3')
// (23, 14, 'neigh_op_bot_7')
// (24, 12, 'neigh_op_tnl_7')
// (24, 13, 'local_g0_7')
// (24, 13, 'lutff_4/in_1')
// (24, 13, 'neigh_op_lft_7')
// (24, 14, 'neigh_op_bnl_7')

reg n3019 = 0;
// (22, 13, 'neigh_op_tnr_0')
// (22, 14, 'local_g3_0')
// (22, 14, 'lutff_1/in_2')
// (22, 14, 'neigh_op_rgt_0')
// (22, 15, 'local_g1_0')
// (22, 15, 'lutff_7/in_2')
// (22, 15, 'neigh_op_bnr_0')
// (23, 13, 'neigh_op_top_0')
// (23, 14, 'lutff_0/out')
// (23, 15, 'neigh_op_bot_0')
// (24, 13, 'neigh_op_tnl_0')
// (24, 14, 'neigh_op_lft_0')
// (24, 15, 'neigh_op_bnl_0')

wire n3020;
// (22, 13, 'neigh_op_tnr_1')
// (22, 14, 'neigh_op_rgt_1')
// (22, 15, 'neigh_op_bnr_1')
// (23, 13, 'neigh_op_top_1')
// (23, 14, 'local_g0_1')
// (23, 14, 'lutff_0/in_1')
// (23, 14, 'lutff_1/out')
// (23, 14, 'lutff_2/in_1')
// (23, 14, 'lutff_4/in_1')
// (23, 14, 'lutff_5/in_0')
// (23, 14, 'lutff_6/in_1')
// (23, 15, 'neigh_op_bot_1')
// (24, 13, 'neigh_op_tnl_1')
// (24, 14, 'neigh_op_lft_1')
// (24, 15, 'neigh_op_bnl_1')

reg n3021 = 0;
// (22, 13, 'neigh_op_tnr_2')
// (22, 14, 'local_g3_2')
// (22, 14, 'lutff_5/in_2')
// (22, 14, 'neigh_op_rgt_2')
// (22, 15, 'neigh_op_bnr_2')
// (23, 13, 'neigh_op_top_2')
// (23, 14, 'local_g3_2')
// (23, 14, 'lutff_2/in_3')
// (23, 14, 'lutff_2/out')
// (23, 15, 'local_g0_2')
// (23, 15, 'lutff_2/in_2')
// (23, 15, 'neigh_op_bot_2')
// (24, 13, 'neigh_op_tnl_2')
// (24, 14, 'neigh_op_lft_2')
// (24, 15, 'neigh_op_bnl_2')

reg n3022 = 0;
// (22, 13, 'neigh_op_tnr_4')
// (22, 14, 'neigh_op_rgt_4')
// (22, 15, 'local_g1_4')
// (22, 15, 'lutff_2/in_1')
// (22, 15, 'lutff_5/in_2')
// (22, 15, 'neigh_op_bnr_4')
// (23, 13, 'neigh_op_top_4')
// (23, 14, 'local_g2_4')
// (23, 14, 'lutff_4/in_2')
// (23, 14, 'lutff_4/out')
// (23, 15, 'neigh_op_bot_4')
// (24, 13, 'neigh_op_tnl_4')
// (24, 14, 'neigh_op_lft_4')
// (24, 15, 'neigh_op_bnl_4')

reg n3023 = 0;
// (22, 13, 'neigh_op_tnr_5')
// (22, 14, 'local_g3_5')
// (22, 14, 'lutff_3/in_1')
// (22, 14, 'neigh_op_rgt_5')
// (22, 15, 'neigh_op_bnr_5')
// (23, 13, 'neigh_op_top_5')
// (23, 14, 'lutff_5/out')
// (23, 15, 'local_g1_5')
// (23, 15, 'lutff_2/in_0')
// (23, 15, 'neigh_op_bot_5')
// (24, 13, 'neigh_op_tnl_5')
// (24, 14, 'neigh_op_lft_5')
// (24, 15, 'neigh_op_bnl_5')

reg n3024 = 0;
// (22, 13, 'neigh_op_tnr_6')
// (22, 14, 'neigh_op_rgt_6')
// (22, 15, 'local_g1_6')
// (22, 15, 'lutff_0/in_1')
// (22, 15, 'lutff_5/in_0')
// (22, 15, 'neigh_op_bnr_6')
// (23, 13, 'neigh_op_top_6')
// (23, 14, 'local_g2_6')
// (23, 14, 'lutff_6/in_0')
// (23, 14, 'lutff_6/out')
// (23, 15, 'neigh_op_bot_6')
// (24, 13, 'neigh_op_tnl_6')
// (24, 14, 'neigh_op_lft_6')
// (24, 15, 'neigh_op_bnl_6')

wire n3025;
// (22, 13, 'sp4_r_v_b_40')
// (22, 14, 'local_g1_5')
// (22, 14, 'lutff_global/s_r')
// (22, 14, 'neigh_op_tnr_0')
// (22, 14, 'sp4_r_v_b_29')
// (22, 15, 'local_g1_5')
// (22, 15, 'lutff_global/s_r')
// (22, 15, 'neigh_op_rgt_0')
// (22, 15, 'sp4_h_r_5')
// (22, 15, 'sp4_r_v_b_16')
// (22, 16, 'neigh_op_bnr_0')
// (22, 16, 'sp4_r_v_b_5')
// (23, 12, 'sp4_v_t_40')
// (23, 13, 'sp4_v_b_40')
// (23, 14, 'local_g0_0')
// (23, 14, 'lutff_2/in_2')
// (23, 14, 'lutff_4/in_0')
// (23, 14, 'lutff_6/in_2')
// (23, 14, 'lutff_7/in_1')
// (23, 14, 'neigh_op_top_0')
// (23, 14, 'sp4_v_b_29')
// (23, 15, 'lutff_0/out')
// (23, 15, 'sp4_h_r_16')
// (23, 15, 'sp4_v_b_16')
// (23, 16, 'neigh_op_bot_0')
// (23, 16, 'sp4_v_b_5')
// (24, 14, 'neigh_op_tnl_0')
// (24, 15, 'neigh_op_lft_0')
// (24, 15, 'sp4_h_r_29')
// (24, 16, 'neigh_op_bnl_0')
// (25, 15, 'sp4_h_r_40')

wire n3026;
// (22, 14, 'lutff_1/cout')
// (22, 14, 'lutff_2/in_3')

wire n3027;
// (22, 14, 'lutff_2/cout')
// (22, 14, 'lutff_3/in_3')

wire n3028;
// (22, 14, 'lutff_3/cout')
// (22, 14, 'lutff_4/in_3')

wire n3029;
// (22, 14, 'lutff_5/cout')
// (22, 14, 'lutff_6/in_3')

wire n3030;
// (22, 14, 'lutff_6/cout')
// (22, 14, 'lutff_7/in_3')

wire n3031;
// (22, 14, 'lutff_7/cout')
// (22, 15, 'carry_in')
// (22, 15, 'carry_in_mux')

wire n3032;
// (22, 14, 'neigh_op_tnr_2')
// (22, 15, 'neigh_op_rgt_2')
// (22, 16, 'neigh_op_bnr_2')
// (23, 14, 'local_g1_2')
// (23, 14, 'lutff_0/in_3')
// (23, 14, 'lutff_5/in_2')
// (23, 14, 'neigh_op_top_2')
// (23, 15, 'local_g1_2')
// (23, 15, 'lutff_0/in_3')
// (23, 15, 'lutff_2/out')
// (23, 16, 'neigh_op_bot_2')
// (24, 14, 'neigh_op_tnl_2')
// (24, 15, 'neigh_op_lft_2')
// (24, 16, 'neigh_op_bnl_2')

reg n3033 = 0;
// (22, 14, 'neigh_op_tnr_6')
// (22, 15, 'neigh_op_rgt_6')
// (22, 16, 'local_g0_6')
// (22, 16, 'lutff_2/in_2')
// (22, 16, 'neigh_op_bnr_6')
// (23, 14, 'neigh_op_top_6')
// (23, 15, 'lutff_6/out')
// (23, 16, 'neigh_op_bot_6')
// (24, 14, 'neigh_op_tnl_6')
// (24, 15, 'neigh_op_lft_6')
// (24, 16, 'neigh_op_bnl_6')

reg n3034 = 0;
// (22, 14, 'sp4_r_v_b_46')
// (22, 15, 'sp4_r_v_b_35')
// (22, 16, 'local_g3_6')
// (22, 16, 'lutff_2/in_1')
// (22, 16, 'sp4_r_v_b_22')
// (22, 17, 'sp4_r_v_b_11')
// (22, 18, 'sp4_r_v_b_38')
// (22, 19, 'neigh_op_tnr_7')
// (22, 19, 'sp4_r_v_b_27')
// (22, 20, 'neigh_op_rgt_7')
// (22, 20, 'sp4_r_v_b_14')
// (22, 21, 'neigh_op_bnr_7')
// (22, 21, 'sp4_r_v_b_3')
// (23, 13, 'sp4_v_t_46')
// (23, 14, 'sp4_v_b_46')
// (23, 15, 'sp4_v_b_35')
// (23, 16, 'sp4_v_b_22')
// (23, 17, 'sp4_v_b_11')
// (23, 17, 'sp4_v_t_38')
// (23, 18, 'sp4_v_b_38')
// (23, 19, 'neigh_op_top_7')
// (23, 19, 'sp4_v_b_27')
// (23, 20, 'lutff_7/out')
// (23, 20, 'sp4_v_b_14')
// (23, 21, 'neigh_op_bot_7')
// (23, 21, 'sp4_v_b_3')
// (24, 19, 'neigh_op_tnl_7')
// (24, 20, 'neigh_op_lft_7')
// (24, 21, 'neigh_op_bnl_7')

wire n3035;
// (22, 15, 'lutff_0/cout')
// (22, 15, 'lutff_1/in_3')

wire n3036;
// (22, 15, 'lutff_2/cout')
// (22, 15, 'lutff_3/in_3')

wire n3037;
// (22, 15, 'lutff_3/cout')
// (22, 15, 'lutff_4/in_3')

reg n3038 = 0;
// (22, 16, 'neigh_op_tnr_0')
// (22, 17, 'neigh_op_rgt_0')
// (22, 18, 'local_g1_0')
// (22, 18, 'lutff_7/in_0')
// (22, 18, 'neigh_op_bnr_0')
// (23, 16, 'neigh_op_top_0')
// (23, 17, 'lutff_0/out')
// (23, 18, 'neigh_op_bot_0')
// (24, 16, 'neigh_op_tnl_0')
// (24, 17, 'neigh_op_lft_0')
// (24, 18, 'neigh_op_bnl_0')

reg n3039 = 0;
// (22, 17, 'neigh_op_tnr_1')
// (22, 18, 'local_g3_1')
// (22, 18, 'lutff_2/in_2')
// (22, 18, 'neigh_op_rgt_1')
// (22, 19, 'neigh_op_bnr_1')
// (23, 17, 'neigh_op_top_1')
// (23, 18, 'lutff_1/out')
// (23, 19, 'neigh_op_bot_1')
// (24, 17, 'neigh_op_tnl_1')
// (24, 18, 'neigh_op_lft_1')
// (24, 19, 'neigh_op_bnl_1')

reg n3040 = 0;
// (22, 18, 'neigh_op_tnr_3')
// (22, 19, 'neigh_op_rgt_3')
// (22, 20, 'neigh_op_bnr_3')
// (23, 18, 'neigh_op_top_3')
// (23, 19, 'local_g2_3')
// (23, 19, 'lutff_1/in_2')
// (23, 19, 'lutff_3/out')
// (23, 20, 'neigh_op_bot_3')
// (24, 18, 'neigh_op_tnl_3')
// (24, 19, 'neigh_op_lft_3')
// (24, 20, 'neigh_op_bnl_3')

reg n3041 = 0;
// (22, 20, 'neigh_op_tnr_4')
// (22, 21, 'local_g3_4')
// (22, 21, 'lutff_4/in_3')
// (22, 21, 'neigh_op_rgt_4')
// (22, 22, 'neigh_op_bnr_4')
// (23, 20, 'neigh_op_top_4')
// (23, 21, 'lutff_4/out')
// (23, 22, 'neigh_op_bot_4')
// (24, 20, 'neigh_op_tnl_4')
// (24, 21, 'neigh_op_lft_4')
// (24, 22, 'neigh_op_bnl_4')

reg n3042 = 0;
// (22, 21, 'local_g0_2')
// (22, 21, 'lutff_4/in_0')
// (22, 21, 'sp4_h_r_10')
// (23, 20, 'neigh_op_tnr_1')
// (23, 21, 'neigh_op_rgt_1')
// (23, 21, 'sp4_h_r_23')
// (23, 22, 'neigh_op_bnr_1')
// (24, 20, 'neigh_op_top_1')
// (24, 21, 'lutff_1/out')
// (24, 21, 'sp4_h_r_34')
// (24, 22, 'neigh_op_bot_1')
// (25, 20, 'neigh_op_tnl_1')
// (25, 21, 'neigh_op_lft_1')
// (25, 21, 'sp4_h_r_47')
// (25, 22, 'neigh_op_bnl_1')

wire n3043;
// (23, 2, 'lutff_1/cout')
// (23, 2, 'lutff_2/in_3')

wire n3044;
// (23, 2, 'lutff_2/cout')
// (23, 2, 'lutff_3/in_3')

wire n3045;
// (23, 2, 'lutff_4/cout')
// (23, 2, 'lutff_5/in_3')

wire n3046;
// (23, 2, 'lutff_6/cout')
// (23, 2, 'lutff_7/in_3')

wire n3047;
// (23, 2, 'lutff_7/cout')
// (23, 3, 'carry_in')
// (23, 3, 'carry_in_mux')
// (23, 3, 'lutff_0/in_3')

wire n3048;
// (23, 3, 'lutff_1/cout')
// (23, 3, 'lutff_2/in_3')

wire n3049;
// (23, 3, 'lutff_3/cout')
// (23, 3, 'lutff_4/in_3')

wire n3050;
// (23, 3, 'lutff_4/cout')
// (23, 3, 'lutff_5/in_3')

wire n3051;
// (23, 12, 'lutff_1/cout')
// (23, 12, 'lutff_2/in_3')

reg n3052 = 0;
// (23, 12, 'neigh_op_tnr_4')
// (23, 13, 'local_g2_4')
// (23, 13, 'lutff_1/in_3')
// (23, 13, 'lutff_7/in_3')
// (23, 13, 'neigh_op_rgt_4')
// (23, 14, 'neigh_op_bnr_4')
// (24, 12, 'neigh_op_top_4')
// (24, 13, 'lutff_4/out')
// (24, 14, 'neigh_op_bot_4')
// (25, 12, 'neigh_op_tnl_4')
// (25, 13, 'neigh_op_lft_4')
// (25, 14, 'neigh_op_bnl_4')

reg n3053 = 0;
// (23, 15, 'neigh_op_tnr_5')
// (23, 16, 'neigh_op_rgt_5')
// (23, 17, 'local_g1_5')
// (23, 17, 'lutff_7/in_3')
// (23, 17, 'neigh_op_bnr_5')
// (24, 15, 'neigh_op_top_5')
// (24, 16, 'lutff_5/out')
// (24, 17, 'neigh_op_bot_5')
// (25, 15, 'neigh_op_tnl_5')
// (25, 16, 'neigh_op_lft_5')
// (25, 17, 'neigh_op_bnl_5')

reg n3054 = 0;
// (23, 16, 'neigh_op_tnr_3')
// (23, 17, 'local_g2_3')
// (23, 17, 'lutff_7/in_0')
// (23, 17, 'neigh_op_rgt_3')
// (23, 18, 'neigh_op_bnr_3')
// (24, 16, 'neigh_op_top_3')
// (24, 17, 'lutff_3/out')
// (24, 18, 'neigh_op_bot_3')
// (25, 16, 'neigh_op_tnl_3')
// (25, 17, 'neigh_op_lft_3')
// (25, 18, 'neigh_op_bnl_3')

reg n3055 = 0;
// (23, 18, 'neigh_op_tnr_0')
// (23, 19, 'local_g2_0')
// (23, 19, 'lutff_1/in_1')
// (23, 19, 'neigh_op_rgt_0')
// (23, 20, 'neigh_op_bnr_0')
// (24, 18, 'neigh_op_top_0')
// (24, 19, 'lutff_0/out')
// (24, 20, 'neigh_op_bot_0')
// (25, 18, 'neigh_op_tnl_0')
// (25, 19, 'neigh_op_lft_0')
// (25, 20, 'neigh_op_bnl_0')

wire open_0;
wire open_1;
wire open_2;
wire open_3;
wire open_4;
wire open_5;
wire open_6;
wire open_7;
wire open_8;
wire open_9;
wire open_10;
wire open_11;
wire open_12;
wire open_13;
wire open_14;
wire open_15;
wire open_16;
wire open_17;
wire open_18;
wire open_19;
wire open_20;
wire open_21;
wire open_22;
wire open_23;
wire open_24;
wire open_25;
wire open_26;
wire open_27;
wire open_28;
wire open_29;
wire open_30;
wire open_31;
wire open_32;
wire open_33;
wire open_34;
wire open_35;
wire open_36;
wire open_37;
wire open_38;
wire open_39;
wire open_40;
wire open_41;
wire open_42;
wire open_43;
wire open_44;
wire open_45;
wire open_46;
wire open_47;
wire open_48;
wire open_49;
wire open_50;
wire open_51;
wire open_52;
wire open_53;
wire open_54;
wire open_55;
wire open_56;
wire open_57;
wire open_58;
wire open_59;
wire open_60;
wire open_61;
wire open_62;
wire open_63;
wire open_64;
wire open_65;
wire open_66;
wire open_67;
wire open_68;
wire open_69;
wire open_70;
wire open_71;
wire open_72;
wire open_73;
wire open_74;
wire open_75;
wire n3056;
// (13, 1, 'lutff_2/cout')

wire n3057;
// (8, 15, 'lutff_5/cout')

wire n3058;
// (9, 20, 'lutff_0/cout')

wire n3059;
// (9, 16, 'lutff_2/cout')

wire n3060;
// (3, 14, 'lutff_0/cout')

wire n3061;
// (1, 6, 'lutff_3/cout')

wire n3062;
// (12, 1, 'lutff_1/cout')

wire n3063;
// (8, 19, 'lutff_1/cout')

wire n3064;
// (1, 21, 'lutff_0/cout')

wire n3065;
// (7, 15, 'lutff_3/cout')

wire n3066;
// (8, 7, 'lutff_4/cout')

wire n3067;
// (7, 8, 'lutff_0/cout')

wire n3068;
// (3, 17, 'lutff_0/cout')

wire n3069;
// (3, 14, 'lutff_3/cout')

wire n3070;
// (4, 18, 'lutff_2/cout')

wire n3071;
// (11, 1, 'lutff_0/cout')

wire n3072;
// (10, 18, 'lutff_0/cout')

wire n3073;
// (7, 15, 'lutff_6/cout')

wire n3074;
// (20, 1, 'lutff_0/cout')

wire n3075;
// (12, 3, 'lutff_4/cout')

wire n3076;
// (11, 1, 'lutff_3/cout')

wire n3077;
// (9, 18, 'lutff_0/cout')

wire n3078;
// (10, 18, 'lutff_3/cout')

wire n3079;
// (1, 8, 'lutff_0/cout')

wire n3080;
// (4, 13, 'lutff_2/cout')

wire n3081;
// (16, 19, 'lutff_0/cout')

wire n3082;
// (17, 11, 'lutff_0/cout')

wire n3083;
// (9, 16, 'lutff_1/cout')

wire n3084;
// (7, 9, 'lutff_5/cout')

wire n3085;
// (8, 19, 'lutff_0/cout')

wire n3086;
// (13, 1, 'lutff_4/cout')

wire n3087;
// (17, 14, 'lutff_0/cout')

wire n3088;
// (8, 7, 'lutff_3/cout')

wire n3089;
// (13, 23, 'lutff_0/cout')

wire n3090;
// (17, 6, 'lutff_1/cout')

wire n3091;
// (9, 16, 'lutff_4/cout')

wire n3092;
// (1, 6, 'lutff_5/cout')

wire n3093;
// (21, 7, 'lutff_0/cout')

wire n3094;
// (18, 1, 'lutff_0/cout')

wire n3095;
// (12, 1, 'lutff_3/cout')

wire n3096;
// (7, 15, 'lutff_5/cout')

wire n3097;
// (4, 18, 'lutff_4/cout')

wire n3098;
// (11, 1, 'lutff_2/cout')

wire n3099;
// (7, 18, 'lutff_6/cout')

wire n3100;
// (10, 18, 'lutff_2/cout')

wire n3101;
// (21, 13, 'lutff_0/cout')

wire n3102;
// (4, 21, 'lutff_0/cout')

wire n3103;
// (5, 6, 'lutff_0/cout')

wire n3104;
// (9, 17, 'lutff_1/cout')

wire n3105;
// (9, 18, 'lutff_2/cout')

wire n3106;
// (10, 18, 'lutff_5/cout')

wire n3107;
// (2, 9, 'lutff_0/cout')

wire n3108;
// (16, 19, 'lutff_2/cout')

wire n3109;
// (20, 14, 'lutff_0/cout')

wire n3110;
// (9, 16, 'lutff_3/cout')

wire n3111;
// (21, 8, 'lutff_0/cout')

wire n3112;
// (8, 19, 'lutff_2/cout')

wire n3113;
// (4, 8, 'lutff_0/cout')

wire n3114;
// (13, 1, 'lutff_6/cout')

wire n3115;
// (17, 18, 'lutff_0/cout')

wire n3116;
// (17, 6, 'lutff_3/cout')

wire n3117;
// (9, 12, 'lutff_0/cout')

wire n3118;
// (9, 16, 'lutff_6/cout')

wire n3119;
// (22, 15, 'lutff_1/cout')

wire n3120;
// (21, 7, 'lutff_2/cout')

wire n3121;
// (12, 1, 'lutff_5/cout')

wire n3122;
// (1, 13, 'lutff_0/cout')

wire n3123;
// (4, 18, 'lutff_6/cout')

wire n3124;
// (11, 1, 'lutff_4/cout')

wire n3125;
// (9, 18, 'lutff_1/cout')

wire n3126;
// (1, 16, 'lutff_0/cout')

wire n3127;
// (10, 18, 'lutff_4/cout')

wire n3128;
// (3, 13, 'lutff_1/cout')

wire n3129;
// (4, 13, 'lutff_3/cout')

wire n3130;
// (8, 17, 'lutff_1/cout')

wire n3131;
// (1, 19, 'lutff_0/cout')

wire n3132;
// (9, 18, 'lutff_4/cout')

wire n3133;
// (13, 1, 'lutff_5/cout')

wire n3134;
// (9, 16, 'lutff_5/cout')

wire n3135;
// (12, 21, 'lutff_0/cout')

wire n3136;
// (21, 8, 'lutff_2/cout')

wire n3137;
// (12, 2, 'lutff_0/cout')

wire n3138;
// (12, 1, 'lutff_4/cout')

wire n3139;
// (8, 19, 'lutff_4/cout')

wire n3140;
// (7, 20, 'lutff_0/cout')

wire n3141;
// (17, 6, 'lutff_5/cout')

wire n3142;
// (12, 12, 'lutff_3/cout')

wire n3143;
// (21, 7, 'lutff_4/cout')

wire n3144;
// (8, 15, 'lutff_1/cout')

wire n3145;
// (1, 17, 'lutff_0/cout')

wire n3146;
// (3, 13, 'lutff_0/cout')

wire n3147;
// (8, 17, 'lutff_0/cout')

wire n3148;
// (17, 19, 'lutff_4/cout')

wire n3149;
// (11, 1, 'lutff_6/cout')

wire n3150;
// (9, 18, 'lutff_3/cout')

wire n3151;
// (10, 18, 'lutff_6/cout')

wire n3152;
// (15, 18, 'lutff_0/cout')

wire n3153;
// (3, 13, 'lutff_3/cout')

wire n3154;
// (13, 2, 'lutff_0/cout')

wire n3155;
// (7, 18, 'lutff_0/cout')

wire n3156;
// (8, 17, 'lutff_3/cout')

wire n3157;
// (23, 2, 'lutff_0/cout')

wire n3158;
// (12, 22, 'lutff_0/cout')

wire n3159;
// (9, 18, 'lutff_6/cout')

wire n3160;
// (8, 19, 'lutff_3/cout')

wire n3161;
// (12, 3, 'lutff_0/cout')

wire n3162;
// (7, 16, 'lutff_1/cout')

wire n3163;
// (23, 2, 'lutff_3/cout')

wire n3164;
// (20, 6, 'lutff_0/cout')

wire n3165;
// (8, 15, 'lutff_0/cout')

wire n3166;
// (7, 19, 'lutff_1/cout')

wire n3167;
// (12, 1, 'lutff_6/cout')

wire n3168;
// (16, 18, 'lutff_0/cout')

wire n3169;
// (8, 19, 'lutff_6/cout')

wire n3170;
// (7, 20, 'lutff_2/cout')

wire n3171;
// (13, 19, 'lutff_0/cout')

wire n3172;
// (15, 16, 'lutff_0/cout')

wire n3173;
// (22, 14, 'lutff_4/cout')

wire n3174;
// (21, 3, 'lutff_0/cout')

wire n3175;
// (21, 7, 'lutff_6/cout')

wire n3176;
// (11, 1, 'lutff_5/cout')

wire n3177;
// (8, 15, 'lutff_3/cout')

wire n3178;
// (17, 13, 'lutff_0/cout')

wire n3179;
// (3, 13, 'lutff_2/cout')

wire n3180;
// (15, 19, 'lutff_0/cout')

wire n3181;
// (4, 21, 'lutff_3/cout')

wire n3182;
// (3, 9, 'lutff_4/cout')

wire n3183;
// (8, 17, 'lutff_2/cout')

wire n3184;
// (17, 19, 'lutff_6/cout')

wire n3185;
// (23, 3, 'lutff_0/cout')

wire n3186;
// (9, 18, 'lutff_5/cout')

wire n3187;
// (2, 21, 'lutff_0/cout')

wire n3188;
// (15, 18, 'lutff_2/cout')

wire n3189;
// (7, 18, 'lutff_2/cout')

wire n3190;
// (13, 17, 'lutff_0/cout')

wire n3191;
// (20, 7, 'lutff_0/cout')

wire n3192;
// (15, 15, 'lutff_0/cout')

wire n3193;
// (8, 19, 'lutff_5/cout')

wire n3194;
// (7, 20, 'lutff_1/cout')

wire n3195;
// (7, 9, 'lutff_0/cout')

wire n3196;
// (13, 20, 'lutff_0/cout')

wire n3197;
// (3, 18, 'lutff_0/cout')

wire n3198;
// (2, 8, 'lutff_0/cout')

wire n3199;
// (4, 19, 'lutff_2/cout')

wire n3200;
// (8, 15, 'lutff_2/cout')

wire n3201;
// (16, 18, 'lutff_2/cout')

wire n3202;
// (7, 20, 'lutff_4/cout')

wire n3203;
// (1, 6, 'lutff_0/cout')

wire n3204;
// (7, 15, 'lutff_0/cout')

wire n3205;
// (8, 7, 'lutff_1/cout')

wire n3206;
// (20, 5, 'lutff_0/cout')

wire n3207;
// (3, 13, 'lutff_4/cout')

wire n3208;
// (15, 19, 'lutff_2/cout')

wire n3209;
// (7, 18, 'lutff_1/cout')

wire n3210;
// (8, 17, 'lutff_4/cout')

wire n3211;
// (8, 9, 'lutff_0/cout')

wire n3212;
// (9, 22, 'lutff_0/cout')

wire n3213;
// (23, 3, 'lutff_2/cout')

wire n3214;
// (20, 8, 'lutff_0/cout')

wire n3215;
// (3, 8, 'lutff_0/cout')

wire n3216;
// (11, 11, 'lutff_0/cout')

wire n3217;
// (15, 18, 'lutff_4/cout')

wire n3218;
// (12, 3, 'lutff_1/cout')

wire n3219;
// (17, 7, 'lutff_1/cout')

wire n3220;
// (7, 18, 'lutff_4/cout')

wire n3221;
// (3, 19, 'lutff_0/cout')

wire n3222;
// (13, 17, 'lutff_2/cout')

wire n3223;
// (20, 7, 'lutff_2/cout')

wire n3224;
// (12, 14, 'lutff_0/cout')

wire n3225;
// (7, 20, 'lutff_3/cout')

wire n3226;
// (13, 1, 'lutff_1/cout')

wire n3227;
// (8, 15, 'lutff_4/cout')

wire n3228;
// (8, 7, 'lutff_0/cout')

wire n3229;
// (16, 18, 'lutff_4/cout')

wire n3230;
// (7, 20, 'lutff_6/cout')

wire n3231;
// (1, 6, 'lutff_2/cout')

wire n3232;
// (12, 1, 'lutff_0/cout')

wire n3233;
// (23, 12, 'lutff_0/cout')

wire n3234;
// (7, 15, 'lutff_2/cout')

wire n3235;
// (3, 13, 'lutff_6/cout')

wire n3236;
// (15, 19, 'lutff_4/cout')

wire n3237;
// (7, 18, 'lutff_3/cout')

wire n3238;
// (8, 17, 'lutff_6/cout')

wire n3239;
// (10, 19, 'lutff_0/cout')

wire n3240;
// (20, 8, 'lutff_2/cout')

wire n3241;
// (11, 11, 'lutff_2/cout')

wire n3242;
// (15, 15, 'lutff_1/cout')

wire n3243;
// (15, 18, 'lutff_6/cout')

wire n3244;
// (12, 3, 'lutff_3/cout')

wire n3245;
// (17, 19, 'lutff_0/cout')

wire n3246;
// (17, 7, 'lutff_3/cout')

wire n3247;
// (13, 17, 'lutff_4/cout')

wire n3248;
// (20, 7, 'lutff_4/cout')

wire n3249;
// (13, 1, 'lutff_0/cout')

wire n3250;
// (18, 6, 'lutff_0/cout')

wire n3251;
// (4, 12, 'lutff_0/cout')

wire n3252;
// (4, 13, 'lutff_1/cout')

wire n3253;
// (7, 20, 'lutff_5/cout')

wire n3254;
// (9, 16, 'lutff_0/cout')

wire n3255;
// (1, 6, 'lutff_1/cout')

wire n3256;
// (2, 19, 'lutff_0/cout')

wire n3257;
// (13, 1, 'lutff_3/cout')

wire n3258;
// (7, 15, 'lutff_1/cout')

wire n3259;
// (8, 15, 'lutff_6/cout')

wire n3260;
// (8, 7, 'lutff_2/cout')

wire n3261;
// (16, 18, 'lutff_6/cout')

wire n3262;
// (13, 15, 'lutff_0/cout')

wire n3263;
// (3, 14, 'lutff_1/cout')

wire n3264;
// (4, 18, 'lutff_0/cout')

wire n3265;
// (8, 17, 'lutff_5/cout')

wire n3266;
// (12, 1, 'lutff_2/cout')

wire n3267;
// (5, 11, 'lutff_0/cout')

wire n3268;
// (1, 20, 'lutff_0/cout')

wire n3269;
// (7, 15, 'lutff_4/cout')

wire n3270;
// (22, 14, 'lutff_0/cout')

wire n3271;
// (12, 3, 'lutff_2/cout')

wire n3272;
// (2, 6, 'lutff_0/cout')

wire n3273;
// (11, 1, 'lutff_1/cout')

wire n3274;
// (7, 18, 'lutff_5/cout')

wire n3275;
// (10, 18, 'lutff_1/cout')

wire n3276;
// (23, 2, 'lutff_5/cout')

wire n3277;
// (20, 8, 'lutff_4/cout')

wire n3278;
// (2, 17, 'lutff_0/cout')

wire n3279;
// (4, 13, 'lutff_0/cout')

wire n3280;
// (12, 3, 'lutff_5/cout')

wire n3281;
// (17, 19, 'lutff_2/cout')

wire n3282;
// (13, 17, 'lutff_6/cout')

wire n3283;
// (1, 8, 'lutff_1/cout')

wire n3284;
// (20, 7, 'lutff_6/cout')

wire n3285;
// (13, 1, 'lutff_2/out')

wire n3286;
// (13, 1, 'lutff_2/lout')

wire n3287;
// (2, 8, 'lutff_3/lout')

wire n3288;
// (4, 19, 'lutff_5/lout')

wire n3289;
// (14, 22, 'lutff_5/lout')

wire n3290;
// (14, 14, 'lutff_1/lout')

wire n3291;
// (3, 7, 'lutff_6/lout')

wire n3292;
// (11, 10, 'lutff_7/lout')

wire n3293;
// (12, 6, 'lutff_5/lout')

wire n3294;
// (15, 13, 'lutff_4/lout')

wire n3295;
// (5, 16, 'lutff_3/lout')

wire n3296;
// (4, 20, 'lutff_6/lout')

wire n3297;
// (4, 12, 'lutff_2/lout')

wire n3298;
// (14, 15, 'lutff_2/lout')

wire n3299;
// (8, 16, 'lutff_1/lout')

wire n3300;
// (2, 4, 'lutff_5/lout')

wire n3301;
// (22, 4, 'lutff_6/lout')

wire n3302;
// (14, 18, 'lutff_7/lout')

wire n3303;
// (11, 2, 'lutff_2/lout')

wire n3304;
// (8, 15, 'lutff_5/out')

wire n3305;
// (8, 15, 'lutff_5/lout')

wire n3306;
// (15, 14, 'lutff_5/lout')

wire n3307;
// (15, 6, 'lutff_1/lout')

wire n3308;
// (5, 9, 'lutff_0/lout')

wire n3309;
// (24, 13, 'lutff_4/lout')

wire n3310;
// (12, 2, 'lutff_7/lout')

wire n3311;
// (5, 8, 'lutff_4/lout')

wire n3312;
// (16, 19, 'lutff_1/out')

wire n3313;
// (16, 19, 'lutff_1/lout')

wire n3314;
// (4, 4, 'lutff_3/lout')

wire n3315;
// (11, 3, 'lutff_3/lout')

wire n3316;
// (16, 18, 'lutff_5/out')

wire n3317;
// (16, 18, 'lutff_5/lout')

wire n3318;
// (1, 18, 'lutff_0/lout')

wire n3319;
// (20, 22, 'lutff_4/lout')

wire n3320;
// (9, 20, 'lutff_0/out')

wire n3321;
// (9, 20, 'lutff_0/lout')

wire n3322;
// (9, 20, 'carry_in_mux')

// Carry-In for (9 20)
assign n3322 = 1;

wire n3323;
// (5, 1, 'lutff_1/lout')

wire n3324;
// (7, 20, 'lutff_7/out')

wire n3325;
// (7, 20, 'lutff_7/lout')

wire n3326;
// (17, 9, 'lutff_4/lout')

wire n3327;
// (7, 12, 'lutff_3/lout')

wire n3328;
// (8, 8, 'lutff_1/lout')

wire n3329;
// (5, 4, 'lutff_6/lout')

wire n3330;
// (16, 11, 'lutff_2/lout')

wire n3331;
// (16, 14, 'lutff_7/lout')

wire n3332;
// (17, 10, 'lutff_5/lout')

wire n3333;
// (7, 13, 'lutff_4/lout')

wire n3334;
// (17, 2, 'lutff_1/lout')

wire n3335;
// (7, 5, 'lutff_0/lout')

wire n3336;
// (5, 5, 'lutff_7/lout')

wire n3337;
// (9, 16, 'lutff_2/out')

wire n3338;
// (9, 16, 'lutff_2/lout')

wire n3339;
// (4, 1, 'lutff_6/lout')

wire n3340;
// (14, 3, 'lutff_4/lout')

wire n3341;
// (8, 4, 'lutff_3/lout')

wire n3342;
// (16, 7, 'lutff_4/lout')

wire n3343;
// (13, 19, 'lutff_5/lout')

wire n3344;
// (20, 18, 'lutff_5/lout')

wire n3345;
// (3, 14, 'lutff_0/out')

wire n3346;
// (3, 14, 'lutff_0/lout')

wire n3347;
// (3, 14, 'carry_in_mux')

// Carry-In for (3 14)
assign n3347 = 1;

wire n3348;
// (1, 14, 'lutff_7/lout')

wire n3349;
// (1, 6, 'lutff_3/out')

wire n3350;
// (1, 6, 'lutff_3/lout')

wire n3351;
// (10, 12, 'lutff_4/lout')

wire n3352;
// (9, 8, 'lutff_3/lout')

wire n3353;
// (13, 20, 'lutff_6/lout')

wire n3354;
// (2, 18, 'lutff_1/lout')

wire n3355;
// (21, 22, 'lutff_5/lout')

wire n3356;
// (11, 17, 'lutff_0/lout')

wire n3357;
// (18, 16, 'lutff_0/lout')

wire n3358;
// (3, 18, 'lutff_6/lout')

wire n3359;
// (10, 5, 'lutff_1/lout')

wire n3360;
// (9, 1, 'lutff_0/lout')

wire n3361;
// (2, 19, 'lutff_2/lout')

wire n3362;
// (7, 1, 'lutff_7/lout')

wire n3363;
// (3, 15, 'lutff_0/lout')

wire n3364;
// (11, 18, 'lutff_1/lout')

wire n3365;
// (11, 21, 'lutff_6/lout')

wire n3366;
// (12, 17, 'lutff_4/lout')

wire n3367;
// (12, 9, 'lutff_0/lout')

wire n3368;
// (3, 10, 'lutff_7/lout')

wire n3369;
// (22, 12, 'lutff_0/lout')

wire n3370;
// (3, 2, 'lutff_3/lout')

wire n3371;
// (18, 11, 'lutff_6/lout')

wire n3372;
// (15, 16, 'lutff_5/lout')

wire n3373;
// (8, 18, 'lutff_0/out')

wire n3374;
// (8, 18, 'lutff_0/lout')

wire n3375;
// (11, 13, 'lutff_7/lout')

wire n3376;
// (18, 12, 'lutff_7/lout')

wire n3377;
// (11, 5, 'lutff_3/lout')

wire n3378;
// (18, 4, 'lutff_3/lout')

wire n3379;
// (12, 1, 'lutff_1/out')

wire n3380;
// (12, 1, 'lutff_1/lout')

wire n3381;
// (5, 19, 'lutff_3/lout')

wire n3382;
// (4, 15, 'lutff_2/lout')

wire n3383;
// (12, 4, 'lutff_6/lout')

wire n3384;
// (8, 19, 'lutff_1/out')

wire n3385;
// (8, 19, 'lutff_1/lout')

wire n3386;
// (2, 7, 'lutff_5/lout')

wire n3387;
// (22, 7, 'lutff_6/lout')

wire n3388;
// (3, 3, 'lutff_3/lout')

wire n3389;
// (21, 3, 'lutff_5/lout')

wire n3390;
// (14, 21, 'lutff_7/lout')

wire n3391;
// (11, 6, 'lutff_4/lout')

wire n3392;
// (15, 17, 'lutff_5/lout')

wire n3393;
// (15, 9, 'lutff_1/lout')

wire n3394;
// (5, 12, 'lutff_0/lout')

wire n3395;
// (17, 21, 'lutff_5/lout')

wire n3396;
// (12, 5, 'lutff_7/lout')

wire n3397;
// (14, 14, 'lutff_4/lout')

wire n3398;
// (14, 6, 'lutff_0/lout')

wire n3399;
// (1, 21, 'lutff_0/out')

wire n3400;
// (1, 21, 'lutff_0/lout')

wire n3401;
// (1, 21, 'carry_in_mux')

// Carry-In for (1 21)
assign n3401 = 1;

wire n3402;
// (23, 12, 'lutff_1/lout')

wire n3403;
// (8, 14, 'lutff_7/lout')

wire n3404;
// (20, 17, 'lutff_0/lout')

wire n3405;
// (7, 15, 'lutff_3/out')

wire n3406;
// (7, 15, 'lutff_3/lout')

wire n3407;
// (5, 7, 'lutff_6/lout')

wire n3408;
// (9, 19, 'lutff_3/lout')

wire n3409;
// (4, 3, 'lutff_5/lout')

wire n3410;
// (8, 7, 'lutff_4/out')

wire n3411;
// (8, 7, 'lutff_4/lout')

wire n3412;
// (16, 9, 'lutff_3/lout')

wire n3413;
// (20, 21, 'lutff_6/lout')

wire n3414;
// (17, 13, 'lutff_5/lout')

wire n3415;
// (17, 5, 'lutff_1/lout')

wire n3416;
// (20, 13, 'lutff_2/lout')

wire n3417;
// (7, 8, 'lutff_0/out')

wire n3418;
// (7, 8, 'lutff_0/lout')

wire n3419;
// (7, 8, 'carry_in_mux')

// Carry-In for (7 8)
assign n3419 = 1;

wire n3420;
// (5, 8, 'lutff_7/lout')

wire n3421;
// (18, 18, 'lutff_0/lout')

wire n3422;
// (4, 4, 'lutff_6/lout')

wire n3423;
// (7, 11, 'lutff_5/lout')

wire n3424;
// (13, 23, 'lutff_1/lout')

wire n3425;
// (16, 10, 'lutff_4/lout')

wire n3426;
// (13, 22, 'lutff_5/lout')

wire n3427;
// (17, 6, 'lutff_2/out')

wire n3428;
// (17, 6, 'lutff_2/lout')

wire n3429;
// (14, 2, 'lutff_7/lout')

wire n3430;
// (3, 17, 'lutff_0/out')

wire n3431;
// (3, 17, 'lutff_0/lout')

wire n3432;
// (3, 17, 'carry_in_mux')

// Carry-In for (3 17)
assign n3432 = 1;

wire n3433;
// (10, 16, 'lutff_0/lout')

wire n3434;
// (1, 17, 'lutff_7/lout')

wire n3435;
// (17, 9, 'lutff_7/lout')

wire n3436;
// (1, 9, 'lutff_3/lout')

wire n3437;
// (7, 4, 'lutff_2/lout')

wire n3438;
// (9, 11, 'lutff_3/lout')

wire n3439;
// (16, 3, 'lutff_1/lout')

wire n3440;
// (13, 15, 'lutff_2/lout')

wire n3441;
// (7, 3, 'lutff_6/lout')

wire n3442;
// (10, 11, 'lutff_7/lout')

wire n3443;
// (13, 18, 'lutff_7/lout')

wire n3444;
// (3, 21, 'lutff_6/lout')

wire n3445;
// (10, 8, 'lutff_1/lout')

wire n3446;
// (22, 22, 'lutff_3/lout')

wire n3447;
// (9, 7, 'lutff_5/lout')

wire n3448;
// (13, 11, 'lutff_4/lout')

wire n3449;
// (21, 21, 'lutff_7/lout')

wire n3450;
// (3, 14, 'lutff_3/lout')

wire n3451;
// (11, 16, 'lutff_2/lout')

wire n3452;
// (12, 12, 'lutff_0/out')

wire n3453;
// (12, 12, 'lutff_0/lout')

wire n3454;
// (12, 12, 'carry_in_mux')

// Carry-In for (12 12)
assign n3454 = 0;

wire n3455;
// (22, 15, 'lutff_0/out')

wire n3456;
// (22, 15, 'lutff_0/lout')

wire n3457;
// (3, 13, 'lutff_7/lout')

wire n3458;
// (10, 12, 'lutff_7/lout')

wire n3459;
// (10, 4, 'lutff_3/lout')

wire n3460;
// (9, 8, 'lutff_6/lout')

wire n3461;
// (2, 18, 'lutff_4/lout')

wire n3462;
// (21, 14, 'lutff_4/lout')

wire n3463;
// (11, 17, 'lutff_3/lout')

wire n3464;
// (8, 21, 'lutff_0/lout')

wire n3465;
// (13, 3, 'lutff_5/lout')

wire n3466;
// (18, 7, 'lutff_3/lout')

wire n3467;
// (15, 20, 'lutff_6/lout')

wire n3468;
// (15, 12, 'lutff_2/lout')

wire n3469;
// (4, 18, 'lutff_2/lout')

wire n3470;
// (2, 10, 'lutff_5/lout')

wire n3471;
// (5, 18, 'lutff_6/lout')

wire n3472;
// (2, 2, 'lutff_1/lout')

wire n3473;
// (21, 6, 'lutff_5/lout')

wire n3474;
// (14, 16, 'lutff_3/lout')

wire n3475;
// (11, 1, 'lutff_0/out')

wire n3476;
// (11, 1, 'lutff_0/lout')

wire n3477;
// (11, 1, 'carry_in_mux')

// Carry-In for (11 1)
assign n3477 = 1;

wire n3478;
// (5, 15, 'lutff_0/lout')

wire n3479;
// (3, 2, 'lutff_6/lout')

wire n3480;
// (23, 15, 'lutff_2/lout')

wire n3481;
// (11, 4, 'lutff_5/lout')

wire n3482;
// (12, 8, 'lutff_7/lout')

wire n3483;
// (2, 3, 'lutff_2/lout')

wire n3484;
// (24, 14, 'lutff_5/lout')

wire n3485;
// (4, 14, 'lutff_4/lout')

wire n3486;
// (14, 9, 'lutff_0/lout')

wire n3487;
// (11, 5, 'lutff_6/lout')

wire n3488;
// (8, 17, 'lutff_7/out')

wire n3489;
// (8, 17, 'lutff_7/lout')

wire n3490;
// (17, 8, 'lutff_2/lout')

wire n3491;
// (10, 18, 'lutff_0/out')

wire n3492;
// (10, 18, 'lutff_0/lout')

wire n3493;
// (10, 18, 'carry_in_mux')

// Carry-In for (10 18)
assign n3493 = 1;

wire n3494;
// (9, 22, 'lutff_3/lout')

wire n3495;
// (17, 11, 'lutff_7/lout')

wire n3496;
// (4, 6, 'lutff_5/lout')

wire n3497;
// (7, 14, 'lutff_6/lout')

wire n3498;
// (8, 10, 'lutff_4/lout')

wire n3499;
// (8, 2, 'lutff_0/lout')

wire n3500;
// (1, 20, 'lutff_2/lout')

wire n3501;
// (14, 4, 'lutff_6/lout')

wire n3502;
// (10, 19, 'lutff_1/lout')

wire n3503;
// (5, 3, 'lutff_3/lout')

wire n3504;
// (23, 3, 'lutff_5/lout')

wire n3505;
// (9, 15, 'lutff_0/lout')

wire n3506;
// (17, 4, 'lutff_4/lout')

wire n3507;
// (8, 3, 'lutff_1/lout')

wire n3508;
// (16, 13, 'lutff_4/lout')

wire n3509;
// (4, 2, 'lutff_7/lout')

wire n3510;
// (16, 5, 'lutff_0/lout')

wire n3511;
// (14, 5, 'lutff_7/lout')

wire n3512;
// (18, 22, 'lutff_1/lout')

wire n3513;
// (1, 12, 'lutff_3/lout')

wire n3514;
// (7, 15, 'lutff_6/out')

wire n3515;
// (7, 15, 'lutff_6/lout')

wire n3516;
// (7, 7, 'lutff_2/lout')

wire n3517;
// (16, 6, 'lutff_1/lout')

wire n3518;
// (10, 14, 'lutff_7/lout')

wire n3519;
// (9, 10, 'lutff_6/lout')

wire n3520;
// (16, 9, 'lutff_6/lout')

wire n3521;
// (1, 5, 'lutff_0/lout')

wire n3522;
// (3, 16, 'lutff_2/lout')

wire n3523;
// (20, 1, 'lutff_0/out')

wire n3524;
// (20, 1, 'lutff_0/lout')

wire n3525;
// (20, 1, 'carry_in_mux')

// Carry-In for (20 1)
assign n3525 = 1;

wire n3526;
// (12, 15, 'lutff_1/lout')

wire n3527;
// (20, 4, 'lutff_5/lout')

wire n3528;
// (13, 14, 'lutff_4/lout')

wire n3529;
// (22, 13, 'lutff_2/lout')

wire n3530;
// (3, 17, 'lutff_3/lout')

wire n3531;
// (1, 9, 'lutff_6/lout')

wire n3532;
// (15, 23, 'lutff_1/lout')

wire n3533;
// (20, 5, 'lutff_6/lout')

wire n3534;
// (9, 11, 'lutff_6/lout')

wire n3535;
// (12, 19, 'lutff_7/lout')

wire n3536;
// (18, 10, 'lutff_4/lout')

wire n3537;
// (9, 3, 'lutff_2/lout')

wire n3538;
// (12, 11, 'lutff_3/lout')

wire n3539;
// (18, 2, 'lutff_0/lout')

wire n3540;
// (13, 7, 'lutff_1/lout')

wire n3541;
// (21, 17, 'lutff_4/lout')

wire n3542;
// (11, 20, 'lutff_3/lout')

wire n3543;
// (2, 13, 'lutff_6/lout')

wire n3544;
// (13, 6, 'lutff_5/lout')

wire n3545;
// (3, 1, 'lutff_0/lout')

wire n3546;
// (22, 14, 'lutff_2/lout')

wire n3547;
// (15, 15, 'lutff_2/out')

wire n3548;
// (15, 15, 'lutff_2/lout')

wire n3549;
// (3, 4, 'lutff_5/lout')

wire n3550;
// (15, 18, 'lutff_7/out')

wire n3551;
// (15, 18, 'lutff_7/lout')

wire n3552;
// (12, 3, 'lutff_4/out')

wire n3553;
// (12, 3, 'lutff_4/lout')

wire n3554;
// (5, 13, 'lutff_2/lout')

wire n3555;
// (4, 17, 'lutff_5/lout')

wire n3556;
// (4, 9, 'lutff_1/lout')

wire n3557;
// (3, 5, 'lutff_6/lout')

wire n3558;
// (16, 23, 'lutff_3/lout')

wire n3559;
// (17, 19, 'lutff_1/out')

wire n3560;
// (17, 19, 'lutff_1/lout')

wire n3561;
// (11, 7, 'lutff_5/lout')

wire n3562;
// (15, 11, 'lutff_4/lout')

wire n3563;
// (2, 6, 'lutff_2/lout')

wire n3564;
// (5, 14, 'lutff_3/lout')

wire n3565;
// (14, 20, 'lutff_4/lout')

wire n3566;
// (8, 21, 'lutff_3/lout')

wire n3567;
// (14, 12, 'lutff_0/lout')

wire n3568;
// (21, 5, 'lutff_7/lout')

wire n3569;
// (17, 20, 'lutff_2/lout')

wire n3570;
// (11, 8, 'lutff_6/lout')

wire n3571;
// (15, 12, 'lutff_5/lout')

wire n3572;
// (15, 4, 'lutff_1/lout')

wire n3573;
// (23, 14, 'lutff_4/lout')

wire n3574;
// (4, 10, 'lutff_1/lout')

wire n3575;
// (14, 13, 'lutff_1/lout')

wire n3576;
// (22, 2, 'lutff_5/lout')

wire n3577;
// (2, 2, 'lutff_4/lout')

wire n3578;
// (16, 24, 'lutff_3/lout')

wire n3579;
// (7, 17, 'lutff_6/lout')

wire n3580;
// (14, 16, 'lutff_6/lout')

wire n3581;
// (11, 1, 'lutff_3/out')

wire n3582;
// (11, 1, 'lutff_3/lout')

wire n3583;
// (8, 13, 'lutff_4/lout')

wire n3584;
// (8, 5, 'lutff_0/lout')

wire n3585;
// (23, 7, 'lutff_1/lout')

wire n3586;
// (9, 18, 'lutff_0/out')

wire n3587;
// (9, 18, 'lutff_0/lout')

wire n3588;
// (9, 18, 'carry_in_mux')

// Carry-In for (9 18)
assign n3588 = 1;

wire n3589;
// (7, 18, 'lutff_7/out')

wire n3590;
// (7, 18, 'lutff_7/lout')

wire n3591;
// (17, 7, 'lutff_4/out')

wire n3592;
// (17, 7, 'lutff_4/lout')

wire n3593;
// (7, 10, 'lutff_3/lout')

wire n3594;
// (9, 21, 'lutff_5/lout')

wire n3595;
// (8, 6, 'lutff_1/lout')

wire n3596;
// (16, 8, 'lutff_0/lout')

wire n3597;
// (20, 20, 'lutff_3/lout')

wire n3598;
// (14, 8, 'lutff_7/lout')

wire n3599;
// (8, 9, 'lutff_6/lout')

wire n3600;
// (17, 8, 'lutff_5/lout')

wire n3601;
// (10, 18, 'lutff_3/out')

wire n3602;
// (10, 18, 'lutff_3/lout')

wire n3603;
// (9, 22, 'lutff_6/lout')

wire n3604;
// (5, 2, 'lutff_5/lout')

wire n3605;
// (23, 2, 'lutff_7/lout')

wire n3606;
// (9, 14, 'lutff_2/lout')

wire n3607;
// (16, 12, 'lutff_6/lout')

wire n3608;
// (16, 4, 'lutff_2/lout')

wire n3609;
// (1, 8, 'lutff_0/out')

wire n3610;
// (1, 8, 'lutff_0/lout')

wire n3611;
// (1, 8, 'carry_in_mux')

// Carry-In for (1 8)
assign n3611 = 1;

wire n3612;
// (13, 17, 'lutff_5/out')

wire n3613;
// (13, 17, 'lutff_5/lout')

wire n3614;
// (8, 1, 'lutff_7/lout')

wire n3615;
// (12, 18, 'lutff_1/lout')

wire n3616;
// (20, 7, 'lutff_5/out')

wire n3617;
// (20, 7, 'lutff_5/lout')

wire n3618;
// (10, 10, 'lutff_4/lout')

wire n3619;
// (10, 2, 'lutff_0/lout')

wire n3620;
// (9, 6, 'lutff_3/lout')

wire n3621;
// (22, 16, 'lutff_2/lout')

wire n3622;
// (13, 9, 'lutff_0/lout')

wire n3623;
// (2, 16, 'lutff_1/lout')

wire n3624;
// (3, 20, 'lutff_3/lout')

wire n3625;
// (21, 20, 'lutff_5/lout')

wire n3626;
// (21, 12, 'lutff_1/lout')

wire n3627;
// (1, 12, 'lutff_6/lout')

wire n3628;
// (1, 4, 'lutff_2/lout')

wire n3629;
// (20, 8, 'lutff_6/lout')

wire n3630;
// (12, 22, 'lutff_7/lout')

wire n3631;
// (18, 13, 'lutff_4/lout')

wire n3632;
// (12, 14, 'lutff_3/lout')

wire n3633;
// (18, 5, 'lutff_0/lout')

wire n3634;
// (22, 17, 'lutff_3/lout')

wire n3635;
// (2, 17, 'lutff_2/lout')

wire n3636;
// (13, 10, 'lutff_1/lout')

wire n3637;
// (9, 2, 'lutff_5/lout')

wire n3638;
// (14, 23, 'lutff_0/out')

wire n3639;
// (14, 23, 'lutff_0/lout')

wire n3640;
// (14, 23, 'carry_in_mux')

// Carry-In for (14 23)
assign n3640 = 1;

wire n3641;
// (21, 16, 'lutff_7/lout')

wire n3642;
// (20, 1, 'lutff_3/lout')

wire n3643;
// (10, 3, 'lutff_0/lout')

wire n3644;
// (18, 6, 'lutff_1/lout')

wire n3645;
// (12, 7, 'lutff_0/lout')

wire n3646;
// (21, 13, 'lutff_1/out')

wire n3647;
// (21, 13, 'lutff_1/lout')

wire n3648;
// (18, 9, 'lutff_6/lout')

wire n3649;
// (12, 6, 'lutff_4/lout')

wire n3650;
// (5, 16, 'lutff_2/lout')

wire n3651;
// (11, 19, 'lutff_5/lout')

wire n3652;
// (4, 20, 'lutff_5/lout')

wire n3653;
// (4, 12, 'lutff_1/out')

wire n3654;
// (4, 12, 'lutff_1/lout')

wire n3655;
// (13, 5, 'lutff_7/lout')

wire n3656;
// (14, 15, 'lutff_1/lout')

wire n3657;
// (8, 16, 'lutff_0/out')

wire n3658;
// (8, 16, 'lutff_0/lout')

wire n3659;
// (2, 4, 'lutff_4/lout')

wire n3660;
// (3, 8, 'lutff_6/lout')

wire n3661;
// (17, 22, 'lutff_1/lout')

wire n3662;
// (18, 2, 'lutff_3/lout')

wire n3663;
// (5, 17, 'lutff_3/lout')

wire n3664;
// (15, 6, 'lutff_0/lout')

wire n3665;
// (4, 13, 'lutff_2/out')

wire n3666;
// (4, 13, 'lutff_2/lout')

wire n3667;
// (12, 2, 'lutff_6/lout')

wire n3668;
// (2, 5, 'lutff_5/lout')

wire n3669;
// (16, 19, 'lutff_0/lout')

wire n3670;
// (4, 16, 'lutff_7/lout')

wire n3671;
// (3, 1, 'lutff_3/lout')

wire n3672;
// (11, 11, 'lutff_6/lout')

wire n3673;
// (11, 3, 'lutff_2/lout')

wire n3674;
// (15, 15, 'lutff_5/lout')

wire n3675;
// (14, 11, 'lutff_3/lout')

wire n3676;
// (14, 19, 'lutff_7/lout')

wire n3677;
// (15, 7, 'lutff_1/lout')

wire n3678;
// (5, 10, 'lutff_0/lout')

wire n3679;
// (7, 21, 'lutff_2/lout')

wire n3680;
// (12, 3, 'lutff_7/lout')

wire n3681;
// (22, 5, 'lutff_5/lout')

wire n3682;
// (5, 13, 'lutff_5/lout')

wire n3683;
// (4, 9, 'lutff_4/lout')

wire n3684;
// (8, 8, 'lutff_0/lout')

wire n3685;
// (17, 11, 'lutff_0/out')

wire n3686;
// (17, 11, 'lutff_0/lout')

wire n3687;
// (17, 11, 'carry_in_mux')

// Carry-In for (17 11)
assign n3687 = 1;

wire n3688;
// (17, 10, 'lutff_4/lout')

wire n3689;
// (7, 13, 'lutff_3/lout')

wire n3690;
// (15, 2, 'lutff_7/lout')

wire n3691;
// (5, 5, 'lutff_6/lout')

wire n3692;
// (9, 16, 'lutff_1/out')

wire n3693;
// (9, 16, 'lutff_1/lout')

wire n3694;
// (4, 1, 'lutff_5/lout')

wire n3695;
// (14, 3, 'lutff_3/lout')

wire n3696;
// (8, 4, 'lutff_2/lout')

wire n3697;
// (16, 15, 'lutff_7/lout')

wire n3698;
// (20, 18, 'lutff_4/lout')

wire n3699;
// (17, 3, 'lutff_1/lout')

wire n3700;
// (7, 6, 'lutff_0/lout')

wire n3701;
// (9, 17, 'lutff_2/lout')

wire n3702;
// (7, 9, 'lutff_5/lout')

wire n3703;
// (8, 5, 'lutff_3/lout')

wire n3704;
// (13, 20, 'lutff_5/lout')

wire n3705;
// (20, 11, 'lutff_1/lout')

wire n3706;
// (10, 14, 'lutff_0/lout')

wire n3707;
// (18, 24, 'lutff_3/lout')

wire n3708;
// (17, 7, 'lutff_7/lout')

wire n3709;
// (3, 18, 'lutff_5/lout')

wire n3710;
// (16, 8, 'lutff_3/lout')

wire n3711;
// (2, 19, 'lutff_1/lout')

wire n3712;
// (7, 1, 'lutff_6/lout')

wire n3713;
// (13, 13, 'lutff_2/lout')

wire n3714;
// (18, 17, 'lutff_0/lout')

wire n3715;
// (1, 7, 'lutff_2/lout')

wire n3716;
// (13, 16, 'lutff_7/lout')

wire n3717;
// (3, 19, 'lutff_6/lout')

wire n3718;
// (20, 3, 'lutff_2/lout')

wire n3719;
// (11, 21, 'lutff_5/lout')

wire n3720;
// (12, 17, 'lutff_3/lout')

wire n3721;
// (20, 6, 'lutff_7/lout')

wire n3722;
// (2, 20, 'lutff_2/lout')

wire n3723;
// (10, 9, 'lutff_6/lout')

wire n3724;
// (9, 5, 'lutff_5/lout')

wire n3725;
// (1, 8, 'lutff_3/lout')

wire n3726;
// (21, 19, 'lutff_7/lout')

wire n3727;
// (3, 11, 'lutff_1/lout')

wire n3728;
// (11, 14, 'lutff_2/lout')

wire n3729;
// (12, 18, 'lutff_4/lout')

wire n3730;
// (12, 10, 'lutff_0/lout')

wire n3731;
// (10, 10, 'lutff_7/lout')

wire n3732;
// (10, 2, 'lutff_3/lout')

wire n3733;
// (18, 12, 'lutff_6/lout')

wire n3734;
// (9, 6, 'lutff_6/lout')

wire n3735;
// (18, 4, 'lutff_2/lout')

wire n3736;
// (22, 16, 'lutff_5/lout')

wire n3737;
// (22, 8, 'lutff_1/lout')

wire n3738;
// (21, 12, 'lutff_4/lout')

wire n3739;
// (21, 4, 'lutff_0/lout')

wire n3740;
// (8, 19, 'lutff_0/out')

wire n3741;
// (8, 19, 'lutff_0/lout')

wire n3742;
// (8, 19, 'carry_in_mux')

// Carry-In for (8 19)
assign n3742 = 1;

wire n3743;
// (3, 3, 'lutff_2/lout')

wire n3744;
// (18, 13, 'lutff_7/lout')

wire n3745;
// (18, 5, 'lutff_3/lout')

wire n3746;
// (5, 20, 'lutff_3/lout')

wire n3747;
// (17, 21, 'lutff_4/lout')

wire n3748;
// (12, 5, 'lutff_6/lout')

wire n3749;
// (8, 20, 'lutff_1/lout')

wire n3750;
// (13, 1, 'lutff_4/out')

wire n3751;
// (13, 1, 'lutff_4/lout')

wire n3752;
// (2, 8, 'lutff_5/lout')

wire n3753;
// (4, 19, 'lutff_7/lout')

wire n3754;
// (14, 14, 'lutff_3/lout')

wire n3755;
// (15, 10, 'lutff_1/lout')

wire n3756;
// (12, 6, 'lutff_7/lout')

wire n3757;
// (15, 13, 'lutff_6/lout')

wire n3758;
// (5, 16, 'lutff_5/lout')

wire n3759;
// (4, 12, 'lutff_4/lout')

wire n3760;
// (14, 15, 'lutff_4/lout')

wire n3761;
// (2, 4, 'lutff_7/lout')

wire n3762;
// (23, 13, 'lutff_1/lout')

wire n3763;
// (17, 14, 'lutff_0/out')

wire n3764;
// (17, 14, 'lutff_0/lout')

wire n3765;
// (17, 14, 'carry_in_mux')

// Carry-In for (17 14)
assign n3765 = 1;

wire n3766;
// (11, 2, 'lutff_4/lout')

wire n3767;
// (8, 15, 'lutff_7/out')

wire n3768;
// (8, 15, 'lutff_7/lout')

wire n3769;
// (8, 7, 'lutff_3/out')

wire n3770;
// (8, 7, 'lutff_3/lout')

wire n3771;
// (15, 6, 'lutff_3/lout')

wire n3772;
// (5, 8, 'lutff_6/lout')

wire n3773;
// (13, 23, 'lutff_0/out')

wire n3774;
// (13, 23, 'lutff_0/lout')

wire n3775;
// (13, 23, 'carry_in_mux')

// Carry-In for (13 23)
assign n3775 = 1;

wire n3776;
// (16, 18, 'lutff_7/out')

wire n3777;
// (16, 18, 'lutff_7/lout')

wire n3778;
// (16, 10, 'lutff_3/lout')

wire n3779;
// (17, 6, 'lutff_1/lout')

wire n3780;
// (14, 2, 'lutff_6/lout')

wire n3781;
// (9, 20, 'lutff_2/lout')

wire n3782;
// (5, 1, 'lutff_3/lout')

wire n3783;
// (17, 9, 'lutff_6/lout')

wire n3784;
// (18, 19, 'lutff_0/lout')

wire n3785;
// (7, 12, 'lutff_5/lout')

wire n3786;
// (7, 4, 'lutff_1/lout')

wire n3787;
// (8, 8, 'lutff_3/lout')

wire n3788;
// (16, 11, 'lutff_4/lout')

wire n3789;
// (16, 3, 'lutff_0/lout')

wire n3790;
// (20, 14, 'lutff_1/out')

wire n3791;
// (20, 14, 'lutff_1/lout')

wire n3792;
// (17, 10, 'lutff_7/lout')

wire n3793;
// (17, 2, 'lutff_3/lout')

wire n3794;
// (3, 21, 'lutff_5/lout')

wire n3795;
// (7, 5, 'lutff_2/lout')

wire n3796;
// (9, 16, 'lutff_4/out')

wire n3797;
// (9, 16, 'lutff_4/lout')

wire n3798;
// (12, 20, 'lutff_4/lout')

wire n3799;
// (14, 3, 'lutff_6/lout')

wire n3800;
// (16, 7, 'lutff_6/lout')

wire n3801;
// (13, 19, 'lutff_7/lout')

wire n3802;
// (3, 14, 'lutff_2/out')

wire n3803;
// (3, 14, 'lutff_2/lout')

wire n3804;
// (1, 6, 'lutff_5/lout')

wire n3805;
// (10, 12, 'lutff_6/lout')

wire n3806;
// (10, 4, 'lutff_2/lout')

wire n3807;
// (9, 8, 'lutff_5/lout')

wire n3808;
// (2, 18, 'lutff_3/lout')

wire n3809;
// (13, 12, 'lutff_4/lout')

wire n3810;
// (13, 4, 'lutff_0/lout')

wire n3811;
// (21, 14, 'lutff_3/lout')

wire n3812;
// (11, 17, 'lutff_2/lout')

wire n3813;
// (12, 13, 'lutff_0/lout')

wire n3814;
// (20, 2, 'lutff_4/lout')

wire n3815;
// (18, 7, 'lutff_2/lout')

wire n3816;
// (22, 19, 'lutff_5/lout')

wire n3817;
// (2, 19, 'lutff_4/lout')

wire n3818;
// (2, 11, 'lutff_0/lout')

wire n3819;
// (21, 15, 'lutff_4/lout')

wire n3820;
// (11, 18, 'lutff_3/lout')

wire n3821;
// (21, 7, 'lutff_0/out')

wire n3822;
// (21, 7, 'lutff_0/lout')

wire n3823;
// (21, 7, 'carry_in_mux')

// Carry-In for (21 7)
assign n3823 = 1;

wire n3824;
// (8, 22, 'lutff_0/lout')

wire n3825;
// (18, 8, 'lutff_3/lout')

wire n3826;
// (12, 9, 'lutff_2/lout')

wire n3827;
// (3, 2, 'lutff_5/lout')

wire n3828;
// (12, 8, 'lutff_6/lout')

wire n3829;
// (15, 16, 'lutff_7/lout')

wire n3830;
// (2, 3, 'lutff_1/lout')

wire n3831;
// (4, 14, 'lutff_3/lout')

wire n3832;
// (14, 17, 'lutff_3/lout')

wire n3833;
// (8, 18, 'lutff_2/lout')

wire n3834;
// (18, 1, 'lutff_0/out')

wire n3835;
// (18, 1, 'lutff_0/lout')

wire n3836;
// (18, 1, 'carry_in_mux')

// Carry-In for (18 1)
assign n3836 = 1;

wire n3837;
// (17, 17, 'lutff_1/lout')

wire n3838;
// (11, 5, 'lutff_5/lout')

wire n3839;
// (12, 1, 'lutff_3/out')

wire n3840;
// (12, 1, 'lutff_3/lout')

wire n3841;
// (5, 19, 'lutff_5/lout')

wire n3842;
// (5, 11, 'lutff_1/lout')

wire n3843;
// (4, 15, 'lutff_4/lout')

wire n3844;
// (4, 7, 'lutff_0/lout')

wire n3845;
// (2, 7, 'lutff_7/lout')

wire n3846;
// (14, 10, 'lutff_0/lout')

wire n3847;
// (3, 3, 'lutff_5/lout')

wire n3848;
// (21, 3, 'lutff_7/lout')

wire n3849;
// (11, 6, 'lutff_6/lout')

wire n3850;
// (15, 9, 'lutff_3/lout')

wire n3851;
// (5, 12, 'lutff_2/lout')

wire n3852;
// (4, 8, 'lutff_1/lout')

wire n3853;
// (14, 6, 'lutff_2/lout')

wire n3854;
// (8, 3, 'lutff_0/lout')

wire n3855;
// (1, 21, 'lutff_2/lout')

wire n3856;
// (15, 1, 'lutff_4/lout')

wire n3857;
// (7, 15, 'lutff_5/out')

wire n3858;
// (7, 15, 'lutff_5/lout')

wire n3859;
// (7, 7, 'lutff_1/lout')

wire n3860;
// (9, 19, 'lutff_5/lout')

wire n3861;
// (4, 3, 'lutff_7/lout')

wire n3862;
// (16, 6, 'lutff_0/lout')

wire n3863;
// (8, 7, 'lutff_6/lout')

wire n3864;
// (16, 9, 'lutff_5/lout')

wire n3865;
// (17, 13, 'lutff_7/lout')

wire n3866;
// (17, 5, 'lutff_3/lout')

wire n3867;
// (20, 13, 'lutff_4/lout')

wire n3868;
// (7, 8, 'lutff_2/lout')

wire n3869;
// (18, 18, 'lutff_2/lout')

wire n3870;
// (16, 10, 'lutff_6/lout')

wire n3871;
// (13, 22, 'lutff_7/lout')

wire n3872;
// (13, 14, 'lutff_3/lout')

wire n3873;
// (3, 17, 'lutff_2/lout')

wire n3874;
// (18, 19, 'lutff_3/lout')

wire n3875;
// (1, 9, 'lutff_5/lout')

wire n3876;
// (20, 5, 'lutff_5/lout')

wire n3877;
// (9, 11, 'lutff_5/lout')

wire n3878;
// (13, 15, 'lutff_4/lout')

wire n3879;
// (13, 7, 'lutff_0/lout')

wire n3880;
// (1, 2, 'lutff_2/lout')

wire n3881;
// (10, 8, 'lutff_3/lout')

wire n3882;
// (12, 20, 'lutff_7/lout')

wire n3883;
// (9, 4, 'lutff_2/lout')

wire n3884;
// (22, 14, 'lutff_1/lout')

wire n3885;
// (2, 14, 'lutff_0/lout')

wire n3886;
// (13, 8, 'lutff_1/lout')

wire n3887;
// (9, 7, 'lutff_7/lout')

wire n3888;
// (13, 11, 'lutff_6/lout')

wire n3889;
// (10, 1, 'lutff_0/lout')

wire n3890;
// (11, 16, 'lutff_4/lout')

wire n3891;
// (12, 12, 'lutff_2/lout')

wire n3892;
// (22, 15, 'lutff_2/out')

wire n3893;
// (22, 15, 'lutff_2/lout')

wire n3894;
// (3, 5, 'lutff_5/lout')

wire n3895;
// (10, 4, 'lutff_5/lout')

wire n3896;
// (15, 19, 'lutff_7/lout')

wire n3897;
// (22, 18, 'lutff_7/lout')

wire n3898;
// (2, 6, 'lutff_1/out')

wire n3899;
// (2, 6, 'lutff_1/lout')

wire n3900;
// (5, 14, 'lutff_2/lout')

wire n3901;
// (21, 14, 'lutff_6/lout')

wire n3902;
// (11, 9, 'lutff_1/lout')

wire n3903;
// (8, 21, 'lutff_2/lout')

wire n3904;
// (13, 3, 'lutff_7/lout')

wire n3905;
// (3, 6, 'lutff_6/lout')

wire n3906;
// (17, 20, 'lutff_1/lout')

wire n3907;
// (11, 8, 'lutff_5/lout')

wire n3908;
// (18, 7, 'lutff_5/lout')

wire n3909;
// (15, 12, 'lutff_4/lout')

wire n3910;
// (15, 4, 'lutff_0/lout')

wire n3911;
// (4, 18, 'lutff_4/lout')

wire n3912;
// (4, 10, 'lutff_0/lout')

wire n3913;
// (8, 22, 'lutff_3/lout')

wire n3914;
// (2, 10, 'lutff_7/lout')

wire n3915;
// (14, 13, 'lutff_0/lout')

wire n3916;
// (22, 2, 'lutff_4/lout')

wire n3917;
// (2, 2, 'lutff_3/lout')

wire n3918;
// (21, 6, 'lutff_7/lout')

wire n3919;
// (11, 1, 'lutff_2/out')

wire n3920;
// (11, 1, 'lutff_2/lout')

wire n3921;
// (5, 15, 'lutff_2/lout')

wire n3922;
// (17, 24, 'lutff_7/lout')

wire n3923;
// (17, 16, 'lutff_3/lout')

wire n3924;
// (11, 4, 'lutff_7/lout')

wire n3925;
// (4, 11, 'lutff_1/lout')

wire n3926;
// (22, 3, 'lutff_5/lout')

wire n3927;
// (2, 3, 'lutff_4/lout')

wire n3928;
// (4, 14, 'lutff_6/lout')

wire n3929;
// (7, 18, 'lutff_6/out')

wire n3930;
// (7, 18, 'lutff_6/lout')

wire n3931;
// (14, 17, 'lutff_6/lout')

wire n3932;
// (14, 9, 'lutff_2/lout')

wire n3933;
// (15, 5, 'lutff_0/lout')

wire n3934;
// (8, 6, 'lutff_0/lout')

wire n3935;
// (20, 20, 'lutff_2/lout')

wire n3936;
// (8, 9, 'lutff_5/lout')

wire n3937;
// (17, 8, 'lutff_4/lout')

wire n3938;
// (10, 18, 'lutff_2/out')

wire n3939;
// (10, 18, 'lutff_2/lout')

wire n3940;
// (9, 22, 'lutff_5/lout')

wire n3941;
// (5, 2, 'lutff_4/lout')

wire n3942;
// (9, 14, 'lutff_1/lout')

wire n3943;
// (4, 6, 'lutff_7/lout')

wire n3944;
// (8, 10, 'lutff_6/lout')

wire n3945;
// (8, 2, 'lutff_2/lout')

wire n3946;
// (1, 20, 'lutff_4/lout')

wire n3947;
// (16, 12, 'lutff_5/lout')

wire n3948;
// (10, 19, 'lutff_3/lout')

wire n3949;
// (5, 3, 'lutff_5/lout')

wire n3950;
// (9, 15, 'lutff_2/lout')

wire n3951;
// (18, 21, 'lutff_2/lout')

wire n3952;
// (17, 4, 'lutff_6/lout')

wire n3953;
// (23, 3, 'lutff_7/lout')

wire n3954;
// (16, 13, 'lutff_6/lout')

wire n3955;
// (16, 5, 'lutff_2/lout')

wire n3956;
// (3, 20, 'lutff_2/lout')

wire n3957;
// (20, 9, 'lutff_1/lout')

wire n3958;
// (18, 22, 'lutff_3/lout')

wire n3959;
// (1, 12, 'lutff_5/lout')

wire n3960;
// (7, 7, 'lutff_4/lout')

wire n3961;
// (12, 22, 'lutff_6/lout')

wire n3962;
// (22, 17, 'lutff_2/lout')

wire n3963;
// (2, 17, 'lutff_1/out')

wire n3964;
// (2, 17, 'lutff_1/lout')

wire n3965;
// (13, 10, 'lutff_0/lout')

wire n3966;
// (10, 6, 'lutff_5/lout')

wire n3967;
// (9, 2, 'lutff_4/lout')

wire n3968;
// (3, 16, 'lutff_4/lout')

wire n3969;
// (20, 1, 'lutff_2/lout')

wire n3970;
// (12, 15, 'lutff_3/lout')

wire n3971;
// (20, 4, 'lutff_7/lout')

wire n3972;
// (10, 7, 'lutff_6/lout')

wire n3973;
// (21, 13, 'lutff_0/out')

wire n3974;
// (21, 13, 'lutff_0/lout')

wire n3975;
// (21, 13, 'carry_in_mux')

// Carry-In for (21 13)
assign n3975 = 1;

wire n3976;
// (24, 21, 'lutff_1/lout')

wire n3977;
// (4, 21, 'lutff_0/out')

wire n3978;
// (4, 21, 'lutff_0/lout')

wire n3979;
// (4, 21, 'carry_in_mux')

// Carry-In for (4 21)
assign n3979 = 1;

wire n3980;
// (13, 14, 'lutff_6/lout')

wire n3981;
// (2, 21, 'lutff_7/lout')

wire n3982;
// (22, 13, 'lutff_4/lout')

wire n3983;
// (3, 17, 'lutff_5/lout')

wire n3984;
// (3, 9, 'lutff_1/lout')

wire n3985;
// (11, 19, 'lutff_4/lout')

wire n3986;
// (18, 10, 'lutff_6/lout')

wire n3987;
// (9, 3, 'lutff_4/lout')

wire n3988;
// (18, 2, 'lutff_2/lout')

wire n3989;
// (21, 17, 'lutff_6/lout')

wire n3990;
// (21, 9, 'lutff_2/lout')

wire n3991;
// (11, 12, 'lutff_1/lout')

wire n3992;
// (13, 6, 'lutff_7/lout')

wire n3993;
// (2, 5, 'lutff_4/lout')

wire n3994;
// (3, 1, 'lutff_2/lout')

wire n3995;
// (14, 19, 'lutff_6/lout')

wire n3996;
// (15, 15, 'lutff_4/lout')

wire n3997;
// (3, 4, 'lutff_7/lout')

wire n3998;
// (15, 7, 'lutff_0/lout')

wire n3999;
// (7, 21, 'lutff_1/lout')

wire n4000;
// (12, 3, 'lutff_6/out')

wire n4001;
// (12, 3, 'lutff_6/lout')

wire n4002;
// (22, 5, 'lutff_4/lout')

wire n4003;
// (5, 13, 'lutff_4/lout')

wire n4004;
// (4, 17, 'lutff_7/lout')

wire n4005;
// (4, 9, 'lutff_3/lout')

wire n4006;
// (15, 8, 'lutff_1/lout')

wire n4007;
// (17, 19, 'lutff_3/out')

wire n4008;
// (17, 19, 'lutff_3/lout')

wire n4009;
// (11, 7, 'lutff_7/lout')

wire n4010;
// (15, 11, 'lutff_6/lout')

wire n4011;
// (2, 6, 'lutff_4/lout')

wire n4012;
// (5, 14, 'lutff_5/lout')

wire n4013;
// (14, 12, 'lutff_2/lout')

wire n4014;
// (17, 12, 'lutff_0/lout')

wire n4015;
// (15, 4, 'lutff_3/lout')

wire n4016;
// (23, 14, 'lutff_6/lout')

wire n4017;
// (5, 6, 'lutff_0/out')

wire n4018;
// (5, 6, 'lutff_0/lout')

wire n4019;
// (5, 6, 'carry_in_mux')

// Carry-In for (5 6)
assign n4019 = 1;

wire n4020;
// (15, 3, 'lutff_7/lout')

wire n4021;
// (22, 2, 'lutff_7/lout')

wire n4022;
// (16, 16, 'lutff_1/lout')

wire n4023;
// (9, 17, 'lutff_1/lout')

wire n4024;
// (13, 21, 'lutff_0/lout')

wire n4025;
// (7, 9, 'lutff_4/lout')

wire n4026;
// (8, 13, 'lutff_6/lout')

wire n4027;
// (8, 5, 'lutff_2/lout')

wire n4028;
// (20, 11, 'lutff_0/lout')

wire n4029;
// (9, 18, 'lutff_2/out')

wire n4030;
// (9, 18, 'lutff_2/lout')

wire n4031;
// (17, 7, 'lutff_6/lout')

wire n4032;
// (7, 10, 'lutff_5/lout')

wire n4033;
// (7, 2, 'lutff_1/lout')

wire n4034;
// (9, 21, 'lutff_7/lout')

wire n4035;
// (8, 6, 'lutff_3/lout')

wire n4036;
// (1, 16, 'lutff_1/lout')

wire n4037;
// (16, 8, 'lutff_2/lout')

wire n4038;
// (20, 20, 'lutff_5/lout')

wire n4039;
// (20, 12, 'lutff_1/lout')

wire n4040;
// (10, 15, 'lutff_0/lout')

wire n4041;
// (17, 8, 'lutff_7/lout')

wire n4042;
// (10, 18, 'lutff_5/out')

wire n4043;
// (10, 18, 'lutff_5/lout')

wire n4044;
// (3, 19, 'lutff_5/lout')

wire n4045;
// (5, 2, 'lutff_7/lout')

wire n4046;
// (9, 14, 'lutff_4/lout')

wire n4047;
// (2, 20, 'lutff_1/lout')

wire n4048;
// (1, 8, 'lutff_2/out')

wire n4049;
// (1, 8, 'lutff_2/lout')

wire n4050;
// (13, 17, 'lutff_7/out')

wire n4051;
// (13, 17, 'lutff_7/lout')

wire n4052;
// (3, 11, 'lutff_0/lout')

wire n4053;
// (1, 11, 'lutff_7/lout')

wire n4054;
// (12, 18, 'lutff_3/lout')

wire n4055;
// (20, 7, 'lutff_7/out')

wire n4056;
// (20, 7, 'lutff_7/lout')

wire n4057;
// (10, 10, 'lutff_6/lout')

wire n4058;
// (10, 2, 'lutff_2/lout')

wire n4059;
// (9, 6, 'lutff_5/lout')

wire n4060;
// (22, 16, 'lutff_4/lout')

wire n4061;
// (2, 16, 'lutff_3/lout')

wire n4062;
// (3, 20, 'lutff_5/lout')

wire n4063;
// (13, 9, 'lutff_2/lout')

wire n4064;
// (3, 12, 'lutff_1/lout')

wire n4065;
// (22, 8, 'lutff_0/lout')

wire n4066;
// (21, 20, 'lutff_7/lout')

wire n4067;
// (21, 12, 'lutff_3/lout')

wire n4068;
// (1, 4, 'lutff_4/lout')

wire n4069;
// (18, 13, 'lutff_6/lout')

wire n4070;
// (12, 14, 'lutff_5/lout')

wire n4071;
// (18, 5, 'lutff_2/lout')

wire n4072;
// (2, 17, 'lutff_4/lout')

wire n4073;
// (13, 10, 'lutff_3/lout')

wire n4074;
// (2, 9, 'lutff_0/out')

wire n4075;
// (2, 9, 'lutff_0/lout')

wire n4076;
// (2, 9, 'carry_in_mux')

// Carry-In for (2 9)
assign n4076 = 1;

wire n4077;
// (9, 2, 'lutff_7/lout')

wire n4078;
// (11, 15, 'lutff_1/lout')

wire n4079;
// (14, 23, 'lutff_2/lout')

wire n4080;
// (8, 20, 'lutff_0/out')

wire n4081;
// (8, 20, 'lutff_0/lout')

wire n4082;
// (10, 3, 'lutff_2/lout')

wire n4083;
// (18, 6, 'lutff_3/lout')

wire n4084;
// (3, 7, 'lutff_7/lout')

wire n4085;
// (21, 13, 'lutff_3/lout')

wire n4086;
// (12, 6, 'lutff_6/lout')

wire n4087;
// (5, 16, 'lutff_4/lout')

wire n4088;
// (4, 20, 'lutff_7/lout')

wire n4089;
// (23, 22, 'lutff_0/lout')

wire n4090;
// (4, 12, 'lutff_3/lout')

wire n4091;
// (14, 15, 'lutff_3/lout')

wire n4092;
// (8, 16, 'lutff_2/lout')

wire n4093;
// (2, 4, 'lutff_6/lout')

wire n4094;
// (22, 4, 'lutff_7/lout')

wire n4095;
// (15, 14, 'lutff_6/lout')

wire n4096;
// (5, 17, 'lutff_5/lout')

wire n4097;
// (15, 6, 'lutff_2/lout')

wire n4098;
// (2, 1, 'lutff_0/lout')

wire n4099;
// (5, 9, 'lutff_1/lout')

wire n4100;
// (4, 13, 'lutff_4/out')

wire n4101;
// (4, 13, 'lutff_4/lout')

wire n4102;
// (4, 5, 'lutff_0/lout')

wire n4103;
// (2, 5, 'lutff_7/lout')

wire n4104;
// (16, 19, 'lutff_2/lout')

wire n4105;
// (11, 3, 'lutff_4/lout')

wire n4106;
// (14, 11, 'lutff_5/lout')

wire n4107;
// (15, 7, 'lutff_3/lout')

wire n4108;
// (20, 22, 'lutff_5/lout')

wire n4109;
// (22, 5, 'lutff_7/lout')

wire n4110;
// (5, 1, 'lutff_2/lout')

wire n4111;
// (8, 8, 'lutff_2/lout')

wire n4112;
// (5, 4, 'lutff_7/lout')

wire n4113;
// (16, 11, 'lutff_3/lout')

wire n4114;
// (20, 14, 'lutff_0/out')

wire n4115;
// (20, 14, 'lutff_0/lout')

wire n4116;
// (20, 14, 'carry_in_mux')

// Carry-In for (20 14)
assign n4116 = 1;

wire n4117;
// (17, 10, 'lutff_6/lout')

wire n4118;
// (7, 13, 'lutff_5/lout')

wire n4119;
// (17, 2, 'lutff_2/lout')

wire n4120;
// (7, 5, 'lutff_1/lout')

wire n4121;
// (9, 16, 'lutff_3/out')

wire n4122;
// (9, 16, 'lutff_3/lout')

wire n4123;
// (1, 19, 'lutff_1/lout')

wire n4124;
// (4, 1, 'lutff_7/lout')

wire n4125;
// (20, 15, 'lutff_1/lout')

wire n4126;
// (14, 3, 'lutff_5/lout')

wire n4127;
// (8, 4, 'lutff_4/lout')

wire n4128;
// (16, 7, 'lutff_5/lout')

wire n4129;
// (20, 18, 'lutff_6/lout')

wire n4130;
// (17, 3, 'lutff_3/lout')

wire n4131;
// (7, 6, 'lutff_2/lout')

wire n4132;
// (10, 13, 'lutff_1/lout')

wire n4133;
// (9, 17, 'lutff_4/lout')

wire n4134;
// (9, 9, 'lutff_0/lout')

wire n4135;
// (7, 9, 'lutff_7/lout')

wire n4136;
// (13, 20, 'lutff_7/lout')

wire n4137;
// (13, 12, 'lutff_3/lout')

wire n4138;
// (20, 11, 'lutff_3/lout')

wire n4139;
// (18, 16, 'lutff_1/lout')

wire n4140;
// (20, 10, 'lutff_7/lout')

wire n4141;
// (3, 18, 'lutff_7/lout')

wire n4142;
// (22, 20, 'lutff_0/lout')

wire n4143;
// (9, 1, 'lutff_1/lout')

wire n4144;
// (2, 19, 'lutff_3/lout')

wire n4145;
// (13, 13, 'lutff_4/lout')

wire n4146;
// (22, 19, 'lutff_4/lout')

wire n4147;
// (3, 15, 'lutff_1/lout')

wire n4148;
// (21, 15, 'lutff_3/lout')

wire n4149;
// (11, 18, 'lutff_2/lout')

wire n4150;
// (1, 7, 'lutff_4/lout')

wire n4151;
// (12, 17, 'lutff_5/lout')

wire n4152;
// (18, 8, 'lutff_2/lout')

wire n4153;
// (2, 20, 'lutff_4/lout')

wire n4154;
// (12, 9, 'lutff_1/lout')

wire n4155;
// (22, 12, 'lutff_1/lout')

wire n4156;
// (2, 12, 'lutff_0/lout')

wire n4157;
// (18, 11, 'lutff_7/lout')

wire n4158;
// (21, 8, 'lutff_0/lout')

wire n4159;
// (9, 5, 'lutff_7/lout')

wire n4160;
// (3, 11, 'lutff_3/lout')

wire n4161;
// (11, 14, 'lutff_4/lout')

wire n4162;
// (12, 10, 'lutff_2/lout')

wire n4163;
// (10, 2, 'lutff_5/lout')

wire n4164;
// (22, 16, 'lutff_7/lout')

wire n4165;
// (5, 19, 'lutff_4/lout')

wire n4166;
// (22, 8, 'lutff_3/lout')

wire n4167;
// (21, 12, 'lutff_6/lout')

wire n4168;
// (21, 4, 'lutff_2/lout')

wire n4169;
// (4, 15, 'lutff_3/lout')

wire n4170;
// (8, 19, 'lutff_2/out')

wire n4171;
// (8, 19, 'lutff_2/lout')

wire n4172;
// (2, 7, 'lutff_6/lout')

wire n4173;
// (3, 3, 'lutff_4/lout')

wire n4174;
// (11, 6, 'lutff_5/lout')

wire n4175;
// (18, 5, 'lutff_5/lout')

wire n4176;
// (5, 20, 'lutff_5/lout')

wire n4177;
// (15, 9, 'lutff_2/lout')

wire n4178;
// (23, 20, 'lutff_7/lout')

wire n4179;
// (5, 12, 'lutff_1/lout')

wire n4180;
// (17, 21, 'lutff_6/lout')

wire n4181;
// (4, 8, 'lutff_0/out')

wire n4182;
// (4, 8, 'lutff_0/lout')

wire n4183;
// (4, 8, 'carry_in_mux')

// Carry-In for (4 8)
assign n4183 = 1;

wire n4184;
// (8, 20, 'lutff_3/lout')

wire n4185;
// (2, 8, 'lutff_7/lout')

wire n4186;
// (13, 1, 'lutff_6/out')

wire n4187;
// (13, 1, 'lutff_6/lout')

wire n4188;
// (16, 22, 'lutff_2/lout')

wire n4189;
// (17, 18, 'lutff_0/out')

wire n4190;
// (17, 18, 'lutff_0/lout')

wire n4191;
// (17, 18, 'carry_in_mux')

// Carry-In for (17 18)
assign n4191 = 1;

wire n4192;
// (14, 14, 'lutff_5/lout')

wire n4193;
// (14, 6, 'lutff_1/lout')

wire n4194;
// (15, 10, 'lutff_3/lout')

wire n4195;
// (23, 12, 'lutff_2/lout')

wire n4196;
// (7, 16, 'lutff_0/out')

wire n4197;
// (7, 16, 'lutff_0/lout')

wire n4198;
// (5, 16, 'lutff_7/lout')

wire n4199;
// (4, 12, 'lutff_6/lout')

wire n4200;
// (14, 15, 'lutff_6/lout')

wire n4201;
// (17, 14, 'lutff_2/lout')

wire n4202;
// (8, 7, 'lutff_5/out')

wire n4203;
// (8, 7, 'lutff_5/lout')

wire n4204;
// (17, 13, 'lutff_6/lout')

wire n4205;
// (20, 21, 'lutff_7/lout')

wire n4206;
// (20, 13, 'lutff_3/lout')

wire n4207;
// (7, 8, 'lutff_1/lout')

wire n4208;
// (14, 7, 'lutff_1/lout')

wire n4209;
// (4, 4, 'lutff_7/lout')

wire n4210;
// (7, 11, 'lutff_6/lout')

wire n4211;
// (13, 23, 'lutff_2/lout')

wire n4212;
// (16, 10, 'lutff_5/lout')

wire n4213;
// (17, 6, 'lutff_3/lout')

wire n4214;
// (16, 2, 'lutff_1/lout')

wire n4215;
// (9, 20, 'lutff_4/lout')

wire n4216;
// (5, 1, 'lutff_5/lout')

wire n4217;
// (9, 12, 'lutff_0/out')

wire n4218;
// (9, 12, 'lutff_0/lout')

wire n4219;
// (9, 12, 'carry_in_mux')

// Carry-In for (9 12)
assign n4219 = 1;

wire n4220;
// (18, 19, 'lutff_2/lout')

wire n4221;
// (7, 12, 'lutff_7/lout')

wire n4222;
// (8, 8, 'lutff_5/lout')

wire n4223;
// (7, 4, 'lutff_3/lout')

wire n4224;
// (16, 11, 'lutff_6/lout')

wire n4225;
// (16, 3, 'lutff_2/lout')

wire n4226;
// (20, 14, 'lutff_3/lout')

wire n4227;
// (17, 2, 'lutff_5/lout')

wire n4228;
// (3, 21, 'lutff_7/lout')

wire n4229;
// (1, 2, 'lutff_1/lout')

wire n4230;
// (9, 16, 'lutff_6/out')

wire n4231;
// (9, 16, 'lutff_6/lout')

wire n4232;
// (13, 8, 'lutff_0/lout')

wire n4233;
// (13, 11, 'lutff_5/lout')

wire n4234;
// (3, 14, 'lutff_4/lout')

wire n4235;
// (1, 6, 'lutff_7/lout')

wire n4236;
// (12, 12, 'lutff_1/lout')

wire n4237;
// (22, 15, 'lutff_1/lout')

wire n4238;
// (2, 15, 'lutff_0/lout')

wire n4239;
// (10, 4, 'lutff_4/lout')

wire n4240;
// (9, 8, 'lutff_7/lout')

wire n4241;
// (21, 11, 'lutff_0/lout')

wire n4242;
// (22, 18, 'lutff_6/lout')

wire n4243;
// (1, 3, 'lutff_1/lout')

wire n4244;
// (2, 18, 'lutff_5/lout')

wire n4245;
// (13, 12, 'lutff_6/lout')

wire n4246;
// (13, 4, 'lutff_2/lout')

wire n4247;
// (21, 14, 'lutff_5/lout')

wire n4248;
// (11, 9, 'lutff_0/lout')

wire n4249;
// (12, 13, 'lutff_2/lout')

wire n4250;
// (20, 2, 'lutff_6/lout')

wire n4251;
// (10, 5, 'lutff_5/lout')

wire n4252;
// (3, 6, 'lutff_5/lout')

wire n4253;
// (24, 19, 'lutff_0/lout')

wire n4254;
// (9, 1, 'lutff_4/lout')

wire n4255;
// (15, 20, 'lutff_7/lout')

wire n4256;
// (22, 19, 'lutff_7/lout')

wire n4257;
// (22, 11, 'lutff_3/lout')

wire n4258;
// (2, 11, 'lutff_2/lout')

wire n4259;
// (21, 7, 'lutff_2/lout')

wire n4260;
// (11, 10, 'lutff_1/lout')

wire n4261;
// (8, 22, 'lutff_2/lout')

wire n4262;
// (18, 8, 'lutff_5/lout')

wire n4263;
// (3, 2, 'lutff_7/lout')

wire n4264;
// (5, 15, 'lutff_1/lout')

wire n4265;
// (17, 16, 'lutff_2/lout')

wire n4266;
// (4, 11, 'lutff_0/lout')

wire n4267;
// (22, 3, 'lutff_4/lout')

wire n4268;
// (2, 3, 'lutff_3/lout')

wire n4269;
// (4, 14, 'lutff_5/lout')

wire n4270;
// (14, 17, 'lutff_5/lout')

wire n4271;
// (8, 18, 'lutff_4/lout')

wire n4272;
// (14, 9, 'lutff_1/lout')

wire n4273;
// (17, 17, 'lutff_3/lout')

wire n4274;
// (11, 5, 'lutff_7/lout')

wire n4275;
// (7, 19, 'lutff_0/out')

wire n4276;
// (7, 19, 'lutff_0/lout')

wire n4277;
// (12, 1, 'lutff_5/out')

wire n4278;
// (12, 1, 'lutff_5/lout')

wire n4279;
// (5, 19, 'lutff_7/lout')

wire n4280;
// (5, 11, 'lutff_3/lout')

wire n4281;
// (4, 15, 'lutff_6/lout')

wire n4282;
// (4, 7, 'lutff_2/lout')

wire n4283;
// (14, 10, 'lutff_2/lout')

wire n4284;
// (8, 11, 'lutff_1/lout')

wire n4285;
// (15, 9, 'lutff_5/lout')

wire n4286;
// (1, 20, 'lutff_3/lout')

wire n4287;
// (5, 4, 'lutff_0/lout')

wire n4288;
// (10, 19, 'lutff_2/lout')

wire n4289;
// (5, 3, 'lutff_4/lout')

wire n4290;
// (16, 14, 'lutff_1/lout')

wire n4291;
// (14, 6, 'lutff_4/lout')

wire n4292;
// (8, 3, 'lutff_2/lout')

wire n4293;
// (16, 13, 'lutff_5/lout')

wire n4294;
// (1, 13, 'lutff_0/out')

wire n4295;
// (1, 13, 'lutff_0/lout')

wire n4296;
// (1, 13, 'carry_in_mux')

// Carry-In for (1 13)
assign n4296 = 1;

wire n4297;
// (20, 17, 'lutff_4/lout')

wire n4298;
// (20, 9, 'lutff_0/lout')

wire n4299;
// (18, 22, 'lutff_2/lout')

wire n4300;
// (7, 15, 'lutff_7/out')

wire n4301;
// (7, 15, 'lutff_7/lout')

wire n4302;
// (7, 7, 'lutff_3/lout')

wire n4303;
// (9, 19, 'lutff_7/lout')

wire n4304;
// (16, 6, 'lutff_2/lout')

wire n4305;
// (16, 9, 'lutff_7/lout')

wire n4306;
// (20, 13, 'lutff_6/lout')

wire n4307;
// (7, 8, 'lutff_4/lout')

wire n4308;
// (20, 10, 'lutff_0/lout')

wire n4309;
// (2, 21, 'lutff_6/lout')

wire n4310;
// (13, 14, 'lutff_5/lout')

wire n4311;
// (3, 17, 'lutff_4/lout')

wire n4312;
// (3, 9, 'lutff_0/out')

wire n4313;
// (3, 9, 'lutff_0/lout')

wire n4314;
// (3, 9, 'carry_in_mux')

// Carry-In for (3 9)
assign n4314 = 0;

wire n4315;
// (18, 19, 'lutff_5/lout')

wire n4316;
// (20, 5, 'lutff_7/lout')

wire n4317;
// (9, 11, 'lutff_7/lout')

wire n4318;
// (4, 22, 'lutff_0/lout')

wire n4319;
// (9, 3, 'lutff_3/lout')

wire n4320;
// (13, 15, 'lutff_6/lout')

wire n4321;
// (13, 7, 'lutff_2/lout')

wire n4322;
// (21, 17, 'lutff_5/lout')

wire n4323;
// (3, 10, 'lutff_1/lout')

wire n4324;
// (11, 20, 'lutff_4/lout')

wire n4325;
// (11, 12, 'lutff_0/lout')

wire n4326;
// (1, 2, 'lutff_4/lout')

wire n4327;
// (18, 11, 'lutff_0/lout')

wire n4328;
// (10, 8, 'lutff_5/lout')

wire n4329;
// (9, 4, 'lutff_4/lout')

wire n4330;
// (22, 22, 'lutff_7/lout')

wire n4331;
// (22, 14, 'lutff_3/lout')

wire n4332;
// (2, 14, 'lutff_2/lout')

wire n4333;
// (21, 18, 'lutff_6/lout')

wire n4334;
// (21, 10, 'lutff_2/lout')

wire n4335;
// (11, 16, 'lutff_6/lout')

wire n4336;
// (12, 12, 'lutff_4/lout')

wire n4337;
// (18, 3, 'lutff_1/lout')

wire n4338;
// (12, 4, 'lutff_0/lout')

wire n4339;
// (3, 5, 'lutff_7/lout')

wire n4340;
// (15, 8, 'lutff_0/lout')

wire n4341;
// (22, 7, 'lutff_0/lout')

wire n4342;
// (15, 11, 'lutff_5/lout')

wire n4343;
// (2, 6, 'lutff_3/lout')

wire n4344;
// (5, 14, 'lutff_4/lout')

wire n4345;
// (8, 21, 'lutff_4/lout')

wire n4346;
// (17, 20, 'lutff_3/lout')

wire n4347;
// (11, 8, 'lutff_7/lout')

wire n4348;
// (15, 12, 'lutff_6/lout')

wire n4349;
// (15, 4, 'lutff_2/lout')

wire n4350;
// (4, 18, 'lutff_6/lout')

wire n4351;
// (4, 10, 'lutff_2/lout')

wire n4352;
// (14, 13, 'lutff_2/lout')

wire n4353;
// (8, 14, 'lutff_1/lout')

wire n4354;
// (2, 2, 'lutff_5/lout')

wire n4355;
// (22, 2, 'lutff_6/lout')

wire n4356;
// (16, 16, 'lutff_0/lout')

wire n4357;
// (14, 16, 'lutff_7/lout')

wire n4358;
// (11, 1, 'lutff_4/out')

wire n4359;
// (11, 1, 'lutff_4/lout')

wire n4360;
// (5, 15, 'lutff_4/lout')

wire n4361;
// (23, 15, 'lutff_6/lout')

wire n4362;
// (5, 7, 'lutff_0/lout')

wire n4363;
// (23, 7, 'lutff_2/lout')

wire n4364;
// (24, 3, 'lutff_0/lout')

wire n4365;
// (22, 3, 'lutff_7/lout')

wire n4366;
// (9, 18, 'lutff_1/out')

wire n4367;
// (9, 18, 'lutff_1/lout')

wire n4368;
// (16, 17, 'lutff_1/lout')

wire n4369;
// (14, 9, 'lutff_4/lout')

wire n4370;
// (8, 6, 'lutff_2/lout')

wire n4371;
// (1, 16, 'lutff_0/out')

wire n4372;
// (1, 16, 'lutff_0/lout')

wire n4373;
// (1, 16, 'carry_in_mux')

// Carry-In for (1 16)
assign n4373 = 1;

wire n4374;
// (20, 20, 'lutff_4/lout')

wire n4375;
// (8, 9, 'lutff_7/lout')

wire n4376;
// (20, 12, 'lutff_0/lout')

wire n4377;
// (17, 8, 'lutff_6/lout')

wire n4378;
// (10, 18, 'lutff_4/out')

wire n4379;
// (10, 18, 'lutff_4/lout')

wire n4380;
// (9, 22, 'lutff_7/lout')

wire n4381;
// (5, 2, 'lutff_6/lout')

wire n4382;
// (9, 14, 'lutff_3/lout')

wire n4383;
// (1, 17, 'lutff_1/out')

wire n4384;
// (1, 17, 'lutff_1/lout')

wire n4385;
// (8, 2, 'lutff_4/lout')

wire n4386;
// (1, 20, 'lutff_6/lout')

wire n4387;
// (16, 12, 'lutff_7/lout')

wire n4388;
// (16, 4, 'lutff_3/lout')

wire n4389;
// (10, 19, 'lutff_5/lout')

wire n4390;
// (7, 3, 'lutff_0/lout')

wire n4391;
// (10, 11, 'lutff_1/lout')

wire n4392;
// (5, 3, 'lutff_7/lout')

wire n4393;
// (9, 15, 'lutff_4/lout')

wire n4394;
// (16, 5, 'lutff_4/lout')

wire n4395;
// (17, 1, 'lutff_2/lout')

wire n4396;
// (3, 20, 'lutff_4/lout')

wire n4397;
// (3, 12, 'lutff_0/lout')

wire n4398;
// (1, 12, 'lutff_7/lout')

wire n4399;
// (18, 14, 'lutff_1/lout')

wire n4400;
// (1, 4, 'lutff_3/lout')

wire n4401;
// (21, 21, 'lutff_1/lout')

wire n4402;
// (12, 14, 'lutff_4/lout')

wire n4403;
// (22, 17, 'lutff_4/lout')

wire n4404;
// (2, 17, 'lutff_3/lout')

wire n4405;
// (13, 10, 'lutff_2/lout')

wire n4406;
// (3, 13, 'lutff_1/out')

wire n4407;
// (3, 13, 'lutff_1/lout')

wire n4408;
// (9, 2, 'lutff_6/lout')

wire n4409;
// (1, 5, 'lutff_4/lout')

wire n4410;
// (11, 15, 'lutff_0/lout')

wire n4411;
// (14, 23, 'lutff_1/lout')

wire n4412;
// (3, 16, 'lutff_6/lout')

wire n4413;
// (20, 1, 'lutff_4/lout')

wire n4414;
// (10, 3, 'lutff_1/lout')

wire n4415;
// (12, 15, 'lutff_5/lout')

wire n4416;
// (18, 6, 'lutff_2/lout')

wire n4417;
// (12, 7, 'lutff_1/lout')

wire n4418;
// (21, 13, 'lutff_2/lout')

wire n4419;
// (4, 21, 'lutff_2/lout')

wire n4420;
// (18, 9, 'lutff_7/lout')

wire n4421;
// (15, 20, 'lutff_0/lout')

wire n4422;
// (3, 9, 'lutff_3/lout')

wire n4423;
// (3, 8, 'lutff_7/lout')

wire n4424;
// (9, 3, 'lutff_6/lout')

wire n4425;
// (5, 17, 'lutff_4/lout')

wire n4426;
// (4, 13, 'lutff_3/out')

wire n4427;
// (4, 13, 'lutff_3/lout')

wire n4428;
// (11, 12, 'lutff_3/lout')

wire n4429;
// (2, 5, 'lutff_6/lout')

wire n4430;
// (3, 1, 'lutff_4/lout')

wire n4431;
// (11, 11, 'lutff_7/lout')

wire n4432;
// (23, 18, 'lutff_1/lout')

wire n4433;
// (14, 11, 'lutff_4/lout')

wire n4434;
// (15, 15, 'lutff_6/lout')

wire n4435;
// (15, 7, 'lutff_2/lout')

wire n4436;
// (5, 10, 'lutff_1/lout')

wire n4437;
// (7, 21, 'lutff_3/lout')

wire n4438;
// (8, 17, 'lutff_1/out')

wire n4439;
// (8, 17, 'lutff_1/lout')

wire n4440;
// (22, 5, 'lutff_6/lout')

wire n4441;
// (5, 13, 'lutff_6/lout')

wire n4442;
// (21, 1, 'lutff_5/lout')

wire n4443;
// (4, 9, 'lutff_5/lout')

wire n4444;
// (15, 8, 'lutff_3/lout')

wire n4445;
// (16, 23, 'lutff_7/lout')

wire n4446;
// (17, 19, 'lutff_5/out')

wire n4447;
// (17, 19, 'lutff_5/lout')

wire n4448;
// (17, 11, 'lutff_1/lout')

wire n4449;
// (7, 14, 'lutff_0/lout')

wire n4450;
// (2, 6, 'lutff_6/lout')

wire n4451;
// (14, 12, 'lutff_4/lout')

wire n4452;
// (14, 4, 'lutff_0/lout')

wire n4453;
// (1, 19, 'lutff_0/out')

wire n4454;
// (1, 19, 'lutff_0/lout')

wire n4455;
// (1, 19, 'carry_in_mux')

// Carry-In for (1 19)
assign n4455 = 1;

wire n4456;
// (8, 12, 'lutff_7/lout')

wire n4457;
// (10, 21, 'lutff_4/lout')

wire n4458;
// (10, 13, 'lutff_0/lout')

wire n4459;
// (9, 17, 'lutff_3/lout')

wire n4460;
// (13, 21, 'lutff_2/lout')

wire n4461;
// (7, 9, 'lutff_6/lout')

wire n4462;
// (8, 5, 'lutff_4/lout')

wire n4463;
// (21, 23, 'lutff_1/lout')

wire n4464;
// (20, 19, 'lutff_6/lout')

wire n4465;
// (20, 11, 'lutff_2/lout')

wire n4466;
// (10, 14, 'lutff_1/lout')

wire n4467;
// (18, 24, 'lutff_4/lout')

wire n4468;
// (9, 18, 'lutff_4/out')

wire n4469;
// (9, 18, 'lutff_4/lout')

wire n4470;
// (9, 10, 'lutff_0/lout')

wire n4471;
// (16, 8, 'lutff_4/lout')

wire n4472;
// (13, 13, 'lutff_3/lout')

wire n4473;
// (20, 12, 'lutff_3/lout')

wire n4474;
// (3, 19, 'lutff_7/lout')

wire n4475;
// (16, 1, 'lutff_1/lout')

wire n4476;
// (2, 20, 'lutff_3/lout')

wire n4477;
// (10, 9, 'lutff_7/lout')

wire n4478;
// (9, 5, 'lutff_6/lout')

wire n4479;
// (1, 8, 'lutff_4/lout')

wire n4480;
// (3, 11, 'lutff_2/lout')

wire n4481;
// (11, 14, 'lutff_3/lout')

wire n4482;
// (12, 18, 'lutff_5/lout')

wire n4483;
// (12, 10, 'lutff_1/lout')

wire n4484;
// (2, 13, 'lutff_0/lout')

wire n4485;
// (10, 2, 'lutff_4/lout')

wire n4486;
// (9, 6, 'lutff_7/lout')

wire n4487;
// (22, 16, 'lutff_6/lout')

wire n4488;
// (2, 16, 'lutff_5/lout')

wire n4489;
// (13, 9, 'lutff_4/lout')

wire n4490;
// (22, 8, 'lutff_2/lout')

wire n4491;
// (3, 12, 'lutff_3/lout')

wire n4492;
// (21, 12, 'lutff_5/lout')

wire n4493;
// (21, 4, 'lutff_1/lout')

wire n4494;
// (1, 4, 'lutff_6/lout')

wire n4495;
// (15, 18, 'lutff_1/out')

wire n4496;
// (15, 18, 'lutff_1/lout')

wire n4497;
// (12, 14, 'lutff_7/lout')

wire n4498;
// (18, 5, 'lutff_4/lout')

wire n4499;
// (5, 20, 'lutff_4/lout')

wire n4500;
// (2, 9, 'lutff_2/lout')

wire n4501;
// (13, 2, 'lutff_1/lout')

wire n4502;
// (11, 15, 'lutff_3/lout')

wire n4503;
// (14, 23, 'lutff_4/lout')

wire n4504;
// (8, 20, 'lutff_2/lout')

wire n4505;
// (2, 8, 'lutff_6/lout')

wire n4506;
// (13, 1, 'lutff_5/out')

wire n4507;
// (13, 1, 'lutff_5/lout')

wire n4508;
// (18, 6, 'lutff_5/lout')

wire n4509;
// (15, 10, 'lutff_2/lout')

wire n4510;
// (21, 5, 'lutff_1/lout')

wire n4511;
// (15, 13, 'lutff_7/lout')

wire n4512;
// (5, 16, 'lutff_6/lout')

wire n4513;
// (4, 12, 'lutff_5/lout')

wire n4514;
// (14, 15, 'lutff_5/lout')

wire n4515;
// (8, 16, 'lutff_4/lout')

wire n4516;
// (17, 22, 'lutff_5/lout')

wire n4517;
// (23, 13, 'lutff_2/lout')

wire n4518;
// (17, 14, 'lutff_1/lout')

wire n4519;
// (11, 2, 'lutff_5/lout')

wire n4520;
// (7, 17, 'lutff_0/lout')

wire n4521;
// (5, 17, 'lutff_7/lout')

wire n4522;
// (15, 6, 'lutff_4/lout')

wire n4523;
// (2, 1, 'lutff_2/lout')

wire n4524;
// (5, 9, 'lutff_3/lout')

wire n4525;
// (4, 13, 'lutff_6/lout')

wire n4526;
// (4, 5, 'lutff_2/lout')

wire n4527;
// (14, 7, 'lutff_0/lout')

wire n4528;
// (16, 19, 'lutff_4/lout')

wire n4529;
// (17, 15, 'lutff_2/lout')

wire n4530;
// (11, 3, 'lutff_6/lout')

wire n4531;
// (14, 11, 'lutff_7/lout')

wire n4532;
// (15, 7, 'lutff_5/lout')

wire n4533;
// (20, 22, 'lutff_7/lout')

wire n4534;
// (14, 8, 'lutff_1/lout')

wire n4535;
// (9, 20, 'lutff_3/lout')

wire n4536;
// (5, 1, 'lutff_4/lout')

wire n4537;
// (7, 12, 'lutff_6/lout')

wire n4538;
// (8, 8, 'lutff_4/lout')

wire n4539;
// (16, 11, 'lutff_5/lout')

wire n4540;
// (23, 2, 'lutff_1/out')

wire n4541;
// (23, 2, 'lutff_1/lout')

wire n4542;
// (20, 14, 'lutff_2/lout')

wire n4543;
// (10, 17, 'lutff_1/lout')

wire n4544;
// (9, 13, 'lutff_0/lout')

wire n4545;
// (7, 13, 'lutff_7/lout')

wire n4546;
// (17, 2, 'lutff_4/lout')

wire n4547;
// (7, 5, 'lutff_3/lout')

wire n4548;
// (8, 1, 'lutff_1/lout')

wire n4549;
// (9, 16, 'lutff_5/out')

wire n4550;
// (9, 16, 'lutff_5/lout')

wire n4551;
// (1, 19, 'lutff_3/lout')

wire n4552;
// (14, 3, 'lutff_7/lout')

wire n4553;
// (8, 4, 'lutff_6/lout')

wire n4554;
// (16, 7, 'lutff_7/lout')

wire n4555;
// (12, 21, 'lutff_0/out')

wire n4556;
// (12, 21, 'lutff_0/lout')

wire n4557;
// (12, 21, 'carry_in_mux')

// Carry-In for (12 21)
assign n4557 = 1;

wire n4558;
// (17, 3, 'lutff_5/lout')

wire n4559;
// (10, 21, 'lutff_7/lout')

wire n4560;
// (10, 13, 'lutff_3/lout')

wire n4561;
// (9, 17, 'lutff_6/lout')

wire n4562;
// (9, 9, 'lutff_2/lout')

wire n4563;
// (21, 23, 'lutff_4/lout')

wire n4564;
// (1, 3, 'lutff_0/lout')

wire n4565;
// (13, 12, 'lutff_5/lout')

wire n4566;
// (13, 4, 'lutff_1/lout')

wire n4567;
// (18, 16, 'lutff_3/lout')

wire n4568;
// (12, 13, 'lutff_1/lout')

wire n4569;
// (10, 5, 'lutff_4/lout')

wire n4570;
// (9, 1, 'lutff_3/lout')

wire n4571;
// (2, 19, 'lutff_5/lout')

wire n4572;
// (13, 13, 'lutff_6/lout')

wire n4573;
// (22, 11, 'lutff_2/lout')

wire n4574;
// (2, 11, 'lutff_1/lout')

wire n4575;
// (3, 15, 'lutff_3/lout')

wire n4576;
// (22, 19, 'lutff_6/lout')

wire n4577;
// (21, 15, 'lutff_5/lout')

wire n4578;
// (21, 7, 'lutff_1/lout')

wire n4579;
// (1, 7, 'lutff_6/lout')

wire n4580;
// (11, 10, 'lutff_0/lout')

wire n4581;
// (12, 17, 'lutff_7/lout')

wire n4582;
// (18, 8, 'lutff_4/lout')

wire n4583;
// (2, 20, 'lutff_6/lout')

wire n4584;
// (12, 9, 'lutff_3/lout')

wire n4585;
// (2, 12, 'lutff_2/lout')

wire n4586;
// (13, 5, 'lutff_1/lout')

wire n4587;
// (21, 8, 'lutff_2/lout')

wire n4588;
// (14, 18, 'lutff_0/lout')

wire n4589;
// (11, 14, 'lutff_6/lout')

wire n4590;
// (18, 1, 'lutff_1/lout')

wire n4591;
// (8, 18, 'lutff_3/lout')

wire n4592;
// (12, 2, 'lutff_0/lout')

wire n4593;
// (17, 17, 'lutff_2/lout')

wire n4594;
// (12, 1, 'lutff_4/out')

wire n4595;
// (12, 1, 'lutff_4/lout')

wire n4596;
// (5, 19, 'lutff_6/lout')

wire n4597;
// (22, 8, 'lutff_5/lout')

wire n4598;
// (5, 11, 'lutff_2/lout')

wire n4599;
// (21, 4, 'lutff_4/lout')

wire n4600;
// (4, 15, 'lutff_5/lout')

wire n4601;
// (4, 7, 'lutff_1/lout')

wire n4602;
// (8, 19, 'lutff_4/out')

wire n4603;
// (8, 19, 'lutff_4/lout')

wire n4604;
// (14, 10, 'lutff_1/lout')

wire n4605;
// (8, 11, 'lutff_0/lout')

wire n4606;
// (11, 6, 'lutff_7/lout')

wire n4607;
// (7, 20, 'lutff_0/out')

wire n4608;
// (7, 20, 'lutff_0/lout')

wire n4609;
// (7, 20, 'carry_in_mux')

// Carry-In for (7 20)
assign n4609 = 1;

wire n4610;
// (5, 20, 'lutff_7/lout')

wire n4611;
// (15, 9, 'lutff_4/lout')

wire n4612;
// (5, 12, 'lutff_3/lout')

wire n4613;
// (4, 8, 'lutff_2/lout')

wire n4614;
// (16, 14, 'lutff_0/lout')

wire n4615;
// (17, 18, 'lutff_2/lout')

wire n4616;
// (14, 14, 'lutff_7/lout')

wire n4617;
// (15, 10, 'lutff_5/lout')

wire n4618;
// (14, 6, 'lutff_3/lout')

wire n4619;
// (15, 2, 'lutff_1/lout')

wire n4620;
// (1, 21, 'lutff_3/lout')

wire n4621;
// (5, 5, 'lutff_0/lout')

wire n4622;
// (7, 16, 'lutff_2/lout')

wire n4623;
// (16, 15, 'lutff_1/lout')

wire n4624;
// (9, 19, 'lutff_6/lout')

wire n4625;
// (1, 14, 'lutff_0/lout')

wire n4626;
// (10, 20, 'lutff_1/lout')

wire n4627;
// (8, 7, 'lutff_7/lout')

wire n4628;
// (17, 5, 'lutff_4/lout')

wire n4629;
// (20, 13, 'lutff_5/lout')

wire n4630;
// (7, 8, 'lutff_3/lout')

wire n4631;
// (13, 23, 'lutff_4/lout')

wire n4632;
// (16, 10, 'lutff_7/lout')

wire n4633;
// (17, 6, 'lutff_5/lout')

wire n4634;
// (16, 2, 'lutff_3/lout')

wire n4635;
// (10, 16, 'lutff_3/lout')

wire n4636;
// (9, 20, 'lutff_6/lout')

wire n4637;
// (5, 1, 'lutff_7/lout')

wire n4638;
// (9, 12, 'lutff_2/lout')

wire n4639;
// (7, 4, 'lutff_5/lout')

wire n4640;
// (13, 15, 'lutff_5/lout')

wire n4641;
// (20, 14, 'lutff_5/lout')

wire n4642;
// (20, 6, 'lutff_1/lout')

wire n4643;
// (10, 9, 'lutff_0/lout')

wire n4644;
// (1, 10, 'lutff_7/lout')

wire n4645;
// (17, 2, 'lutff_7/lout')

wire n4646;
// (1, 2, 'lutff_3/lout')

wire n4647;
// (10, 8, 'lutff_4/lout')

wire n4648;
// (9, 4, 'lutff_3/lout')

wire n4649;
// (2, 14, 'lutff_1/lout')

wire n4650;
// (13, 8, 'lutff_2/lout')

wire n4651;
// (18, 12, 'lutff_0/lout')

wire n4652;
// (13, 11, 'lutff_7/lout')

wire n4653;
// (11, 16, 'lutff_5/lout')

wire n4654;
// (10, 1, 'lutff_1/lout')

wire n4655;
// (12, 12, 'lutff_3/lout')

wire n4656;
// (22, 15, 'lutff_3/lout')

wire n4657;
// (2, 15, 'lutff_2/lout')

wire n4658;
// (10, 4, 'lutff_6/lout')

wire n4659;
// (1, 3, 'lutff_3/lout')

wire n4660;
// (2, 18, 'lutff_7/lout')

wire n4661;
// (14, 21, 'lutff_0/lout')

wire n4662;
// (13, 4, 'lutff_4/lout')

wire n4663;
// (21, 14, 'lutff_7/lout')

wire n4664;
// (11, 17, 'lutff_6/lout')

wire n4665;
// (11, 9, 'lutff_2/lout')

wire n4666;
// (12, 13, 'lutff_4/lout')

wire n4667;
// (12, 5, 'lutff_0/lout')

wire n4668;
// (3, 6, 'lutff_7/lout')

wire n4669;
// (10, 5, 'lutff_7/lout')

wire n4670;
// (4, 19, 'lutff_1/lout')

wire n4671;
// (9, 1, 'lutff_6/lout')

wire n4672;
// (14, 22, 'lutff_1/lout')

wire n4673;
// (2, 11, 'lutff_4/lout')

wire n4674;
// (4, 18, 'lutff_5/out')

wire n4675;
// (4, 18, 'lutff_5/lout')

wire n4676;
// (21, 7, 'lutff_4/lout')

wire n4677;
// (8, 14, 'lutff_0/lout')

wire n4678;
// (18, 8, 'lutff_7/lout')

wire n4679;
// (5, 15, 'lutff_3/lout')

wire n4680;
// (17, 16, 'lutff_4/lout')

wire n4681;
// (4, 11, 'lutff_2/lout')

wire n4682;
// (8, 15, 'lutff_1/out')

wire n4683;
// (8, 15, 'lutff_1/lout')

wire n4684;
// (2, 3, 'lutff_5/lout')

wire n4685;
// (22, 3, 'lutff_6/lout')

wire n4686;
// (4, 14, 'lutff_7/lout')

wire n4687;
// (16, 17, 'lutff_0/lout')

wire n4688;
// (8, 18, 'lutff_6/lout')

wire n4689;
// (14, 9, 'lutff_3/lout')

wire n4690;
// (15, 5, 'lutff_1/lout')

wire n4691;
// (5, 8, 'lutff_0/lout')

wire n4692;
// (17, 17, 'lutff_5/lout')

wire n4693;
// (12, 1, 'lutff_7/out')

wire n4694;
// (12, 1, 'lutff_7/lout')

wire n4695;
// (16, 18, 'lutff_1/lout')

wire n4696;
// (4, 7, 'lutff_4/lout')

wire n4697;
// (14, 10, 'lutff_4/lout')

wire n4698;
// (14, 2, 'lutff_0/lout')

wire n4699;
// (16, 21, 'lutff_6/lout')

wire n4700;
// (1, 17, 'lutff_0/out')

wire n4701;
// (1, 17, 'lutff_0/lout')

wire n4702;
// (1, 17, 'carry_in_mux')

// Carry-In for (1 17)
assign n4702 = 1;

wire n4703;
// (23, 8, 'lutff_1/lout')

wire n4704;
// (17, 9, 'lutff_0/lout')

wire n4705;
// (8, 10, 'lutff_7/lout')

wire n4706;
// (8, 2, 'lutff_3/lout')

wire n4707;
// (1, 20, 'lutff_5/lout')

wire n4708;
// (10, 19, 'lutff_4/lout')

wire n4709;
// (10, 11, 'lutff_0/lout')

wire n4710;
// (5, 3, 'lutff_6/lout')

wire n4711;
// (9, 15, 'lutff_3/lout')

wire n4712;
// (17, 4, 'lutff_7/lout')

wire n4713;
// (13, 18, 'lutff_0/lout')

wire n4714;
// (8, 3, 'lutff_4/lout')

wire n4715;
// (1, 21, 'lutff_6/lout')

wire n4716;
// (16, 13, 'lutff_7/lout')

wire n4717;
// (16, 5, 'lutff_3/lout')

wire n4718;
// (1, 13, 'lutff_2/lout')

wire n4719;
// (17, 1, 'lutff_1/lout')

wire n4720;
// (20, 9, 'lutff_2/lout')

wire n4721;
// (18, 22, 'lutff_4/lout')

wire n4722;
// (18, 14, 'lutff_0/lout')

wire n4723;
// (13, 19, 'lutff_1/lout')

wire n4724;
// (7, 7, 'lutff_5/lout')

wire n4725;
// (21, 21, 'lutff_0/lout')

wire n4726;
// (16, 6, 'lutff_4/lout')

wire n4727;
// (10, 12, 'lutff_0/lout')

wire n4728;
// (3, 13, 'lutff_0/out')

wire n4729;
// (3, 13, 'lutff_0/lout')

wire n4730;
// (3, 13, 'carry_in_mux')

// Carry-In for (3 13)
assign n4730 = 1;

wire n4731;
// (17, 5, 'lutff_7/lout')

wire n4732;
// (1, 5, 'lutff_3/lout')

wire n4733;
// (3, 16, 'lutff_5/lout')

wire n4734;
// (18, 18, 'lutff_6/lout')

wire n4735;
// (12, 15, 'lutff_4/lout')

wire n4736;
// (10, 7, 'lutff_7/lout')

wire n4737;
// (4, 21, 'lutff_1/out')

wire n4738;
// (4, 21, 'lutff_1/lout')

wire n4739;
// (16, 2, 'lutff_6/lout')

wire n4740;
// (13, 14, 'lutff_7/lout')

wire n4741;
// (3, 17, 'lutff_6/lout')

wire n4742;
// (3, 9, 'lutff_2/lout')

wire n4743;
// (18, 10, 'lutff_7/lout')

wire n4744;
// (9, 3, 'lutff_5/lout')

wire n4745;
// (12, 11, 'lutff_6/lout')

wire n4746;
// (13, 7, 'lutff_4/lout')

wire n4747;
// (21, 17, 'lutff_7/lout')

wire n4748;
// (11, 20, 'lutff_6/lout')

wire n4749;
// (1, 2, 'lutff_6/lout')

wire n4750;
// (12, 8, 'lutff_0/lout')

wire n4751;
// (15, 16, 'lutff_1/out')

wire n4752;
// (15, 16, 'lutff_1/lout')

wire n4753;
// (10, 8, 'lutff_7/lout')

wire n4754;
// (9, 4, 'lutff_6/lout')

wire n4755;
// (22, 14, 'lutff_5/out')

wire n4756;
// (22, 14, 'lutff_5/lout')

wire n4757;
// (2, 14, 'lutff_4/lout')

wire n4758;
// (22, 6, 'lutff_1/lout')

wire n4759;
// (11, 13, 'lutff_3/lout')

wire n4760;
// (21, 2, 'lutff_0/lout')

wire n4761;
// (8, 17, 'lutff_0/out')

wire n4762;
// (8, 17, 'lutff_0/lout')

wire n4763;
// (8, 17, 'carry_in_mux')

// Carry-In for (8 17)
assign n4763 = 1;

wire n4764;
// (23, 19, 'lutff_1/lout')

wire n4765;
// (12, 4, 'lutff_2/lout')

wire n4766;
// (15, 8, 'lutff_2/lout')

wire n4767;
// (22, 7, 'lutff_2/lout')

wire n4768;
// (17, 19, 'lutff_4/lout')

wire n4769;
// (15, 11, 'lutff_7/lout')

wire n4770;
// (2, 6, 'lutff_5/lout')

wire n4771;
// (5, 14, 'lutff_6/lout')

wire n4772;
// (8, 21, 'lutff_6/lout')

wire n4773;
// (14, 12, 'lutff_3/lout')

wire n4774;
// (17, 20, 'lutff_5/lout')

wire n4775;
// (17, 12, 'lutff_1/lout')

wire n4776;
// (15, 4, 'lutff_4/lout')

wire n4777;
// (23, 14, 'lutff_7/lout')

wire n4778;
// (5, 6, 'lutff_1/lout')

wire n4779;
// (14, 13, 'lutff_4/lout')

wire n4780;
// (4, 2, 'lutff_0/lout')

wire n4781;
// (8, 14, 'lutff_3/lout')

wire n4782;
// (2, 2, 'lutff_7/lout')

wire n4783;
// (14, 5, 'lutff_0/lout')

wire n4784;
// (16, 16, 'lutff_2/lout')

wire n4785;
// (13, 21, 'lutff_1/lout')

wire n4786;
// (8, 13, 'lutff_7/lout')

wire n4787;
// (11, 1, 'lutff_6/out')

wire n4788;
// (11, 1, 'lutff_6/lout')

wire n4789;
// (5, 7, 'lutff_2/lout')

wire n4790;
// (4, 3, 'lutff_1/lout')

wire n4791;
// (9, 18, 'lutff_3/out')

wire n4792;
// (9, 18, 'lutff_3/lout')

wire n4793;
// (16, 17, 'lutff_3/lout')

wire n4794;
// (7, 2, 'lutff_2/lout')

wire n4795;
// (8, 6, 'lutff_4/lout')

wire n4796;
// (1, 16, 'lutff_2/lout')

wire n4797;
// (20, 20, 'lutff_6/lout')

wire n4798;
// (10, 15, 'lutff_1/lout')

wire n4799;
// (13, 22, 'lutff_1/lout')

wire n4800;
// (10, 18, 'lutff_6/out')

wire n4801;
// (10, 18, 'lutff_6/lout')

wire n4802;
// (9, 14, 'lutff_5/lout')

wire n4803;
// (8, 2, 'lutff_6/lout')

wire n4804;
// (16, 4, 'lutff_5/lout')

wire n4805;
// (12, 19, 'lutff_0/lout')

wire n4806;
// (7, 3, 'lutff_2/lout')

wire n4807;
// (10, 11, 'lutff_3/lout')

wire n4808;
// (16, 5, 'lutff_6/lout')

wire n4809;
// (2, 16, 'lutff_4/lout')

wire n4810;
// (3, 20, 'lutff_6/lout')

wire n4811;
// (13, 9, 'lutff_3/lout')

wire n4812;
// (3, 12, 'lutff_2/lout')

wire n4813;
// (18, 14, 'lutff_3/lout')

wire n4814;
// (1, 4, 'lutff_5/lout')

wire n4815;
// (15, 18, 'lutff_0/out')

wire n4816;
// (15, 18, 'lutff_0/lout')

wire n4817;
// (15, 18, 'carry_in_mux')

// Carry-In for (15 18)
assign n4817 = 1;

wire n4818;
// (12, 14, 'lutff_6/lout')

wire n4819;
// (22, 17, 'lutff_6/lout')

wire n4820;
// (2, 17, 'lutff_5/lout')

wire n4821;
// (13, 10, 'lutff_4/lout')

wire n4822;
// (2, 9, 'lutff_1/lout')

wire n4823;
// (3, 13, 'lutff_3/out')

wire n4824;
// (3, 13, 'lutff_3/lout')

wire n4825;
// (13, 2, 'lutff_0/lout')

wire n4826;
// (11, 15, 'lutff_2/lout')

wire n4827;
// (1, 5, 'lutff_6/lout')

wire n4828;
// (14, 23, 'lutff_3/lout')

wire n4829;
// (15, 19, 'lutff_1/out')

wire n4830;
// (15, 19, 'lutff_1/lout')

wire n4831;
// (10, 3, 'lutff_3/lout')

wire n4832;
// (12, 15, 'lutff_7/lout')

wire n4833;
// (18, 6, 'lutff_4/lout')

wire n4834;
// (12, 7, 'lutff_3/lout')

wire n4835;
// (13, 3, 'lutff_1/lout')

wire n4836;
// (21, 13, 'lutff_4/lout')

wire n4837;
// (4, 21, 'lutff_4/out')

wire n4838;
// (4, 21, 'lutff_4/lout')

wire n4839;
// (21, 5, 'lutff_0/lout')

wire n4840;
// (8, 16, 'lutff_3/lout')

wire n4841;
// (21, 6, 'lutff_1/lout')

wire n4842;
// (18, 2, 'lutff_6/lout')

wire n4843;
// (15, 14, 'lutff_7/lout')

wire n4844;
// (5, 9, 'lutff_2/lout')

wire n4845;
// (4, 13, 'lutff_5/lout')

wire n4846;
// (11, 4, 'lutff_1/lout')

wire n4847;
// (4, 5, 'lutff_1/lout')

wire n4848;
// (3, 1, 'lutff_6/lout')

wire n4849;
// (16, 19, 'lutff_3/out')

wire n4850;
// (16, 19, 'lutff_3/lout')

wire n4851;
// (17, 15, 'lutff_1/lout')

wire n4852;
// (11, 3, 'lutff_5/lout')

wire n4853;
// (14, 11, 'lutff_6/lout')

wire n4854;
// (7, 18, 'lutff_0/out')

wire n4855;
// (7, 18, 'lutff_0/lout')

wire n4856;
// (7, 18, 'carry_in_mux')

// Carry-In for (7 18)
assign n4856 = 1;

wire n4857;
// (15, 7, 'lutff_4/lout')

wire n4858;
// (23, 17, 'lutff_7/lout')

wire n4859;
// (5, 10, 'lutff_3/lout')

wire n4860;
// (7, 21, 'lutff_5/lout')

wire n4861;
// (8, 17, 'lutff_3/out')

wire n4862;
// (8, 17, 'lutff_3/lout')

wire n4863;
// (14, 8, 'lutff_0/lout')

wire n4864;
// (4, 9, 'lutff_7/lout')

wire n4865;
// (15, 8, 'lutff_5/lout')

wire n4866;
// (17, 19, 'lutff_7/out')

wire n4867;
// (17, 19, 'lutff_7/lout')

wire n4868;
// (17, 11, 'lutff_3/lout')

wire n4869;
// (23, 2, 'lutff_0/out')

wire n4870;
// (23, 2, 'lutff_0/lout')

wire n4871;
// (23, 2, 'carry_in_mux')

// Carry-In for (23 2)
assign n4871 = 1;

wire n4872;
// (4, 6, 'lutff_1/lout')

wire n4873;
// (7, 14, 'lutff_2/lout')

wire n4874;
// (16, 20, 'lutff_3/lout')

wire n4875;
// (7, 13, 'lutff_6/lout')

wire n4876;
// (14, 12, 'lutff_6/lout')

wire n4877;
// (14, 4, 'lutff_2/lout')

wire n4878;
// (8, 1, 'lutff_0/lout')

wire n4879;
// (1, 19, 'lutff_2/lout')

wire n4880;
// (23, 3, 'lutff_1/out')

wire n4881;
// (23, 3, 'lutff_1/lout')

wire n4882;
// (8, 4, 'lutff_5/lout')

wire n4883;
// (20, 18, 'lutff_7/lout')

wire n4884;
// (17, 3, 'lutff_4/lout')

wire n4885;
// (10, 13, 'lutff_2/lout')

wire n4886;
// (9, 17, 'lutff_5/lout')

wire n4887;
// (9, 9, 'lutff_1/lout')

wire n4888;
// (13, 21, 'lutff_4/lout')

wire n4889;
// (8, 5, 'lutff_6/lout')

wire n4890;
// (12, 22, 'lutff_0/out')

wire n4891;
// (12, 22, 'lutff_0/lout')

wire n4892;
// (12, 22, 'carry_in_mux')

// Carry-In for (12 22)
assign n4892 = 1;

wire n4893;
// (20, 11, 'lutff_4/lout')

wire n4894;
// (10, 14, 'lutff_3/lout')

wire n4895;
// (9, 18, 'lutff_6/out')

wire n4896;
// (9, 18, 'lutff_6/lout')

wire n4897;
// (9, 10, 'lutff_2/lout')

wire n4898;
// (22, 20, 'lutff_1/lout')

wire n4899;
// (7, 2, 'lutff_5/lout')

wire n4900;
// (21, 16, 'lutff_0/lout')

wire n4901;
// (16, 8, 'lutff_6/lout')

wire n4902;
// (13, 13, 'lutff_5/lout')

wire n4903;
// (3, 15, 'lutff_2/lout')

wire n4904;
// (20, 4, 'lutff_1/lout')

wire n4905;
// (18, 17, 'lutff_3/lout')

wire n4906;
// (1, 7, 'lutff_5/lout')

wire n4907;
// (12, 17, 'lutff_6/lout')

wire n4908;
// (2, 20, 'lutff_5/lout')

wire n4909;
// (22, 12, 'lutff_2/lout')

wire n4910;
// (2, 12, 'lutff_1/lout')

wire n4911;
// (13, 5, 'lutff_0/lout')

wire n4912;
// (21, 8, 'lutff_1/out')

wire n4913;
// (21, 8, 'lutff_1/lout')

wire n4914;
// (1, 8, 'lutff_6/lout')

wire n4915;
// (11, 14, 'lutff_5/lout')

wire n4916;
// (12, 18, 'lutff_7/lout')

wire n4917;
// (2, 13, 'lutff_2/lout')

wire n4918;
// (13, 6, 'lutff_1/lout')

wire n4919;
// (10, 2, 'lutff_6/lout')

wire n4920;
// (4, 16, 'lutff_0/lout')

wire n4921;
// (2, 16, 'lutff_7/lout')

wire n4922;
// (13, 9, 'lutff_6/lout')

wire n4923;
// (14, 19, 'lutff_0/out')

wire n4924;
// (14, 19, 'lutff_0/lout')

wire n4925;
// (14, 19, 'carry_in_mux')

// Carry-In for (14 19)
assign n4925 = 0;

wire n4926;
// (3, 12, 'lutff_5/lout')

wire n4927;
// (21, 12, 'lutff_7/lout')

wire n4928;
// (22, 8, 'lutff_4/lout')

wire n4929;
// (3, 4, 'lutff_1/lout')

wire n4930;
// (21, 4, 'lutff_3/lout')

wire n4931;
// (15, 18, 'lutff_3/out')

wire n4932;
// (15, 18, 'lutff_3/lout')

wire n4933;
// (8, 19, 'lutff_3/out')

wire n4934;
// (8, 19, 'lutff_3/lout')

wire n4935;
// (12, 3, 'lutff_0/out')

wire n4936;
// (12, 3, 'lutff_0/lout')

wire n4937;
// (12, 3, 'carry_in_mux')

// Carry-In for (12 3)
assign n4937 = 1;

wire n4938;
// (18, 5, 'lutff_6/lout')

wire n4939;
// (5, 20, 'lutff_6/lout')

wire n4940;
// (17, 21, 'lutff_7/lout')

wire n4941;
// (11, 15, 'lutff_5/lout')

wire n4942;
// (11, 7, 'lutff_1/lout')

wire n4943;
// (8, 20, 'lutff_4/lout')

wire n4944;
// (13, 1, 'lutff_7/out')

wire n4945;
// (13, 1, 'lutff_7/lout')

wire n4946;
// (17, 18, 'lutff_1/lout')

wire n4947;
// (14, 14, 'lutff_6/lout')

wire n4948;
// (15, 10, 'lutff_4/lout')

wire n4949;
// (15, 2, 'lutff_0/lout')

wire n4950;
// (7, 16, 'lutff_1/lout')

wire n4951;
// (16, 15, 'lutff_0/lout')

wire n4952;
// (14, 15, 'lutff_7/lout')

wire n4953;
// (8, 16, 'lutff_6/lout')

wire n4954;
// (15, 3, 'lutff_1/lout')

wire n4955;
// (17, 14, 'lutff_3/lout')

wire n4956;
// (7, 17, 'lutff_2/lout')

wire n4957;
// (15, 6, 'lutff_6/lout')

wire n4958;
// (2, 1, 'lutff_4/lout')

wire n4959;
// (5, 9, 'lutff_5/lout')

wire n4960;
// (4, 5, 'lutff_4/lout')

wire n4961;
// (14, 7, 'lutff_2/lout')

wire n4962;
// (16, 19, 'lutff_6/lout')

wire n4963;
// (13, 23, 'lutff_3/lout')

wire n4964;
// (17, 7, 'lutff_0/out')

wire n4965;
// (17, 7, 'lutff_0/lout')

wire n4966;
// (1, 18, 'lutff_5/lout')

wire n4967;
// (17, 6, 'lutff_4/out')

wire n4968;
// (17, 6, 'lutff_4/lout')

wire n4969;
// (10, 16, 'lutff_2/lout')

wire n4970;
// (9, 20, 'lutff_5/lout')

wire n4971;
// (9, 12, 'lutff_1/lout')

wire n4972;
// (13, 16, 'lutff_0/lout')

wire n4973;
// (7, 4, 'lutff_4/lout')

wire n4974;
// (8, 8, 'lutff_6/lout')

wire n4975;
// (16, 11, 'lutff_7/lout')

wire n4976;
// (23, 2, 'lutff_3/lout')

wire n4977;
// (16, 3, 'lutff_3/lout')

wire n4978;
// (20, 14, 'lutff_4/lout')

wire n4979;
// (20, 6, 'lutff_0/out')

wire n4980;
// (20, 6, 'lutff_0/lout')

wire n4981;
// (20, 6, 'carry_in_mux')

// Carry-In for (20 6)
assign n4981 = 1;

wire n4982;
// (9, 13, 'lutff_2/lout')

wire n4983;
// (17, 2, 'lutff_6/lout')

wire n4984;
// (22, 23, 'lutff_1/lout')

wire n4985;
// (13, 17, 'lutff_1/out')

wire n4986;
// (13, 17, 'lutff_1/lout')

wire n4987;
// (7, 5, 'lutff_5/lout')

wire n4988;
// (8, 1, 'lutff_3/lout')

wire n4989;
// (9, 16, 'lutff_7/out')

wire n4990;
// (9, 16, 'lutff_7/lout')

wire n4991;
// (20, 15, 'lutff_5/lout')

wire n4992;
// (20, 7, 'lutff_1/out')

wire n4993;
// (20, 7, 'lutff_1/lout')

wire n4994;
// (10, 10, 'lutff_0/lout')

wire n4995;
// (18, 20, 'lutff_3/lout')

wire n4996;
// (12, 21, 'lutff_2/lout')

wire n4997;
// (17, 3, 'lutff_7/lout')

wire n4998;
// (3, 14, 'lutff_5/lout')

wire n4999;
// (10, 13, 'lutff_5/lout')

wire n5000;
// (9, 9, 'lutff_4/lout')

wire n5001;
// (2, 15, 'lutff_1/lout')

wire n5002;
// (18, 13, 'lutff_0/lout')

wire n5003;
// (1, 3, 'lutff_2/lout')

wire n5004;
// (13, 12, 'lutff_7/lout')

wire n5005;
// (2, 18, 'lutff_6/lout')

wire n5006;
// (13, 4, 'lutff_3/lout')

wire n5007;
// (11, 17, 'lutff_5/lout')

wire n5008;
// (18, 16, 'lutff_5/lout')

wire n5009;
// (12, 13, 'lutff_3/lout')

wire n5010;
// (4, 19, 'lutff_0/lout')

wire n5011;
// (9, 1, 'lutff_5/lout')

wire n5012;
// (2, 19, 'lutff_7/lout')

wire n5013;
// (14, 22, 'lutff_0/lout')

wire n5014;
// (22, 11, 'lutff_4/lout')

wire n5015;
// (2, 11, 'lutff_3/lout')

wire n5016;
// (3, 15, 'lutff_5/lout')

wire n5017;
// (3, 7, 'lutff_1/lout')

wire n5018;
// (11, 18, 'lutff_6/lout')

wire n5019;
// (21, 7, 'lutff_3/out')

wire n5020;
// (21, 7, 'lutff_3/lout')

wire n5021;
// (11, 10, 'lutff_2/lout')

wire n5022;
// (12, 6, 'lutff_0/lout')

wire n5023;
// (24, 20, 'lutff_2/lout')

wire n5024;
// (4, 20, 'lutff_1/lout')

wire n5025;
// (18, 8, 'lutff_6/lout')

wire n5026;
// (12, 9, 'lutff_5/lout')

wire n5027;
// (2, 12, 'lutff_4/lout')

wire n5028;
// (13, 5, 'lutff_3/lout')

wire n5029;
// (22, 4, 'lutff_1/lout')

wire n5030;
// (2, 4, 'lutff_0/lout')

wire n5031;
// (21, 8, 'lutff_4/lout')

wire n5032;
// (14, 18, 'lutff_2/lout')

wire n5033;
// (8, 15, 'lutff_0/out')

wire n5034;
// (8, 15, 'lutff_0/lout')

wire n5035;
// (8, 15, 'carry_in_mux')

// Carry-In for (8 15)
assign n5035 = 1;

wire n5036;
// (18, 1, 'lutff_3/lout')

wire n5037;
// (8, 18, 'lutff_5/lout')

wire n5038;
// (17, 17, 'lutff_4/lout')

wire n5039;
// (7, 19, 'lutff_1/lout')

wire n5040;
// (12, 1, 'lutff_6/out')

wire n5041;
// (12, 1, 'lutff_6/lout')

wire n5042;
// (5, 11, 'lutff_4/lout')

wire n5043;
// (4, 15, 'lutff_7/lout')

wire n5044;
// (16, 18, 'lutff_0/out')

wire n5045;
// (16, 18, 'lutff_0/lout')

wire n5046;
// (16, 18, 'carry_in_mux')

// Carry-In for (16 18)
assign n5046 = 1;

wire n5047;
// (23, 17, 'lutff_0/lout')

wire n5048;
// (4, 7, 'lutff_3/lout')

wire n5049;
// (8, 19, 'lutff_6/out')

wire n5050;
// (8, 19, 'lutff_6/lout')

wire n5051;
// (14, 10, 'lutff_3/lout')

wire n5052;
// (8, 11, 'lutff_2/lout')

wire n5053;
// (7, 20, 'lutff_2/out')

wire n5054;
// (7, 20, 'lutff_2/lout')

wire n5055;
// (15, 9, 'lutff_6/lout')

wire n5056;
// (5, 12, 'lutff_5/lout')

wire n5057;
// (5, 4, 'lutff_1/lout')

wire n5058;
// (4, 8, 'lutff_4/lout')

wire n5059;
// (16, 22, 'lutff_6/lout')

wire n5060;
// (16, 14, 'lutff_2/lout')

wire n5061;
// (17, 18, 'lutff_4/lout')

wire n5062;
// (17, 10, 'lutff_0/out')

wire n5063;
// (17, 10, 'lutff_0/lout')

wire n5064;
// (17, 10, 'carry_in_mux')

// Carry-In for (17 10)
assign n5064 = 1;

wire n5065;
// (14, 6, 'lutff_5/lout')

wire n5066;
// (8, 3, 'lutff_3/lout')

wire n5067;
// (1, 21, 'lutff_5/lout')

wire n5068;
// (15, 2, 'lutff_3/lout')

wire n5069;
// (1, 13, 'lutff_1/lout')

wire n5070;
// (20, 17, 'lutff_5/lout')

wire n5071;
// (13, 19, 'lutff_0/out')

wire n5072;
// (13, 19, 'lutff_0/lout')

wire n5073;
// (13, 19, 'carry_in_mux')

// Carry-In for (13 19)
assign n5073 = 1;

wire n5074;
// (23, 13, 'lutff_7/lout')

wire n5075;
// (16, 6, 'lutff_3/lout')

wire n5076;
// (17, 5, 'lutff_6/lout')

wire n5077;
// (20, 13, 'lutff_7/lout')

wire n5078;
// (13, 20, 'lutff_1/out')

wire n5079;
// (13, 20, 'lutff_1/lout')

wire n5080;
// (7, 8, 'lutff_5/lout')

wire n5081;
// (13, 23, 'lutff_6/lout')

wire n5082;
// (20, 10, 'lutff_1/lout')

wire n5083;
// (3, 18, 'lutff_1/lout')

wire n5084;
// (17, 6, 'lutff_7/lout')

wire n5085;
// (16, 2, 'lutff_5/lout')

wire n5086;
// (7, 1, 'lutff_2/lout')

wire n5087;
// (9, 12, 'lutff_4/lout')

wire n5088;
// (7, 4, 'lutff_7/lout')

wire n5089;
// (4, 22, 'lutff_1/lout')

wire n5090;
// (16, 3, 'lutff_6/lout')

wire n5091;
// (11, 21, 'lutff_1/lout')

wire n5092;
// (13, 15, 'lutff_7/lout')

wire n5093;
// (13, 7, 'lutff_3/lout')

wire n5094;
// (20, 6, 'lutff_3/lout')

wire n5095;
// (18, 11, 'lutff_1/lout')

wire n5096;
// (15, 16, 'lutff_0/out')

wire n5097;
// (15, 16, 'lutff_0/lout')

wire n5098;
// (15, 16, 'carry_in_mux')

// Carry-In for (15 16)
assign n5098 = 1;

wire n5099;
// (10, 8, 'lutff_6/lout')

wire n5100;
// (9, 4, 'lutff_5/lout')

wire n5101;
// (22, 14, 'lutff_4/lout')

wire n5102;
// (2, 14, 'lutff_3/lout')

wire n5103;
// (13, 8, 'lutff_4/lout')

wire n5104;
// (10, 1, 'lutff_3/lout')

wire n5105;
// (11, 16, 'lutff_7/lout')

wire n5106;
// (12, 12, 'lutff_5/lout')

wire n5107;
// (18, 3, 'lutff_2/lout')

wire n5108;
// (22, 15, 'lutff_5/lout')

wire n5109;
// (2, 15, 'lutff_4/lout')

wire n5110;
// (12, 4, 'lutff_1/lout')

wire n5111;
// (22, 7, 'lutff_1/lout')

wire n5112;
// (2, 7, 'lutff_0/lout')

wire n5113;
// (21, 11, 'lutff_4/lout')

wire n5114;
// (24, 18, 'lutff_3/lout')

wire n5115;
// (21, 3, 'lutff_0/out')

wire n5116;
// (21, 3, 'lutff_0/lout')

wire n5117;
// (21, 3, 'carry_in_mux')

// Carry-In for (21 3)
assign n5117 = 1;

wire n5118;
// (15, 17, 'lutff_0/lout')

wire n5119;
// (13, 4, 'lutff_6/lout')

wire n5120;
// (17, 21, 'lutff_0/lout')

wire n5121;
// (11, 9, 'lutff_4/lout')

wire n5122;
// (8, 21, 'lutff_5/lout')

wire n5123;
// (12, 5, 'lutff_2/lout')

wire n5124;
// (17, 20, 'lutff_4/lout')

wire n5125;
// (15, 12, 'lutff_7/lout')

wire n5126;
// (4, 18, 'lutff_7/out')

wire n5127;
// (4, 18, 'lutff_7/lout')

wire n5128;
// (21, 7, 'lutff_6/lout')

wire n5129;
// (4, 10, 'lutff_3/lout')

wire n5130;
// (14, 13, 'lutff_3/lout')

wire n5131;
// (8, 14, 'lutff_2/lout')

wire n5132;
// (2, 2, 'lutff_6/lout')

wire n5133;
// (11, 1, 'lutff_5/out')

wire n5134;
// (11, 1, 'lutff_5/lout')

wire n5135;
// (5, 15, 'lutff_5/lout')

wire n5136;
// (5, 7, 'lutff_1/lout')

wire n5137;
// (17, 16, 'lutff_6/lout')

wire n5138;
// (4, 11, 'lutff_4/lout')

wire n5139;
// (4, 3, 'lutff_0/lout')

wire n5140;
// (8, 15, 'lutff_3/out')

wire n5141;
// (8, 15, 'lutff_3/lout')

wire n5142;
// (2, 3, 'lutff_7/lout')

wire n5143;
// (17, 13, 'lutff_0/out')

wire n5144;
// (17, 13, 'lutff_0/lout')

wire n5145;
// (17, 13, 'carry_in_mux')

// Carry-In for (17 13)
assign n5145 = 1;

wire n5146;
// (14, 9, 'lutff_5/lout')

wire n5147;
// (15, 5, 'lutff_3/lout')

wire n5148;
// (5, 8, 'lutff_2/lout')

wire n5149;
// (17, 17, 'lutff_7/lout')

wire n5150;
// (7, 19, 'lutff_4/lout')

wire n5151;
// (4, 4, 'lutff_1/lout')

wire n5152;
// (7, 11, 'lutff_0/lout')

wire n5153;
// (5, 11, 'lutff_7/lout')

wire n5154;
// (16, 18, 'lutff_3/out')

wire n5155;
// (16, 18, 'lutff_3/lout')

wire n5156;
// (4, 7, 'lutff_6/lout')

wire n5157;
// (13, 22, 'lutff_0/lout')

wire n5158;
// (14, 10, 'lutff_6/lout')

wire n5159;
// (14, 2, 'lutff_2/lout')

wire n5160;
// (1, 17, 'lutff_2/lout')

wire n5161;
// (17, 9, 'lutff_2/lout')

wire n5162;
// (8, 2, 'lutff_5/lout')

wire n5163;
// (1, 20, 'lutff_7/lout')

wire n5164;
// (7, 3, 'lutff_1/lout')

wire n5165;
// (10, 11, 'lutff_2/lout')

wire n5166;
// (9, 15, 'lutff_5/lout')

wire n5167;
// (13, 18, 'lutff_2/lout')

wire n5168;
// (3, 21, 'lutff_1/lout')

wire n5169;
// (8, 3, 'lutff_6/lout')

wire n5170;
// (1, 13, 'lutff_4/lout')

wire n5171;
// (17, 1, 'lutff_3/lout')

wire n5172;
// (20, 9, 'lutff_4/lout')

wire n5173;
// (18, 14, 'lutff_2/lout')

wire n5174;
// (9, 7, 'lutff_0/lout')

wire n5175;
// (7, 7, 'lutff_7/lout')

wire n5176;
// (21, 21, 'lutff_2/lout')

wire n5177;
// (16, 6, 'lutff_6/lout')

wire n5178;
// (3, 13, 'lutff_2/out')

wire n5179;
// (3, 13, 'lutff_2/lout')

wire n5180;
// (10, 12, 'lutff_2/lout')

wire n5181;
// (1, 5, 'lutff_5/lout')

wire n5182;
// (15, 19, 'lutff_0/lout')

wire n5183;
// (3, 16, 'lutff_7/lout')

wire n5184;
// (21, 22, 'lutff_3/lout')

wire n5185;
// (22, 18, 'lutff_0/lout')

wire n5186;
// (12, 15, 'lutff_6/lout')

wire n5187;
// (12, 7, 'lutff_2/lout')

wire n5188;
// (13, 3, 'lutff_0/lout')

wire n5189;
// (4, 21, 'lutff_3/lout')

wire n5190;
// (18, 15, 'lutff_2/lout')

wire n5191;
// (22, 13, 'lutff_7/lout')

wire n5192;
// (3, 9, 'lutff_4/lout')

wire n5193;
// (11, 19, 'lutff_7/lout')

wire n5194;
// (2, 10, 'lutff_0/lout')

wire n5195;
// (5, 18, 'lutff_1/lout')

wire n5196;
// (9, 3, 'lutff_7/lout')

wire n5197;
// (21, 6, 'lutff_0/lout')

wire n5198;
// (18, 2, 'lutff_5/lout')

wire n5199;
// (13, 7, 'lutff_6/lout')

wire n5200;
// (3, 2, 'lutff_1/lout')

wire n5201;
// (11, 12, 'lutff_4/lout')

wire n5202;
// (12, 8, 'lutff_2/lout')

wire n5203;
// (11, 4, 'lutff_0/lout')

wire n5204;
// (15, 16, 'lutff_3/lout')

wire n5205;
// (3, 1, 'lutff_5/lout')

wire n5206;
// (22, 14, 'lutff_7/lout')

wire n5207;
// (15, 15, 'lutff_7/lout')

wire n5208;
// (5, 10, 'lutff_2/lout')

wire n5209;
// (7, 21, 'lutff_4/lout')

wire n5210;
// (11, 5, 'lutff_1/lout')

wire n5211;
// (8, 17, 'lutff_2/out')

wire n5212;
// (8, 17, 'lutff_2/lout')

wire n5213;
// (5, 13, 'lutff_7/lout')

wire n5214;
// (23, 19, 'lutff_3/lout')

wire n5215;
// (4, 9, 'lutff_6/lout')

wire n5216;
// (15, 8, 'lutff_4/lout')

wire n5217;
// (17, 19, 'lutff_6/lout')

wire n5218;
// (17, 11, 'lutff_2/lout')

wire n5219;
// (4, 6, 'lutff_0/lout')

wire n5220;
// (7, 14, 'lutff_1/lout')

wire n5221;
// (2, 6, 'lutff_7/lout')

wire n5222;
// (16, 20, 'lutff_2/lout')

wire n5223;
// (14, 12, 'lutff_5/lout')

wire n5224;
// (14, 4, 'lutff_1/lout')

wire n5225;
// (17, 20, 'lutff_7/lout')

wire n5226;
// (17, 12, 'lutff_3/lout')

wire n5227;
// (23, 3, 'lutff_0/lout')

wire n5228;
// (15, 4, 'lutff_6/lout')

wire n5229;
// (5, 6, 'lutff_3/lout')

wire n5230;
// (14, 13, 'lutff_6/lout')

wire n5231;
// (4, 2, 'lutff_2/lout')

wire n5232;
// (14, 5, 'lutff_2/lout')

wire n5233;
// (16, 16, 'lutff_4/lout')

wire n5234;
// (13, 21, 'lutff_3/lout')

wire n5235;
// (8, 5, 'lutff_5/lout')

wire n5236;
// (24, 3, 'lutff_4/lout')

wire n5237;
// (10, 14, 'lutff_2/lout')

wire n5238;
// (9, 18, 'lutff_5/out')

wire n5239;
// (9, 18, 'lutff_5/lout')

wire n5240;
// (9, 10, 'lutff_1/lout')

wire n5241;
// (16, 9, 'lutff_1/lout')

wire n5242;
// (7, 2, 'lutff_4/lout')

wire n5243;
// (8, 6, 'lutff_6/lout')

wire n5244;
// (16, 8, 'lutff_5/lout')

wire n5245;
// (10, 15, 'lutff_3/lout')

wire n5246;
// (20, 4, 'lutff_0/lout')

wire n5247;
// (18, 17, 'lutff_2/lout')

wire n5248;
// (13, 22, 'lutff_3/lout')

wire n5249;
// (2, 21, 'lutff_0/out')

wire n5250;
// (2, 21, 'lutff_0/lout')

wire n5251;
// (2, 21, 'carry_in_mux')

// Carry-In for (2 21)
assign n5251 = 1;

wire n5252;
// (9, 14, 'lutff_7/lout')

wire n5253;
// (20, 5, 'lutff_1/out')

wire n5254;
// (20, 5, 'lutff_1/lout')

wire n5255;
// (16, 4, 'lutff_7/lout')

wire n5256;
// (1, 8, 'lutff_5/lout')

wire n5257;
// (9, 11, 'lutff_1/lout')

wire n5258;
// (7, 3, 'lutff_4/lout')

wire n5259;
// (12, 18, 'lutff_6/lout')

wire n5260;
// (2, 13, 'lutff_1/lout')

wire n5261;
// (13, 6, 'lutff_0/lout')

wire n5262;
// (2, 16, 'lutff_6/lout')

wire n5263;
// (13, 9, 'lutff_5/lout')

wire n5264;
// (3, 12, 'lutff_4/lout')

wire n5265;
// (1, 4, 'lutff_7/lout')

wire n5266;
// (15, 18, 'lutff_2/lout')

wire n5267;
// (4, 17, 'lutff_0/lout')

wire n5268;
// (2, 17, 'lutff_7/lout')

wire n5269;
// (13, 10, 'lutff_6/lout')

wire n5270;
// (13, 2, 'lutff_2/lout')

wire n5271;
// (2, 9, 'lutff_3/lout')

wire n5272;
// (3, 13, 'lutff_5/out')

wire n5273;
// (3, 13, 'lutff_5/lout')

wire n5274;
// (3, 5, 'lutff_1/lout')

wire n5275;
// (11, 15, 'lutff_4/lout')

wire n5276;
// (14, 23, 'lutff_5/lout')

wire n5277;
// (11, 7, 'lutff_0/lout')

wire n5278;
// (15, 19, 'lutff_3/out')

wire n5279;
// (15, 19, 'lutff_3/lout')

wire n5280;
// (10, 3, 'lutff_5/lout')

wire n5281;
// (18, 6, 'lutff_6/lout')

wire n5282;
// (12, 7, 'lutff_5/lout')

wire n5283;
// (22, 9, 'lutff_3/lout')

wire n5284;
// (21, 13, 'lutff_6/lout')

wire n5285;
// (4, 21, 'lutff_6/lout')

wire n5286;
// (21, 5, 'lutff_2/lout')

wire n5287;
// (8, 16, 'lutff_5/lout')

wire n5288;
// (15, 3, 'lutff_0/lout')

wire n5289;
// (17, 22, 'lutff_6/lout')

wire n5290;
// (22, 2, 'lutff_0/lout')

wire n5291;
// (7, 17, 'lutff_1/lout')

wire n5292;
// (15, 6, 'lutff_5/lout')

wire n5293;
// (5, 9, 'lutff_4/lout')

wire n5294;
// (4, 13, 'lutff_7/lout')

wire n5295;
// (4, 5, 'lutff_3/lout')

wire n5296;
// (16, 19, 'lutff_5/lout')

wire n5297;
// (17, 15, 'lutff_3/lout')

wire n5298;
// (11, 3, 'lutff_7/lout')

wire n5299;
// (7, 18, 'lutff_2/out')

wire n5300;
// (7, 18, 'lutff_2/lout')

wire n5301;
// (15, 7, 'lutff_6/lout')

wire n5302;
// (9, 21, 'lutff_0/lout')

wire n5303;
// (7, 21, 'lutff_7/lout')

wire n5304;
// (14, 8, 'lutff_2/lout')

wire n5305;
// (8, 9, 'lutff_1/lout')

wire n5306;
// (20, 23, 'lutff_3/lout')

wire n5307;
// (17, 8, 'lutff_0/lout')

wire n5308;
// (5, 2, 'lutff_0/lout')

wire n5309;
// (23, 2, 'lutff_2/lout')

wire n5310;
// (4, 6, 'lutff_3/lout')

wire n5311;
// (17, 11, 'lutff_5/lout')

wire n5312;
// (9, 13, 'lutff_1/lout')

wire n5313;
// (16, 12, 'lutff_1/lout')

wire n5314;
// (13, 17, 'lutff_0/out')

wire n5315;
// (13, 17, 'lutff_0/lout')

wire n5316;
// (13, 17, 'carry_in_mux')

// Carry-In for (13 17)
assign n5316 = 1;

wire n5317;
// (7, 5, 'lutff_4/lout')

wire n5318;
// (14, 4, 'lutff_4/lout')

wire n5319;
// (8, 1, 'lutff_2/lout')

wire n5320;
// (1, 19, 'lutff_4/lout')

wire n5321;
// (23, 3, 'lutff_3/out')

wire n5322;
// (23, 3, 'lutff_3/lout')

wire n5323;
// (1, 11, 'lutff_0/lout')

wire n5324;
// (8, 4, 'lutff_7/lout')

wire n5325;
// (20, 7, 'lutff_0/out')

wire n5326;
// (20, 7, 'lutff_0/lout')

wire n5327;
// (20, 7, 'carry_in_mux')

// Carry-In for (20 7)
assign n5327 = 1;

wire n5328;
// (12, 21, 'lutff_1/lout')

wire n5329;
// (17, 3, 'lutff_6/lout')

wire n5330;
// (7, 6, 'lutff_5/lout')

wire n5331;
// (10, 13, 'lutff_4/lout')

wire n5332;
// (9, 17, 'lutff_7/lout')

wire n5333;
// (9, 9, 'lutff_3/lout')

wire n5334;
// (13, 21, 'lutff_6/lout')

wire n5335;
// (1, 12, 'lutff_1/lout')

wire n5336;
// (20, 8, 'lutff_1/out')

wire n5337;
// (20, 8, 'lutff_1/lout')

wire n5338;
// (12, 22, 'lutff_2/lout')

wire n5339;
// (20, 11, 'lutff_6/lout')

wire n5340;
// (10, 14, 'lutff_5/lout')

wire n5341;
// (10, 6, 'lutff_1/lout')

wire n5342;
// (18, 16, 'lutff_4/lout')

wire n5343;
// (9, 10, 'lutff_4/lout')

wire n5344;
// (9, 2, 'lutff_0/lout')

wire n5345;
// (22, 20, 'lutff_3/lout')

wire n5346;
// (7, 2, 'lutff_7/lout')

wire n5347;
// (21, 24, 'lutff_6/lout')

wire n5348;
// (2, 19, 'lutff_6/lout')

wire n5349;
// (13, 13, 'lutff_7/lout')

wire n5350;
// (3, 15, 'lutff_4/lout')

wire n5351;
// (20, 4, 'lutff_3/lout')

wire n5352;
// (3, 7, 'lutff_0/lout')

wire n5353;
// (11, 18, 'lutff_5/lout')

wire n5354;
// (18, 9, 'lutff_1/lout')

wire n5355;
// (4, 20, 'lutff_0/lout')

wire n5356;
// (2, 20, 'lutff_7/lout')

wire n5357;
// (12, 9, 'lutff_4/lout')

wire n5358;
// (22, 12, 'lutff_4/lout')

wire n5359;
// (2, 12, 'lutff_3/lout')

wire n5360;
// (13, 5, 'lutff_2/lout')

wire n5361;
// (3, 8, 'lutff_1/lout')

wire n5362;
// (21, 8, 'lutff_3/out')

wire n5363;
// (21, 8, 'lutff_3/lout')

wire n5364;
// (14, 18, 'lutff_1/lout')

wire n5365;
// (3, 11, 'lutff_6/lout')

wire n5366;
// (11, 14, 'lutff_7/lout')

wire n5367;
// (18, 1, 'lutff_2/lout')

wire n5368;
// (2, 13, 'lutff_4/lout')

wire n5369;
// (13, 6, 'lutff_3/lout')

wire n5370;
// (2, 5, 'lutff_0/lout')

wire n5371;
// (4, 16, 'lutff_2/lout')

wire n5372;
// (11, 11, 'lutff_1/out')

wire n5373;
// (11, 11, 'lutff_1/lout')

wire n5374;
// (14, 19, 'lutff_2/lout')

wire n5375;
// (22, 8, 'lutff_6/lout')

wire n5376;
// (15, 15, 'lutff_0/out')

wire n5377;
// (15, 15, 'lutff_0/lout')

wire n5378;
// (15, 15, 'carry_in_mux')

// Carry-In for (15 15)
assign n5378 = 1;

wire n5379;
// (3, 4, 'lutff_3/lout')

wire n5380;
// (21, 4, 'lutff_5/lout')

wire n5381;
// (15, 18, 'lutff_5/out')

wire n5382;
// (15, 18, 'lutff_5/lout')

wire n5383;
// (8, 19, 'lutff_5/out')

wire n5384;
// (8, 19, 'lutff_5/lout')

wire n5385;
// (22, 5, 'lutff_0/lout')

wire n5386;
// (7, 20, 'lutff_1/out')

wire n5387;
// (7, 20, 'lutff_1/lout')

wire n5388;
// (4, 8, 'lutff_3/lout')

wire n5389;
// (8, 20, 'lutff_6/lout')

wire n5390;
// (11, 7, 'lutff_3/lout')

wire n5391;
// (17, 18, 'lutff_3/lout')

wire n5392;
// (15, 10, 'lutff_6/lout')

wire n5393;
// (15, 2, 'lutff_2/lout')

wire n5394;
// (5, 5, 'lutff_1/lout')

wire n5395;
// (4, 1, 'lutff_0/lout')

wire n5396;
// (16, 15, 'lutff_2/lout')

wire n5397;
// (15, 3, 'lutff_3/lout')

wire n5398;
// (23, 13, 'lutff_6/lout')

wire n5399;
// (17, 14, 'lutff_5/lout')

wire n5400;
// (1, 14, 'lutff_1/lout')

wire n5401;
// (7, 17, 'lutff_4/lout')

wire n5402;
// (7, 9, 'lutff_0/out')

wire n5403;
// (7, 9, 'lutff_0/lout')

wire n5404;
// (7, 9, 'carry_in_mux')

// Carry-In for (7 9)
assign n5404 = 1;

wire n5405;
// (2, 1, 'lutff_6/lout')

wire n5406;
// (13, 20, 'lutff_0/out')

wire n5407;
// (13, 20, 'lutff_0/lout')

wire n5408;
// (13, 20, 'carry_in_mux')

// Carry-In for (13 20)
assign n5408 = 1;

wire n5409;
// (14, 7, 'lutff_4/lout')

wire n5410;
// (13, 23, 'lutff_5/lout')

wire n5411;
// (3, 18, 'lutff_0/out')

wire n5412;
// (3, 18, 'lutff_0/lout')

wire n5413;
// (3, 18, 'carry_in_mux')

// Carry-In for (3 18)
assign n5413 = 1;

wire n5414;
// (17, 6, 'lutff_6/out')

wire n5415;
// (17, 6, 'lutff_6/lout')

wire n5416;
// (10, 16, 'lutff_4/lout')

wire n5417;
// (7, 1, 'lutff_1/lout')

wire n5418;
// (9, 20, 'lutff_7/lout')

wire n5419;
// (9, 12, 'lutff_3/lout')

wire n5420;
// (7, 4, 'lutff_6/lout')

wire n5421;
// (3, 19, 'lutff_1/lout')

wire n5422;
// (20, 14, 'lutff_6/lout')

wire n5423;
// (10, 17, 'lutff_5/lout')

wire n5424;
// (20, 6, 'lutff_2/lout')

wire n5425;
// (10, 9, 'lutff_1/lout')

wire n5426;
// (9, 13, 'lutff_4/lout')

wire n5427;
// (9, 5, 'lutff_0/lout')

wire n5428;
// (7, 5, 'lutff_7/lout')

wire n5429;
// (20, 7, 'lutff_3/out')

wire n5430;
// (20, 7, 'lutff_3/lout')

wire n5431;
// (13, 8, 'lutff_3/lout')

wire n5432;
// (18, 12, 'lutff_1/lout')

wire n5433;
// (3, 14, 'lutff_7/lout')

wire n5434;
// (10, 1, 'lutff_2/lout')

wire n5435;
// (22, 15, 'lutff_4/lout')

wire n5436;
// (2, 15, 'lutff_3/lout')

wire n5437;
// (10, 4, 'lutff_7/lout')

wire n5438;
// (21, 11, 'lutff_3/lout')

wire n5439;
// (14, 21, 'lutff_1/lout')

wire n5440;
// (1, 3, 'lutff_4/lout')

wire n5441;
// (13, 4, 'lutff_5/lout')

wire n5442;
// (11, 17, 'lutff_7/lout')

wire n5443;
// (11, 9, 'lutff_3/lout')

wire n5444;
// (12, 13, 'lutff_5/lout')

wire n5445;
// (12, 5, 'lutff_1/lout')

wire n5446;
// (2, 8, 'lutff_0/out')

wire n5447;
// (2, 8, 'lutff_0/lout')

wire n5448;
// (2, 8, 'carry_in_mux')

// Carry-In for (2 8)
assign n5448 = 1;

wire n5449;
// (4, 19, 'lutff_2/lout')

wire n5450;
// (9, 1, 'lutff_7/lout')

wire n5451;
// (2, 11, 'lutff_5/lout')

wire n5452;
// (21, 7, 'lutff_5/out')

wire n5453;
// (21, 7, 'lutff_5/lout')

wire n5454;
// (11, 10, 'lutff_4/lout')

wire n5455;
// (15, 21, 'lutff_5/lout')

wire n5456;
// (12, 6, 'lutff_2/lout')

wire n5457;
// (15, 13, 'lutff_1/lout')

wire n5458;
// (5, 16, 'lutff_0/lout')

wire n5459;
// (12, 9, 'lutff_7/lout')

wire n5460;
// (22, 12, 'lutff_7/lout')

wire n5461;
// (22, 4, 'lutff_3/lout')

wire n5462;
// (2, 4, 'lutff_2/lout')

wire n5463;
// (21, 8, 'lutff_6/lout')

wire n5464;
// (4, 11, 'lutff_3/lout')

wire n5465;
// (8, 15, 'lutff_2/out')

wire n5466;
// (8, 15, 'lutff_2/lout')

wire n5467;
// (2, 3, 'lutff_6/lout')

wire n5468;
// (8, 18, 'lutff_7/lout')

wire n5469;
// (18, 1, 'lutff_5/lout')

wire n5470;
// (15, 5, 'lutff_2/lout')

wire n5471;
// (5, 8, 'lutff_1/lout')

wire n5472;
// (4, 4, 'lutff_0/lout')

wire n5473;
// (16, 18, 'lutff_2/lout')

wire n5474;
// (4, 7, 'lutff_5/lout')

wire n5475;
// (14, 10, 'lutff_5/lout')

wire n5476;
// (8, 11, 'lutff_4/lout')

wire n5477;
// (14, 2, 'lutff_1/lout')

wire n5478;
// (16, 21, 'lutff_7/lout')

wire n5479;
// (23, 8, 'lutff_2/lout')

wire n5480;
// (7, 20, 'lutff_4/out')

wire n5481;
// (7, 20, 'lutff_4/lout')

wire n5482;
// (17, 9, 'lutff_1/lout')

wire n5483;
// (5, 12, 'lutff_7/lout')

wire n5484;
// (5, 4, 'lutff_3/lout')

wire n5485;
// (4, 8, 'lutff_6/lout')

wire n5486;
// (16, 14, 'lutff_4/lout')

wire n5487;
// (17, 10, 'lutff_2/lout')

wire n5488;
// (14, 6, 'lutff_7/lout')

wire n5489;
// (3, 21, 'lutff_0/lout')

wire n5490;
// (8, 3, 'lutff_5/lout')

wire n5491;
// (1, 21, 'lutff_7/lout')

wire n5492;
// (15, 2, 'lutff_5/lout')

wire n5493;
// (18, 23, 'lutff_1/lout')

wire n5494;
// (1, 13, 'lutff_3/lout')

wire n5495;
// (20, 17, 'lutff_7/lout')

wire n5496;
// (14, 3, 'lutff_1/lout')

wire n5497;
// (12, 23, 'lutff_4/lout')

wire n5498;
// (13, 19, 'lutff_2/lout')

wire n5499;
// (7, 7, 'lutff_6/lout')

wire n5500;
// (1, 14, 'lutff_4/lout')

wire n5501;
// (16, 6, 'lutff_5/lout')

wire n5502;
// (1, 6, 'lutff_0/out')

wire n5503;
// (1, 6, 'lutff_0/lout')

wire n5504;
// (1, 6, 'carry_in_mux')

// Carry-In for (1 6)
assign n5504 = 1;

wire n5505;
// (10, 20, 'lutff_5/lout')

wire n5506;
// (10, 12, 'lutff_1/lout')

wire n5507;
// (9, 8, 'lutff_0/lout')

wire n5508;
// (13, 20, 'lutff_3/lout')

wire n5509;
// (7, 8, 'lutff_7/lout')

wire n5510;
// (18, 18, 'lutff_7/lout')

wire n5511;
// (20, 10, 'lutff_3/lout')

wire n5512;
// (16, 2, 'lutff_7/lout')

wire n5513;
// (12, 16, 'lutff_0/lout')

wire n5514;
// (3, 17, 'lutff_7/lout')

wire n5515;
// (10, 16, 'lutff_7/lout')

wire n5516;
// (22, 19, 'lutff_0/lout')

wire n5517;
// (9, 12, 'lutff_6/lout')

wire n5518;
// (5, 18, 'lutff_0/lout')

wire n5519;
// (11, 21, 'lutff_3/lout')

wire n5520;
// (12, 11, 'lutff_7/lout')

wire n5521;
// (13, 7, 'lutff_5/lout')

wire n5522;
// (3, 10, 'lutff_4/lout')

wire n5523;
// (3, 2, 'lutff_0/lout')

wire n5524;
// (18, 11, 'lutff_3/lout')

wire n5525;
// (1, 2, 'lutff_7/lout')

wire n5526;
// (12, 8, 'lutff_1/lout')

wire n5527;
// (15, 16, 'lutff_2/lout')

wire n5528;
// (9, 4, 'lutff_7/lout')

wire n5529;
// (22, 14, 'lutff_6/lout')

wire n5530;
// (2, 14, 'lutff_5/lout')

wire n5531;
// (13, 8, 'lutff_6/lout')

wire n5532;
// (21, 10, 'lutff_5/lout')

wire n5533;
// (21, 2, 'lutff_1/lout')

wire n5534;
// (11, 13, 'lutff_4/lout')

wire n5535;
// (11, 5, 'lutff_0/lout')

wire n5536;
// (5, 19, 'lutff_0/lout')

wire n5537;
// (10, 1, 'lutff_5/lout')

wire n5538;
// (12, 12, 'lutff_7/lout')

wire n5539;
// (22, 15, 'lutff_7/lout')

wire n5540;
// (2, 15, 'lutff_6/lout')

wire n5541;
// (12, 4, 'lutff_3/lout')

wire n5542;
// (22, 7, 'lutff_3/lout')

wire n5543;
// (2, 7, 'lutff_2/lout')

wire n5544;
// (21, 11, 'lutff_6/lout')

wire n5545;
// (21, 3, 'lutff_2/lout')

wire n5546;
// (11, 6, 'lutff_1/lout')

wire n5547;
// (5, 14, 'lutff_7/lout')

wire n5548;
// (8, 21, 'lutff_7/lout')

wire n5549;
// (17, 20, 'lutff_6/lout')

wire n5550;
// (15, 4, 'lutff_5/lout')

wire n5551;
// (5, 6, 'lutff_2/lout')

wire n5552;
// (4, 10, 'lutff_5/lout')

wire n5553;
// (14, 13, 'lutff_5/lout')

wire n5554;
// (4, 2, 'lutff_1/lout')

wire n5555;
// (8, 14, 'lutff_4/lout')

wire n5556;
// (14, 5, 'lutff_1/lout')

wire n5557;
// (16, 24, 'lutff_7/lout')

wire n5558;
// (16, 16, 'lutff_3/lout')

wire n5559;
// (11, 1, 'lutff_7/out')

wire n5560;
// (11, 1, 'lutff_7/lout')

wire n5561;
// (7, 15, 'lutff_0/out')

wire n5562;
// (7, 15, 'lutff_0/lout')

wire n5563;
// (7, 15, 'carry_in_mux')

// Carry-In for (7 15)
assign n5563 = 1;

wire n5564;
// (5, 15, 'lutff_7/lout')

wire n5565;
// (5, 7, 'lutff_3/lout')

wire n5566;
// (9, 19, 'lutff_0/out')

wire n5567;
// (9, 19, 'lutff_0/lout')

wire n5568;
// (4, 11, 'lutff_6/lout')

wire n5569;
// (4, 3, 'lutff_2/lout')

wire n5570;
// (8, 7, 'lutff_1/out')

wire n5571;
// (8, 7, 'lutff_1/lout')

wire n5572;
// (16, 9, 'lutff_0/lout')

wire n5573;
// (20, 21, 'lutff_3/lout')

wire n5574;
// (14, 9, 'lutff_7/lout')

wire n5575;
// (17, 13, 'lutff_2/lout')

wire n5576;
// (8, 6, 'lutff_5/lout')

wire n5577;
// (15, 5, 'lutff_5/lout')

wire n5578;
// (20, 20, 'lutff_7/lout')

wire n5579;
// (7, 11, 'lutff_2/lout')

wire n5580;
// (10, 15, 'lutff_2/lout')

wire n5581;
// (16, 10, 'lutff_1/lout')

wire n5582;
// (13, 22, 'lutff_2/lout')

wire n5583;
// (10, 18, 'lutff_7/out')

wire n5584;
// (10, 18, 'lutff_7/lout')

wire n5585;
// (14, 2, 'lutff_4/lout')

wire n5586;
// (1, 17, 'lutff_4/lout')

wire n5587;
// (1, 9, 'lutff_0/lout')

wire n5588;
// (8, 2, 'lutff_7/lout')

wire n5589;
// (20, 5, 'lutff_0/out')

wire n5590;
// (20, 5, 'lutff_0/lout')

wire n5591;
// (20, 5, 'carry_in_mux')

// Carry-In for (20 5)
assign n5591 = 1;

wire n5592;
// (12, 19, 'lutff_1/lout')

wire n5593;
// (7, 3, 'lutff_3/lout')

wire n5594;
// (10, 11, 'lutff_4/lout')

wire n5595;
// (18, 21, 'lutff_7/lout')

wire n5596;
// (9, 15, 'lutff_7/lout')

wire n5597;
// (1, 10, 'lutff_1/lout')

wire n5598;
// (13, 18, 'lutff_4/lout')

wire n5599;
// (3, 21, 'lutff_3/lout')

wire n5600;
// (1, 13, 'lutff_6/lout')

wire n5601;
// (16, 5, 'lutff_7/lout')

wire n5602;
// (17, 1, 'lutff_5/lout')

wire n5603;
// (20, 9, 'lutff_6/lout')

wire n5604;
// (18, 14, 'lutff_4/lout')

wire n5605;
// (9, 7, 'lutff_2/lout')

wire n5606;
// (13, 11, 'lutff_1/lout')

wire n5607;
// (21, 21, 'lutff_4/lout')

wire n5608;
// (2, 17, 'lutff_6/lout')

wire n5609;
// (13, 10, 'lutff_5/lout')

wire n5610;
// (3, 13, 'lutff_4/out')

wire n5611;
// (3, 13, 'lutff_4/lout')

wire n5612;
// (3, 5, 'lutff_0/lout')

wire n5613;
// (10, 4, 'lutff_0/lout')

wire n5614;
// (1, 5, 'lutff_7/lout')

wire n5615;
// (15, 19, 'lutff_2/lout')

wire n5616;
// (22, 18, 'lutff_2/lout')

wire n5617;
// (10, 3, 'lutff_4/lout')

wire n5618;
// (21, 14, 'lutff_1/lout')

wire n5619;
// (12, 7, 'lutff_4/lout')

wire n5620;
// (13, 3, 'lutff_2/lout')

wire n5621;
// (21, 13, 'lutff_5/lout')

wire n5622;
// (3, 6, 'lutff_1/lout')

wire n5623;
// (4, 21, 'lutff_5/lout')

wire n5624;
// (11, 8, 'lutff_0/lout')

wire n5625;
// (15, 20, 'lutff_3/lout')

wire n5626;
// (3, 9, 'lutff_6/lout')

wire n5627;
// (17, 23, 'lutff_1/lout')

wire n5628;
// (22, 10, 'lutff_3/lout')

wire n5629;
// (2, 10, 'lutff_2/lout')

wire n5630;
// (5, 18, 'lutff_3/lout')

wire n5631;
// (21, 6, 'lutff_2/lout')

wire n5632;
// (18, 2, 'lutff_7/lout')

wire n5633;
// (21, 9, 'lutff_7/lout')

wire n5634;
// (17, 24, 'lutff_2/lout')

wire n5635;
// (11, 12, 'lutff_6/lout')

wire n5636;
// (12, 8, 'lutff_4/lout')

wire n5637;
// (11, 4, 'lutff_2/lout')

wire n5638;
// (3, 1, 'lutff_7/lout')

wire n5639;
// (22, 3, 'lutff_0/lout')

wire n5640;
// (4, 14, 'lutff_1/lout')

wire n5641;
// (7, 18, 'lutff_1/out')

wire n5642;
// (7, 18, 'lutff_1/lout')

wire n5643;
// (22, 6, 'lutff_5/lout')

wire n5644;
// (5, 10, 'lutff_4/lout')

wire n5645;
// (21, 2, 'lutff_4/lout')

wire n5646;
// (7, 21, 'lutff_6/lout')

wire n5647;
// (8, 17, 'lutff_4/out')

wire n5648;
// (8, 17, 'lutff_4/lout')

wire n5649;
// (8, 9, 'lutff_0/out')

wire n5650;
// (8, 9, 'lutff_0/lout')

wire n5651;
// (8, 9, 'carry_in_mux')

// Carry-In for (8 9)
assign n5651 = 1;

wire n5652;
// (18, 3, 'lutff_7/lout')

wire n5653;
// (15, 8, 'lutff_6/lout')

wire n5654;
// (9, 22, 'lutff_0/out')

wire n5655;
// (9, 22, 'lutff_0/lout')

wire n5656;
// (9, 22, 'carry_in_mux')

// Carry-In for (9 22)
assign n5656 = 1;

wire n5657;
// (4, 6, 'lutff_2/lout')

wire n5658;
// (8, 10, 'lutff_1/lout')

wire n5659;
// (16, 20, 'lutff_4/lout')

wire n5660;
// (16, 12, 'lutff_0/lout')

wire n5661;
// (14, 12, 'lutff_7/lout')

wire n5662;
// (14, 4, 'lutff_3/lout')

wire n5663;
// (5, 3, 'lutff_0/lout')

wire n5664;
// (23, 3, 'lutff_2/lout')

wire n5665;
// (17, 12, 'lutff_5/lout')

wire n5666;
// (17, 4, 'lutff_1/lout')

wire n5667;
// (5, 6, 'lutff_5/lout')

wire n5668;
// (16, 13, 'lutff_1/lout')

wire n5669;
// (4, 2, 'lutff_4/lout')

wire n5670;
// (7, 6, 'lutff_4/lout')

wire n5671;
// (14, 5, 'lutff_4/lout')

wire n5672;
// (16, 16, 'lutff_6/lout')

wire n5673;
// (1, 12, 'lutff_0/lout')

wire n5674;
// (8, 5, 'lutff_7/lout')

wire n5675;
// (20, 8, 'lutff_0/lout')

wire n5676;
// (12, 22, 'lutff_1/lout')

wire n5677;
// (20, 11, 'lutff_5/lout')

wire n5678;
// (10, 14, 'lutff_4/lout')

wire n5679;
// (9, 18, 'lutff_7/out')

wire n5680;
// (9, 18, 'lutff_7/lout')

wire n5681;
// (9, 10, 'lutff_3/lout')

wire n5682;
// (22, 20, 'lutff_2/lout')

wire n5683;
// (7, 2, 'lutff_6/lout')

wire n5684;
// (21, 16, 'lutff_1/lout')

wire n5685;
// (16, 8, 'lutff_7/lout')

wire n5686;
// (20, 12, 'lutff_6/lout')

wire n5687;
// (10, 15, 'lutff_5/lout')

wire n5688;
// (10, 7, 'lutff_1/lout')

wire n5689;
// (18, 9, 'lutff_0/lout')

wire n5690;
// (22, 21, 'lutff_3/lout')

wire n5691;
// (2, 21, 'lutff_2/lout')

wire n5692;
// (20, 5, 'lutff_3/lout')

wire n5693;
// (3, 8, 'lutff_0/out')

wire n5694;
// (3, 8, 'lutff_0/lout')

wire n5695;
// (3, 8, 'carry_in_mux')

// Carry-In for (3 8)
assign n5695 = 1;

wire n5696;
// (1, 8, 'lutff_7/lout')

wire n5697;
// (18, 10, 'lutff_1/lout')

wire n5698;
// (12, 11, 'lutff_0/lout')

wire n5699;
// (21, 17, 'lutff_1/lout')

wire n5700;
// (12, 10, 'lutff_4/lout')

wire n5701;
// (13, 6, 'lutff_2/lout')

wire n5702;
// (10, 2, 'lutff_7/lout')

wire n5703;
// (11, 11, 'lutff_0/out')

wire n5704;
// (11, 11, 'lutff_0/lout')

wire n5705;
// (11, 11, 'carry_in_mux')

// Carry-In for (11 11)
assign n5705 = 1;

wire n5706;
// (13, 9, 'lutff_7/lout')

wire n5707;
// (14, 19, 'lutff_1/lout')

wire n5708;
// (3, 12, 'lutff_6/lout')

wire n5709;
// (3, 4, 'lutff_2/lout')

wire n5710;
// (15, 18, 'lutff_4/lout')

wire n5711;
// (12, 3, 'lutff_1/out')

wire n5712;
// (12, 3, 'lutff_1/lout')

wire n5713;
// (24, 17, 'lutff_3/lout')

wire n5714;
// (4, 17, 'lutff_2/lout')

wire n5715;
// (18, 5, 'lutff_7/lout')

wire n5716;
// (2, 9, 'lutff_5/lout')

wire n5717;
// (13, 2, 'lutff_4/lout')

wire n5718;
// (3, 5, 'lutff_3/lout')

wire n5719;
// (11, 15, 'lutff_6/lout')

wire n5720;
// (16, 23, 'lutff_0/lout')

wire n5721;
// (11, 7, 'lutff_2/lout')

wire n5722;
// (8, 20, 'lutff_5/lout')

wire n5723;
// (15, 19, 'lutff_5/lout')

wire n5724;
// (15, 11, 'lutff_1/lout')

wire n5725;
// (10, 3, 'lutff_7/lout')

wire n5726;
// (23, 21, 'lutff_4/lout')

wire n5727;
// (5, 14, 'lutff_0/lout')

wire n5728;
// (12, 7, 'lutff_7/lout')

wire n5729;
// (21, 5, 'lutff_4/lout')

wire n5730;
// (11, 8, 'lutff_3/lout')

wire n5731;
// (23, 14, 'lutff_1/lout')

wire n5732;
// (8, 16, 'lutff_7/lout')

wire n5733;
// (15, 3, 'lutff_2/lout')

wire n5734;
// (22, 2, 'lutff_2/lout')

wire n5735;
// (17, 14, 'lutff_4/lout')

wire n5736;
// (7, 17, 'lutff_3/lout')

wire n5737;
// (15, 6, 'lutff_7/lout')

wire n5738;
// (8, 13, 'lutff_1/lout')

wire n5739;
// (2, 1, 'lutff_5/lout')

wire n5740;
// (5, 9, 'lutff_6/lout')

wire n5741;
// (4, 5, 'lutff_5/lout')

wire n5742;
// (14, 7, 'lutff_3/lout')

wire n5743;
// (16, 19, 'lutff_7/lout')

wire n5744;
// (23, 6, 'lutff_2/lout')

wire n5745;
// (17, 7, 'lutff_1/lout')

wire n5746;
// (7, 18, 'lutff_4/out')

wire n5747;
// (7, 18, 'lutff_4/lout')

wire n5748;
// (5, 10, 'lutff_7/lout')

wire n5749;
// (9, 21, 'lutff_2/lout')

wire n5750;
// (20, 20, 'lutff_0/lout')

wire n5751;
// (14, 8, 'lutff_4/lout')

wire n5752;
// (8, 9, 'lutff_3/lout')

wire n5753;
// (13, 16, 'lutff_1/lout')

wire n5754;
// (8, 8, 'lutff_7/lout')

wire n5755;
// (3, 19, 'lutff_0/out')

wire n5756;
// (3, 19, 'lutff_0/lout')

wire n5757;
// (3, 19, 'carry_in_mux')

// Carry-In for (3 19)
assign n5757 = 1;

wire n5758;
// (5, 2, 'lutff_2/lout')

wire n5759;
// (23, 2, 'lutff_4/out')

wire n5760;
// (23, 2, 'lutff_4/lout')

wire n5761;
// (10, 17, 'lutff_4/lout')

wire n5762;
// (9, 13, 'lutff_3/lout')

wire n5763;
// (16, 12, 'lutff_3/lout')

wire n5764;
// (13, 17, 'lutff_2/lout')

wire n5765;
// (7, 5, 'lutff_6/lout')

wire n5766;
// (8, 1, 'lutff_4/lout')

wire n5767;
// (1, 19, 'lutff_6/lout')

wire n5768;
// (1, 11, 'lutff_2/lout')

wire n5769;
// (20, 7, 'lutff_2/lout')

wire n5770;
// (10, 10, 'lutff_1/lout')

wire n5771;
// (12, 21, 'lutff_3/lout')

wire n5772;
// (7, 6, 'lutff_7/lout')

wire n5773;
// (10, 13, 'lutff_6/lout')

wire n5774;
// (3, 20, 'lutff_0/lout')

wire n5775;
// (21, 20, 'lutff_2/lout')

wire n5776;
// (9, 9, 'lutff_5/lout')

wire n5777;
// (20, 8, 'lutff_3/out')

wire n5778;
// (20, 8, 'lutff_3/lout')

wire n5779;
// (21, 23, 'lutff_7/lout')

wire n5780;
// (12, 22, 'lutff_4/lout')

wire n5781;
// (18, 13, 'lutff_1/lout')

wire n5782;
// (12, 14, 'lutff_0/out')

wire n5783;
// (12, 14, 'lutff_0/lout')

wire n5784;
// (12, 14, 'carry_in_mux')

// Carry-In for (12 14)
assign n5784 = 1;

wire n5785;
// (10, 6, 'lutff_3/lout')

wire n5786;
// (18, 16, 'lutff_6/lout')

wire n5787;
// (9, 2, 'lutff_2/lout')

wire n5788;
// (21, 16, 'lutff_4/lout')

wire n5789;
// (3, 15, 'lutff_6/lout')

wire n5790;
// (3, 7, 'lutff_2/lout')

wire n5791;
// (11, 10, 'lutff_3/lout')

wire n5792;
// (18, 9, 'lutff_3/lout')

wire n5793;
// (12, 6, 'lutff_1/lout')

wire n5794;
// (15, 13, 'lutff_0/lout')

wire n5795;
// (4, 20, 'lutff_2/lout')

wire n5796;
// (12, 9, 'lutff_6/lout')

wire n5797;
// (2, 12, 'lutff_5/lout')

wire n5798;
// (13, 5, 'lutff_4/lout')

wire n5799;
// (22, 4, 'lutff_2/lout')

wire n5800;
// (3, 8, 'lutff_3/lout')

wire n5801;
// (2, 4, 'lutff_1/lout')

wire n5802;
// (21, 8, 'lutff_5/lout')

wire n5803;
// (14, 18, 'lutff_3/lout')

wire n5804;
// (15, 14, 'lutff_1/lout')

wire n5805;
// (5, 17, 'lutff_0/lout')

wire n5806;
// (12, 10, 'lutff_7/lout')

wire n5807;
// (18, 1, 'lutff_4/lout')

wire n5808;
// (12, 2, 'lutff_3/lout')

wire n5809;
// (2, 5, 'lutff_2/lout')

wire n5810;
// (24, 16, 'lutff_5/lout')

wire n5811;
// (4, 16, 'lutff_4/lout')

wire n5812;
// (11, 11, 'lutff_3/out')

wire n5813;
// (11, 11, 'lutff_3/lout')

wire n5814;
// (14, 19, 'lutff_4/lout')

wire n5815;
// (14, 11, 'lutff_0/lout')

wire n5816;
// (21, 4, 'lutff_7/lout')

wire n5817;
// (8, 19, 'lutff_7/out')

wire n5818;
// (8, 19, 'lutff_7/lout')

wire n5819;
// (20, 22, 'lutff_0/lout')

wire n5820;
// (8, 11, 'lutff_3/lout')

wire n5821;
// (22, 5, 'lutff_2/lout')

wire n5822;
// (21, 1, 'lutff_1/lout')

wire n5823;
// (7, 20, 'lutff_3/out')

wire n5824;
// (7, 20, 'lutff_3/lout')

wire n5825;
// (15, 9, 'lutff_7/lout')

wire n5826;
// (5, 12, 'lutff_6/lout')

wire n5827;
// (5, 4, 'lutff_2/lout')

wire n5828;
// (4, 8, 'lutff_5/lout')

wire n5829;
// (16, 14, 'lutff_3/lout')

wire n5830;
// (17, 18, 'lutff_5/lout')

wire n5831;
// (17, 10, 'lutff_1/lout')

wire n5832;
// (14, 6, 'lutff_6/lout')

wire n5833;
// (7, 13, 'lutff_0/lout')

wire n5834;
// (15, 2, 'lutff_4/lout')

wire n5835;
// (5, 5, 'lutff_3/lout')

wire n5836;
// (4, 1, 'lutff_2/lout')

wire n5837;
// (14, 3, 'lutff_0/lout')

wire n5838;
// (16, 15, 'lutff_4/lout')

wire n5839;
// (16, 7, 'lutff_0/lout')

wire n5840;
// (20, 18, 'lutff_1/lout')

wire n5841;
// (15, 3, 'lutff_5/lout')

wire n5842;
// (17, 14, 'lutff_7/lout')

wire n5843;
// (1, 14, 'lutff_3/lout')

wire n5844;
// (7, 9, 'lutff_2/lout')

wire n5845;
// (13, 20, 'lutff_2/lout')

wire n5846;
// (7, 8, 'lutff_6/lout')

wire n5847;
// (14, 7, 'lutff_6/lout')

wire n5848;
// (13, 23, 'lutff_7/lout')

wire n5849;
// (3, 18, 'lutff_2/lout')

wire n5850;
// (10, 16, 'lutff_6/lout')

wire n5851;
// (7, 1, 'lutff_3/lout')

wire n5852;
// (18, 19, 'lutff_7/lout')

wire n5853;
// (9, 12, 'lutff_5/lout')

wire n5854;
// (1, 15, 'lutff_3/lout')

wire n5855;
// (13, 16, 'lutff_4/lout')

wire n5856;
// (3, 19, 'lutff_3/lout')

wire n5857;
// (11, 21, 'lutff_2/lout')

wire n5858;
// (16, 3, 'lutff_7/lout')

wire n5859;
// (12, 17, 'lutff_0/lout')

wire n5860;
// (10, 17, 'lutff_7/lout')

wire n5861;
// (20, 6, 'lutff_4/lout')

wire n5862;
// (10, 9, 'lutff_3/lout')

wire n5863;
// (9, 13, 'lutff_6/lout')

wire n5864;
// (18, 11, 'lutff_2/lout')

wire n5865;
// (9, 5, 'lutff_2/lout')

wire n5866;
// (21, 19, 'lutff_4/lout')

wire n5867;
// (13, 8, 'lutff_5/lout')

wire n5868;
// (18, 20, 'lutff_7/lout')

wire n5869;
// (18, 12, 'lutff_3/lout')

wire n5870;
// (10, 1, 'lutff_4/lout')

wire n5871;
// (12, 12, 'lutff_6/lout')

wire n5872;
// (22, 15, 'lutff_6/lout')

wire n5873;
// (2, 7, 'lutff_1/lout')

wire n5874;
// (21, 11, 'lutff_5/lout')

wire n5875;
// (21, 3, 'lutff_1/out')

wire n5876;
// (21, 3, 'lutff_1/lout')

wire n5877;
// (1, 3, 'lutff_6/lout')

wire n5878;
// (14, 21, 'lutff_3/lout')

wire n5879;
// (11, 6, 'lutff_0/lout')

wire n5880;
// (13, 4, 'lutff_7/lout')

wire n5881;
// (5, 20, 'lutff_0/lout')

wire n5882;
// (17, 21, 'lutff_1/lout')

wire n5883;
// (11, 9, 'lutff_5/lout')

wire n5884;
// (12, 13, 'lutff_7/lout')

wire n5885;
// (12, 5, 'lutff_3/lout')

wire n5886;
// (2, 8, 'lutff_2/lout')

wire n5887;
// (13, 1, 'lutff_1/out')

wire n5888;
// (13, 1, 'lutff_1/lout')

wire n5889;
// (4, 19, 'lutff_4/lout')

wire n5890;
// (14, 22, 'lutff_4/lout')

wire n5891;
// (2, 11, 'lutff_7/lout')

wire n5892;
// (14, 14, 'lutff_0/lout')

wire n5893;
// (3, 7, 'lutff_5/lout')

wire n5894;
// (21, 7, 'lutff_7/out')

wire n5895;
// (21, 7, 'lutff_7/lout')

wire n5896;
// (11, 10, 'lutff_6/lout')

wire n5897;
// (8, 22, 'lutff_7/lout')

wire n5898;
// (15, 13, 'lutff_3/lout')

wire n5899;
// (5, 15, 'lutff_6/lout')

wire n5900;
// (22, 4, 'lutff_5/lout')

wire n5901;
// (4, 11, 'lutff_5/lout')

wire n5902;
// (11, 2, 'lutff_1/lout')

wire n5903;
// (8, 15, 'lutff_4/out')

wire n5904;
// (8, 15, 'lutff_4/lout')

wire n5905;
// (8, 7, 'lutff_0/out')

wire n5906;
// (8, 7, 'lutff_0/lout')

wire n5907;
// (8, 7, 'carry_in_mux')

// Carry-In for (8 7)
assign n5907 = 1;

wire n5908;
// (17, 13, 'lutff_1/lout')

wire n5909;
// (20, 21, 'lutff_2/lout')

wire n5910;
// (14, 9, 'lutff_6/lout')

wire n5911;
// (15, 5, 'lutff_4/lout')

wire n5912;
// (5, 8, 'lutff_3/lout')

wire n5913;
// (4, 4, 'lutff_2/lout')

wire n5914;
// (7, 11, 'lutff_1/lout')

wire n5915;
// (16, 18, 'lutff_4/lout')

wire n5916;
// (4, 7, 'lutff_7/lout')

wire n5917;
// (16, 10, 'lutff_0/lout')

wire n5918;
// (14, 10, 'lutff_7/lout')

wire n5919;
// (8, 11, 'lutff_6/lout')

wire n5920;
// (14, 2, 'lutff_3/lout')

wire n5921;
// (5, 1, 'lutff_0/lout')

wire n5922;
// (7, 20, 'lutff_6/out')

wire n5923;
// (7, 20, 'lutff_6/lout')

wire n5924;
// (17, 9, 'lutff_3/lout')

wire n5925;
// (7, 12, 'lutff_2/lout')

wire n5926;
// (5, 4, 'lutff_5/lout')

wire n5927;
// (16, 11, 'lutff_1/lout')

wire n5928;
// (10, 19, 'lutff_7/lout')

wire n5929;
// (16, 14, 'lutff_6/lout')

wire n5930;
// (9, 15, 'lutff_6/lout')

wire n5931;
// (1, 10, 'lutff_0/lout')

wire n5932;
// (17, 2, 'lutff_0/lout')

wire n5933;
// (3, 21, 'lutff_2/lout')

wire n5934;
// (8, 3, 'lutff_7/lout')

wire n5935;
// (1, 13, 'lutff_5/lout')

wire n5936;
// (12, 20, 'lutff_1/lout')

wire n5937;
// (20, 9, 'lutff_5/lout')

wire n5938;
// (9, 7, 'lutff_1/lout')

wire n5939;
// (13, 19, 'lutff_4/lout')

wire n5940;
// (21, 21, 'lutff_3/lout')

wire n5941;
// (1, 14, 'lutff_6/lout')

wire n5942;
// (16, 6, 'lutff_7/lout')

wire n5943;
// (1, 6, 'lutff_2/out')

wire n5944;
// (1, 6, 'lutff_2/lout')

wire n5945;
// (10, 20, 'lutff_7/lout')

wire n5946;
// (10, 12, 'lutff_3/lout')

wire n5947;
// (9, 8, 'lutff_2/lout')

wire n5948;
// (22, 18, 'lutff_1/lout')

wire n5949;
// (2, 18, 'lutff_0/lout')

wire n5950;
// (13, 12, 'lutff_1/lout')

wire n5951;
// (21, 14, 'lutff_0/lout')

wire n5952;
// (20, 10, 'lutff_5/lout')

wire n5953;
// (3, 6, 'lutff_0/lout')

wire n5954;
// (10, 5, 'lutff_0/lout')

wire n5955;
// (12, 16, 'lutff_2/lout')

wire n5956;
// (15, 20, 'lutff_2/lout')

wire n5957;
// (3, 9, 'lutff_5/lout')

wire n5958;
// (2, 10, 'lutff_1/lout')

wire n5959;
// (18, 8, 'lutff_0/lout')

wire n5960;
// (13, 7, 'lutff_7/lout')

wire n5961;
// (3, 2, 'lutff_2/lout')

wire n5962;
// (11, 12, 'lutff_5/lout')

wire n5963;
// (18, 11, 'lutff_5/lout')

wire n5964;
// (12, 8, 'lutff_3/lout')

wire n5965;
// (15, 16, 'lutff_4/lout')

wire n5966;
// (4, 14, 'lutff_0/lout')

wire n5967;
// (2, 14, 'lutff_7/lout')

wire n5968;
// (21, 2, 'lutff_3/lout')

wire n5969;
// (11, 5, 'lutff_2/lout')

wire n5970;
// (12, 1, 'lutff_0/out')

wire n5971;
// (12, 1, 'lutff_0/lout')

wire n5972;
// (12, 1, 'carry_in_mux')

// Carry-In for (12 1)
assign n5972 = 1;

wire n5973;
// (5, 19, 'lutff_2/lout')

wire n5974;
// (10, 1, 'lutff_7/lout')

wire n5975;
// (4, 15, 'lutff_1/lout')

wire n5976;
// (12, 4, 'lutff_5/lout')

wire n5977;
// (22, 7, 'lutff_5/lout')

wire n5978;
// (2, 7, 'lutff_4/lout')

wire n5979;
// (21, 3, 'lutff_4/lout')

wire n5980;
// (14, 21, 'lutff_6/lout')

wire n5981;
// (11, 6, 'lutff_3/lout')

wire n5982;
// (8, 10, 'lutff_0/lout')

wire n5983;
// (15, 9, 'lutff_0/lout')

wire n5984;
// (17, 12, 'lutff_4/lout')

wire n5985;
// (17, 4, 'lutff_0/lout')

wire n5986;
// (15, 4, 'lutff_7/lout')

wire n5987;
// (5, 6, 'lutff_4/lout')

wire n5988;
// (4, 10, 'lutff_7/lout')

wire n5989;
// (16, 13, 'lutff_0/lout')

wire n5990;
// (14, 13, 'lutff_7/lout')

wire n5991;
// (4, 2, 'lutff_3/lout')

wire n5992;
// (8, 14, 'lutff_6/lout')

wire n5993;
// (14, 5, 'lutff_3/lout')

wire n5994;
// (23, 12, 'lutff_0/out')

wire n5995;
// (23, 12, 'lutff_0/lout')

wire n5996;
// (23, 12, 'carry_in_mux')

// Carry-In for (23 12)
assign n5996 = 1;

wire n5997;
// (7, 15, 'lutff_2/out')

wire n5998;
// (7, 15, 'lutff_2/lout')

wire n5999;
// (5, 7, 'lutff_5/lout')

wire n6000;
// (9, 19, 'lutff_2/lout')

wire n6001;
// (4, 3, 'lutff_4/lout')

wire n6002;
// (16, 9, 'lutff_2/lout')

wire n6003;
// (17, 13, 'lutff_4/lout')

wire n6004;
// (17, 5, 'lutff_0/lout')

wire n6005;
// (20, 13, 'lutff_1/lout')

wire n6006;
// (8, 6, 'lutff_7/lout')

wire n6007;
// (15, 5, 'lutff_7/lout')

wire n6008;
// (10, 15, 'lutff_4/lout')

wire n6009;
// (10, 7, 'lutff_0/lout')

wire n6010;
// (13, 22, 'lutff_4/lout')

wire n6011;
// (2, 21, 'lutff_1/lout')

wire n6012;
// (13, 14, 'lutff_0/lout')

wire n6013;
// (1, 17, 'lutff_6/lout')

wire n6014;
// (1, 9, 'lutff_2/lout')

wire n6015;
// (20, 5, 'lutff_2/lout')

wire n6016;
// (9, 11, 'lutff_2/lout')

wire n6017;
// (12, 19, 'lutff_3/lout')

wire n6018;
// (18, 10, 'lutff_0/lout')

wire n6019;
// (13, 15, 'lutff_1/lout')

wire n6020;
// (7, 3, 'lutff_5/lout')

wire n6021;
// (10, 11, 'lutff_6/lout')

wire n6022;
// (13, 18, 'lutff_6/lout')

wire n6023;
// (10, 8, 'lutff_0/lout')

wire n6024;
// (21, 21, 'lutff_6/lout')

wire n6025;
// (4, 17, 'lutff_1/lout')

wire n6026;
// (11, 16, 'lutff_1/lout')

wire n6027;
// (13, 10, 'lutff_7/lout')

wire n6028;
// (2, 9, 'lutff_4/lout')

wire n6029;
// (13, 2, 'lutff_3/lout')

wire n6030;
// (3, 13, 'lutff_6/lout')

wire n6031;
// (3, 5, 'lutff_2/lout')

wire n6032;
// (14, 23, 'lutff_6/lout')

wire n6033;
// (15, 19, 'lutff_4/lout')

wire n6034;
// (15, 11, 'lutff_0/lout')

wire n6035;
// (10, 3, 'lutff_6/lout')

wire n6036;
// (12, 7, 'lutff_6/lout')

wire n6037;
// (14, 20, 'lutff_0/lout')

wire n6038;
// (22, 9, 'lutff_4/lout')

wire n6039;
// (13, 3, 'lutff_4/lout')

wire n6040;
// (21, 13, 'lutff_7/lout')

wire n6041;
// (3, 6, 'lutff_3/lout')

wire n6042;
// (21, 5, 'lutff_3/lout')

wire n6043;
// (4, 21, 'lutff_7/lout')

wire n6044;
// (11, 8, 'lutff_2/lout')

wire n6045;
// (15, 20, 'lutff_5/lout')

wire n6046;
// (15, 12, 'lutff_1/lout')

wire n6047;
// (23, 14, 'lutff_0/lout')

wire n6048;
// (4, 18, 'lutff_1/out')

wire n6049;
// (4, 18, 'lutff_1/lout')

wire n6050;
// (22, 10, 'lutff_5/lout')

wire n6051;
// (2, 10, 'lutff_4/lout')

wire n6052;
// (22, 2, 'lutff_1/lout')

wire n6053;
// (2, 2, 'lutff_0/lout')

wire n6054;
// (21, 6, 'lutff_4/lout')

wire n6055;
// (8, 13, 'lutff_0/lout')

wire n6056;
// (11, 4, 'lutff_4/lout')

wire n6057;
// (22, 3, 'lutff_2/lout')

wire n6058;
// (17, 15, 'lutff_4/lout')

wire n6059;
// (7, 18, 'lutff_3/out')

wire n6060;
// (7, 18, 'lutff_3/lout')

wire n6061;
// (22, 6, 'lutff_7/lout')

wire n6062;
// (15, 7, 'lutff_7/lout')

wire n6063;
// (9, 21, 'lutff_1/lout')

wire n6064;
// (8, 17, 'lutff_6/out')

wire n6065;
// (8, 17, 'lutff_6/lout')

wire n6066;
// (14, 8, 'lutff_3/lout')

wire n6067;
// (8, 9, 'lutff_2/lout')

wire n6068;
// (23, 11, 'lutff_3/lout')

wire n6069;
// (20, 23, 'lutff_4/lout')

wire n6070;
// (17, 8, 'lutff_1/lout')

wire n6071;
// (9, 22, 'lutff_2/lout')

wire n6072;
// (17, 11, 'lutff_6/lout')

wire n6073;
// (4, 6, 'lutff_4/lout')

wire n6074;
// (8, 10, 'lutff_3/lout')

wire n6075;
// (14, 1, 'lutff_0/lout')

wire n6076;
// (16, 20, 'lutff_6/lout')

wire n6077;
// (1, 20, 'lutff_1/lout')

wire n6078;
// (16, 12, 'lutff_2/lout')

wire n6079;
// (14, 4, 'lutff_5/lout')

wire n6080;
// (10, 19, 'lutff_0/lout')

wire n6081;
// (1, 19, 'lutff_5/lout')

wire n6082;
// (5, 3, 'lutff_2/lout')

wire n6083;
// (23, 3, 'lutff_4/lout')

wire n6084;
// (17, 4, 'lutff_3/lout')

wire n6085;
// (5, 6, 'lutff_7/lout')

wire n6086;
// (16, 13, 'lutff_3/lout')

wire n6087;
// (4, 2, 'lutff_6/lout')

wire n6088;
// (14, 5, 'lutff_6/lout')

wire n6089;
// (1, 12, 'lutff_2/lout')

wire n6090;
// (13, 21, 'lutff_7/lout')

wire n6091;
// (20, 8, 'lutff_2/lout')

wire n6092;
// (12, 22, 'lutff_3/lout')

wire n6093;
// (20, 11, 'lutff_7/lout')

wire n6094;
// (10, 14, 'lutff_6/lout')

wire n6095;
// (10, 6, 'lutff_2/lout')

wire n6096;
// (9, 10, 'lutff_5/lout')

wire n6097;
// (9, 2, 'lutff_1/lout')

wire n6098;
// (22, 20, 'lutff_4/lout')

wire n6099;
// (3, 16, 'lutff_1/lout')

wire n6100;
// (21, 16, 'lutff_3/lout')

wire n6101;
// (12, 15, 'lutff_0/lout')

wire n6102;
// (20, 4, 'lutff_4/lout')

wire n6103;
// (10, 15, 'lutff_7/lout')

wire n6104;
// (10, 7, 'lutff_3/lout')

wire n6105;
// (18, 17, 'lutff_6/lout')

wire n6106;
// (18, 9, 'lutff_2/lout')

wire n6107;
// (3, 8, 'lutff_2/lout')

wire n6108;
// (18, 10, 'lutff_3/lout')

wire n6109;
// (9, 3, 'lutff_1/lout')

wire n6110;
// (15, 22, 'lutff_4/lout')

wire n6111;
// (3, 11, 'lutff_7/lout')

wire n6112;
// (15, 14, 'lutff_0/lout')

wire n6113;
// (21, 17, 'lutff_3/lout')

wire n6114;
// (2, 13, 'lutff_5/lout')

wire n6115;
// (12, 2, 'lutff_2/lout')

wire n6116;
// (13, 6, 'lutff_4/lout')

wire n6117;
// (4, 16, 'lutff_3/lout')

wire n6118;
// (11, 11, 'lutff_2/lout')

wire n6119;
// (14, 19, 'lutff_3/lout')

wire n6120;
// (22, 8, 'lutff_7/lout')

wire n6121;
// (15, 15, 'lutff_1/out')

wire n6122;
// (15, 15, 'lutff_1/lout')

wire n6123;
// (3, 4, 'lutff_4/lout')

wire n6124;
// (21, 4, 'lutff_6/lout')

wire n6125;
// (15, 18, 'lutff_6/lout')

wire n6126;
// (12, 3, 'lutff_3/out')

wire n6127;
// (12, 3, 'lutff_3/lout')

wire n6128;
// (22, 5, 'lutff_1/lout')

wire n6129;
// (5, 13, 'lutff_1/lout')

wire n6130;
// (4, 17, 'lutff_4/lout')

wire n6131;
// (21, 1, 'lutff_0/lout')

wire n6132;
// (2, 9, 'lutff_7/lout')

wire n6133;
// (13, 2, 'lutff_6/lout')

wire n6134;
// (17, 19, 'lutff_0/out')

wire n6135;
// (17, 19, 'lutff_0/lout')

wire n6136;
// (17, 19, 'carry_in_mux')

// Carry-In for (17 19)
assign n6136 = 1;

wire n6137;
// (11, 7, 'lutff_4/lout')

wire n6138;
// (8, 20, 'lutff_7/lout')

wire n6139;
// (15, 11, 'lutff_3/lout')

wire n6140;
// (14, 20, 'lutff_3/lout')

wire n6141;
// (15, 10, 'lutff_7/lout')

wire n6142;
// (22, 9, 'lutff_7/lout')

wire n6143;
// (21, 5, 'lutff_6/lout')

wire n6144;
// (5, 5, 'lutff_2/lout')

wire n6145;
// (4, 1, 'lutff_1/lout')

wire n6146;
// (8, 12, 'lutff_2/lout')

wire n6147;
// (16, 15, 'lutff_3/lout')

wire n6148;
// (20, 18, 'lutff_0/lout')

wire n6149;
// (15, 3, 'lutff_4/lout')

wire n6150;
// (17, 14, 'lutff_6/lout')

wire n6151;
// (7, 17, 'lutff_5/lout')

wire n6152;
// (7, 9, 'lutff_1/lout')

wire n6153;
// (2, 1, 'lutff_7/lout')

wire n6154;
// (8, 13, 'lutff_3/lout')

wire n6155;
// (4, 5, 'lutff_7/lout')

wire n6156;
// (20, 19, 'lutff_1/lout')

wire n6157;
// (14, 7, 'lutff_5/lout')

wire n6158;
// (17, 15, 'lutff_7/lout')

wire n6159;
// (17, 7, 'lutff_3/lout')

wire n6160;
// (9, 21, 'lutff_4/lout')

wire n6161;
// (14, 8, 'lutff_6/lout')

wire n6162;
// (1, 15, 'lutff_2/lout')

wire n6163;
// (13, 16, 'lutff_3/lout')

wire n6164;
// (3, 19, 'lutff_2/lout')

wire n6165;
// (23, 2, 'lutff_6/out')

wire n6166;
// (23, 2, 'lutff_6/lout')

wire n6167;
// (20, 14, 'lutff_7/lout')

wire n6168;
// (10, 9, 'lutff_2/lout')

wire n6169;
// (9, 13, 'lutff_5/lout')

wire n6170;
// (9, 5, 'lutff_1/lout')

wire n6171;
// (13, 17, 'lutff_4/lout')

wire n6172;
// (16, 4, 'lutff_1/lout')

wire n6173;
// (8, 1, 'lutff_6/lout')

wire n6174;
// (21, 19, 'lutff_3/lout')

wire n6175;
// (12, 18, 'lutff_0/lout')

wire n6176;
// (20, 7, 'lutff_4/lout')

wire n6177;
// (10, 10, 'lutff_3/lout')

wire n6178;
// (12, 21, 'lutff_5/lout')

wire n6179;
// (18, 12, 'lutff_2/lout')

wire n6180;
// (9, 6, 'lutff_2/lout')

wire n6181;
// (2, 16, 'lutff_0/lout')

wire n6182;
// (21, 20, 'lutff_4/lout')

wire n6183;
// (9, 9, 'lutff_7/lout')

wire n6184;
// (21, 12, 'lutff_0/lout')

wire n6185;
// (1, 4, 'lutff_1/lout')

wire n6186;
// (20, 8, 'lutff_5/lout')

wire n6187;
// (18, 13, 'lutff_3/lout')

wire n6188;
// (1, 3, 'lutff_5/lout')

wire n6189;
// (12, 14, 'lutff_2/lout')

wire n6190;
// (12, 13, 'lutff_6/lout')

wire n6191;
// (22, 20, 'lutff_7/lout')

wire n6192;
// (2, 8, 'lutff_1/out')

wire n6193;
// (2, 8, 'lutff_1/lout')

wire n6194;
// (13, 1, 'lutff_0/out')

wire n6195;
// (13, 1, 'lutff_0/lout')

wire n6196;
// (13, 1, 'carry_in_mux')

// Carry-In for (13 1)
assign n6196 = 1;

wire n6197;
// (4, 19, 'lutff_3/out')

wire n6198;
// (4, 19, 'lutff_3/lout')

wire n6199;
// (14, 22, 'lutff_3/lout')

wire n6200;
// (18, 6, 'lutff_0/out')

wire n6201;
// (18, 6, 'lutff_0/lout')

wire n6202;
// (18, 6, 'carry_in_mux')

// Carry-In for (18 6)
assign n6202 = 1;

wire n6203;
// (2, 11, 'lutff_6/lout')

wire n6204;
// (3, 7, 'lutff_4/lout')

wire n6205;
// (11, 10, 'lutff_5/lout')

wire n6206;
// (18, 9, 'lutff_5/lout')

wire n6207;
// (12, 6, 'lutff_3/lout')

wire n6208;
// (15, 13, 'lutff_2/lout')

wire n6209;
// (4, 20, 'lutff_4/lout')

wire n6210;
// (4, 12, 'lutff_0/out')

wire n6211;
// (4, 12, 'lutff_0/lout')

wire n6212;
// (4, 12, 'carry_in_mux')

// Carry-In for (4 12)
assign n6212 = 1;

wire n6213;
// (2, 12, 'lutff_7/lout')

wire n6214;
// (13, 5, 'lutff_6/lout')

wire n6215;
// (14, 15, 'lutff_0/lout')

wire n6216;
// (2, 4, 'lutff_3/lout')

wire n6217;
// (3, 8, 'lutff_5/lout')

wire n6218;
// (21, 8, 'lutff_7/lout')

wire n6219;
// (22, 4, 'lutff_4/lout')

wire n6220;
// (14, 18, 'lutff_5/lout')

wire n6221;
// (11, 2, 'lutff_0/lout')

wire n6222;
// (15, 14, 'lutff_3/lout')

wire n6223;
// (4, 13, 'lutff_1/out')

wire n6224;
// (4, 13, 'lutff_1/lout')

wire n6225;
// (4, 16, 'lutff_6/lout')

wire n6226;
// (11, 11, 'lutff_5/lout')

wire n6227;
// (11, 3, 'lutff_1/lout')

wire n6228;
// (14, 11, 'lutff_2/lout')

wire n6229;
// (8, 11, 'lutff_5/lout')

wire n6230;
// (7, 20, 'lutff_5/out')

wire n6231;
// (7, 20, 'lutff_5/lout')

wire n6232;
// (7, 12, 'lutff_1/lout')

wire n6233;
// (5, 4, 'lutff_4/lout')

wire n6234;
// (4, 8, 'lutff_7/lout')

wire n6235;
// (16, 11, 'lutff_0/lout')

wire n6236;
// (16, 14, 'lutff_5/lout')

wire n6237;
// (17, 18, 'lutff_7/lout')

wire n6238;
// (17, 10, 'lutff_3/lout')

wire n6239;
// (7, 13, 'lutff_2/lout')

wire n6240;
// (15, 2, 'lutff_6/lout')

wire n6241;
// (5, 5, 'lutff_5/lout')

wire n6242;
// (9, 16, 'lutff_0/out')

wire n6243;
// (9, 16, 'lutff_0/lout')

wire n6244;
// (9, 16, 'carry_in_mux')

// Carry-In for (9 16)
assign n6244 = 1;

wire n6245;
// (7, 16, 'lutff_7/lout')

wire n6246;
// (4, 1, 'lutff_4/lout')

wire n6247;
// (14, 3, 'lutff_2/lout')

wire n6248;
// (8, 4, 'lutff_1/lout')

wire n6249;
// (16, 15, 'lutff_6/lout')

wire n6250;
// (16, 7, 'lutff_2/lout')

wire n6251;
// (13, 19, 'lutff_3/lout')

wire n6252;
// (20, 18, 'lutff_3/lout')

wire n6253;
// (17, 3, 'lutff_0/lout')

wire n6254;
// (23, 5, 'lutff_6/lout')

wire n6255;
// (1, 14, 'lutff_5/lout')

wire n6256;
// (1, 6, 'lutff_1/out')

wire n6257;
// (1, 6, 'lutff_1/lout')

wire n6258;
// (10, 20, 'lutff_6/lout')

wire n6259;
// (9, 8, 'lutff_1/lout')

wire n6260;
// (13, 20, 'lutff_4/lout')

wire n6261;
// (13, 12, 'lutff_0/lout')

wire n6262;
// (3, 18, 'lutff_4/lout')

wire n6263;
// (20, 2, 'lutff_0/lout')

wire n6264;
// (12, 16, 'lutff_1/lout')

wire n6265;
// (22, 19, 'lutff_1/lout')

wire n6266;
// (2, 19, 'lutff_0/out')

wire n6267;
// (2, 19, 'lutff_0/lout')

wire n6268;
// (2, 19, 'carry_in_mux')

// Carry-In for (2 19)
assign n6268 = 1;

wire n6269;
// (7, 1, 'lutff_5/lout')

wire n6270;
// (13, 13, 'lutff_1/lout')

wire n6271;
// (9, 12, 'lutff_7/lout')

wire n6272;
// (21, 15, 'lutff_0/lout')

wire n6273;
// (1, 7, 'lutff_1/lout')

wire n6274;
// (13, 16, 'lutff_6/lout')

wire n6275;
// (20, 3, 'lutff_1/lout')

wire n6276;
// (11, 21, 'lutff_4/lout')

wire n6277;
// (12, 17, 'lutff_2/lout')

wire n6278;
// (20, 6, 'lutff_6/lout')

wire n6279;
// (10, 9, 'lutff_5/lout')

wire n6280;
// (18, 11, 'lutff_4/lout')

wire n6281;
// (9, 5, 'lutff_4/lout')

wire n6282;
// (11, 14, 'lutff_1/lout')

wire n6283;
// (2, 14, 'lutff_6/lout')

wire n6284;
// (13, 8, 'lutff_7/lout')

wire n6285;
// (11, 13, 'lutff_5/lout')

wire n6286;
// (18, 12, 'lutff_5/lout')

wire n6287;
// (18, 4, 'lutff_1/lout')

wire n6288;
// (5, 19, 'lutff_1/lout')

wire n6289;
// (10, 1, 'lutff_6/lout')

wire n6290;
// (24, 15, 'lutff_1/lout')

wire n6291;
// (4, 15, 'lutff_0/lout')

wire n6292;
// (2, 15, 'lutff_7/lout')

wire n6293;
// (12, 4, 'lutff_4/lout')

wire n6294;
// (22, 7, 'lutff_4/lout')

wire n6295;
// (2, 7, 'lutff_3/lout')

wire n6296;
// (3, 3, 'lutff_1/lout')

wire n6297;
// (21, 3, 'lutff_3/lout')

wire n6298;
// (14, 21, 'lutff_5/lout')

wire n6299;
// (11, 6, 'lutff_2/lout')

wire n6300;
// (5, 20, 'lutff_2/lout')

wire n6301;
// (17, 21, 'lutff_3/lout')

wire n6302;
// (11, 9, 'lutff_7/lout')

wire n6303;
// (12, 5, 'lutff_5/lout')

wire n6304;
// (2, 8, 'lutff_4/lout')

wire n6305;
// (13, 1, 'lutff_3/out')

wire n6306;
// (13, 1, 'lutff_3/lout')

wire n6307;
// (4, 19, 'lutff_6/lout')

wire n6308;
// (14, 22, 'lutff_6/lout')

wire n6309;
// (14, 14, 'lutff_2/lout')

wire n6310;
// (15, 10, 'lutff_0/lout')

wire n6311;
// (8, 14, 'lutff_5/lout')

wire n6312;
// (15, 13, 'lutff_5/lout')

wire n6313;
// (23, 16, 'lutff_6/lout')

wire n6314;
// (7, 15, 'lutff_1/out')

wire n6315;
// (7, 15, 'lutff_1/lout')

wire n6316;
// (5, 7, 'lutff_4/lout')

wire n6317;
// (9, 19, 'lutff_1/lout')

wire n6318;
// (4, 11, 'lutff_7/lout')

wire n6319;
// (23, 13, 'lutff_0/lout')

wire n6320;
// (11, 2, 'lutff_3/lout')

wire n6321;
// (4, 3, 'lutff_3/lout')

wire n6322;
// (8, 15, 'lutff_6/out')

wire n6323;
// (8, 15, 'lutff_6/lout')

wire n6324;
// (8, 7, 'lutff_2/out')

wire n6325;
// (8, 7, 'lutff_2/lout')

wire n6326;
// (16, 17, 'lutff_5/lout')

wire n6327;
// (17, 13, 'lutff_3/lout')

wire n6328;
// (20, 13, 'lutff_0/lout')

wire n6329;
// (15, 5, 'lutff_6/lout')

wire n6330;
// (5, 8, 'lutff_5/lout')

wire n6331;
// (7, 19, 'lutff_7/lout')

wire n6332;
// (16, 18, 'lutff_6/lout')

wire n6333;
// (16, 10, 'lutff_2/lout')

wire n6334;
// (17, 6, 'lutff_0/out')

wire n6335;
// (17, 6, 'lutff_0/lout')

wire n6336;
// (17, 6, 'carry_in_mux')

// Carry-In for (17 6)
assign n6336 = 0;

wire n6337;
// (14, 2, 'lutff_5/lout')

wire n6338;
// (9, 20, 'lutff_1/out')

wire n6339;
// (9, 20, 'lutff_1/lout')

wire n6340;
// (1, 17, 'lutff_5/lout')

wire n6341;
// (17, 9, 'lutff_5/lout')

wire n6342;
// (7, 12, 'lutff_4/lout')

wire n6343;
// (7, 4, 'lutff_0/lout')

wire n6344;
// (13, 15, 'lutff_0/out')

wire n6345;
// (13, 15, 'lutff_0/lout')

wire n6346;
// (13, 15, 'carry_in_mux')

// Carry-In for (13 15)
assign n6346 = 1;

wire n6347;
// (10, 11, 'lutff_5/lout')

wire n6348;
// (13, 18, 'lutff_5/lout')

wire n6349;
// (3, 21, 'lutff_4/lout')

wire n6350;
// (1, 13, 'lutff_7/lout')

wire n6351;
// (20, 9, 'lutff_7/lout')

wire n6352;
// (21, 18, 'lutff_0/lout')

wire n6353;
// (13, 19, 'lutff_6/lout')

wire n6354;
// (13, 11, 'lutff_2/lout')

wire n6355;
// (21, 21, 'lutff_5/lout')

wire n6356;
// (3, 14, 'lutff_1/out')

wire n6357;
// (3, 14, 'lutff_1/lout')

wire n6358;
// (11, 16, 'lutff_0/lout')

wire n6359;
// (1, 6, 'lutff_4/out')

wire n6360;
// (1, 6, 'lutff_4/lout')

wire n6361;
// (10, 12, 'lutff_5/lout')

wire n6362;
// (10, 4, 'lutff_1/lout')

wire n6363;
// (9, 8, 'lutff_4/lout')

wire n6364;
// (22, 18, 'lutff_3/lout')

wire n6365;
// (2, 18, 'lutff_2/lout')

wire n6366;
// (21, 14, 'lutff_2/lout')

wire n6367;
// (13, 3, 'lutff_3/lout')

wire n6368;
// (3, 6, 'lutff_2/lout')

wire n6369;
// (18, 15, 'lutff_5/lout')

wire n6370;
// (3, 9, 'lutff_7/lout')

wire n6371;
// (15, 12, 'lutff_0/lout')

wire n6372;
// (17, 23, 'lutff_2/lout')

wire n6373;
// (4, 18, 'lutff_0/out')

wire n6374;
// (4, 18, 'lutff_0/lout')

wire n6375;
// (4, 18, 'carry_in_mux')

// Carry-In for (4 18)
assign n6375 = 1;

wire n6376;
// (22, 10, 'lutff_4/lout')

wire n6377;
// (2, 10, 'lutff_3/lout')

wire n6378;
// (5, 18, 'lutff_4/lout')

wire n6379;
// (21, 6, 'lutff_3/lout')

wire n6380;
// (14, 16, 'lutff_1/lout')

wire n6381;
// (3, 2, 'lutff_4/lout')

wire n6382;
// (11, 12, 'lutff_7/lout')

wire n6383;
// (23, 15, 'lutff_0/lout')

wire n6384;
// (11, 4, 'lutff_3/lout')

wire n6385;
// (12, 8, 'lutff_5/lout')

wire n6386;
// (15, 16, 'lutff_6/lout')

wire n6387;
// (2, 3, 'lutff_0/lout')

wire n6388;
// (4, 14, 'lutff_2/lout')

wire n6389;
// (8, 18, 'lutff_1/lout')

wire n6390;
// (21, 2, 'lutff_5/lout')

wire n6391;
// (11, 5, 'lutff_4/lout')

wire n6392;
// (8, 17, 'lutff_5/out')

wire n6393;
// (8, 17, 'lutff_5/lout')

wire n6394;
// (12, 1, 'lutff_2/out')

wire n6395;
// (12, 1, 'lutff_2/lout')

wire n6396;
// (5, 11, 'lutff_0/out')

wire n6397;
// (5, 11, 'lutff_0/lout')

wire n6398;
// (5, 11, 'carry_in_mux')

// Carry-In for (5 11)
assign n6398 = 1;

wire n6399;
// (12, 4, 'lutff_7/lout')

wire n6400;
// (15, 8, 'lutff_7/lout')

wire n6401;
// (22, 7, 'lutff_7/lout')

wire n6402;
// (9, 22, 'lutff_1/lout')

wire n6403;
// (21, 3, 'lutff_6/lout')

wire n6404;
// (16, 21, 'lutff_1/lout')

wire n6405;
// (7, 14, 'lutff_4/lout')

wire n6406;
// (8, 10, 'lutff_2/lout')

wire n6407;
// (1, 20, 'lutff_0/out')

wire n6408;
// (1, 20, 'lutff_0/lout')

wire n6409;
// (1, 20, 'carry_in_mux')

// Carry-In for (1 20)
assign n6409 = 1;

wire n6410;
// (5, 3, 'lutff_1/lout')

wire n6411;
// (17, 4, 'lutff_2/lout')

wire n6412;
// (5, 6, 'lutff_6/lout')

wire n6413;
// (1, 21, 'lutff_1/lout')

wire n6414;
// (16, 13, 'lutff_2/lout')

wire n6415;
// (4, 2, 'lutff_5/lout')

wire n6416;
// (14, 5, 'lutff_5/lout')

wire n6417;
// (16, 16, 'lutff_7/lout')

wire n6418;
// (7, 15, 'lutff_4/out')

wire n6419;
// (7, 15, 'lutff_4/lout')

wire n6420;
// (7, 7, 'lutff_0/lout')

wire n6421;
// (5, 7, 'lutff_7/lout')

wire n6422;
// (9, 19, 'lutff_4/lout')

wire n6423;
// (4, 3, 'lutff_6/lout')

wire n6424;
// (16, 9, 'lutff_4/lout')

wire n6425;
// (17, 5, 'lutff_2/lout')

wire n6426;
// (3, 16, 'lutff_0/lout')

wire n6427;
// (18, 18, 'lutff_1/lout')

wire n6428;
// (20, 12, 'lutff_7/lout')

wire n6429;
// (10, 15, 'lutff_6/lout')

wire n6430;
// (10, 7, 'lutff_2/lout')

wire n6431;
// (13, 22, 'lutff_6/lout')

wire n6432;
// (22, 21, 'lutff_4/lout')

wire n6433;
// (2, 21, 'lutff_3/lout')

wire n6434;
// (13, 14, 'lutff_2/lout')

wire n6435;
// (22, 13, 'lutff_0/lout')

wire n6436;
// (3, 17, 'lutff_1/lout')

wire n6437;
// (16, 1, 'lutff_5/lout')

wire n6438;
// (9, 11, 'lutff_4/lout')

wire n6439;
// (18, 10, 'lutff_2/lout')

wire n6440;
// (9, 3, 'lutff_0/lout')

wire n6441;
// (12, 11, 'lutff_1/lout')

wire n6442;
// (7, 3, 'lutff_7/lout')

wire n6443;
// (13, 15, 'lutff_3/lout')

wire n6444;
// (11, 20, 'lutff_1/lout')

wire n6445;
// (10, 8, 'lutff_2/lout')

wire n6446;
// (9, 4, 'lutff_1/lout')

wire n6447;
// (22, 22, 'lutff_4/lout')

wire n6448;
// (22, 14, 'lutff_0/out')

wire n6449;
// (22, 14, 'lutff_0/lout')

wire n6450;
// (22, 14, 'carry_in_mux')

// Carry-In for (22 14)
assign n6450 = 1;

wire n6451;
// (21, 18, 'lutff_3/lout')

wire n6452;
// (9, 7, 'lutff_6/lout')

wire n6453;
// (12, 3, 'lutff_2/out')

wire n6454;
// (12, 3, 'lutff_2/lout')

wire n6455;
// (5, 13, 'lutff_0/lout')

wire n6456;
// (4, 17, 'lutff_3/lout')

wire n6457;
// (11, 16, 'lutff_3/lout')

wire n6458;
// (2, 9, 'lutff_6/lout')

wire n6459;
// (13, 2, 'lutff_5/lout')

wire n6460;
// (3, 5, 'lutff_4/lout')

wire n6461;
// (11, 15, 'lutff_7/lout')

wire n6462;
// (15, 11, 'lutff_2/lout')

wire n6463;
// (2, 6, 'lutff_0/out')

wire n6464;
// (2, 6, 'lutff_0/lout')

wire n6465;
// (2, 6, 'carry_in_mux')

// Carry-In for (2 6)
assign n6465 = 1;

wire n6466;
// (5, 14, 'lutff_1/lout')

wire n6467;
// (14, 20, 'lutff_2/lout')

wire n6468;
// (8, 21, 'lutff_1/lout')

wire n6469;
// (13, 3, 'lutff_6/lout')

wire n6470;
// (22, 9, 'lutff_6/lout')

wire n6471;
// (21, 5, 'lutff_5/lout')

wire n6472;
// (17, 20, 'lutff_0/lout')

wire n6473;
// (11, 8, 'lutff_4/lout')

wire n6474;
// (15, 12, 'lutff_3/lout')

wire n6475;
// (23, 14, 'lutff_2/lout')

wire n6476;
// (4, 18, 'lutff_3/out')

wire n6477;
// (4, 18, 'lutff_3/lout')

wire n6478;
// (2, 10, 'lutff_6/lout')

wire n6479;
// (22, 2, 'lutff_3/lout')

wire n6480;
// (2, 2, 'lutff_2/lout')

wire n6481;
// (21, 6, 'lutff_6/lout')

wire n6482;
// (11, 1, 'lutff_1/out')

wire n6483;
// (11, 1, 'lutff_1/lout')

wire n6484;
// (8, 13, 'lutff_2/lout')

wire n6485;
// (5, 9, 'lutff_7/lout')

wire n6486;
// (4, 5, 'lutff_6/lout')

wire n6487;
// (11, 4, 'lutff_6/lout')

wire n6488;
// (7, 18, 'lutff_5/out')

wire n6489;
// (7, 18, 'lutff_5/lout')

wire n6490;
// (17, 7, 'lutff_2/out')

wire n6491;
// (17, 7, 'lutff_2/lout')

wire n6492;
// (7, 10, 'lutff_1/lout')

wire n6493;
// (9, 21, 'lutff_3/lout')

wire n6494;
// (20, 20, 'lutff_1/lout')

wire n6495;
// (14, 8, 'lutff_5/lout')

wire n6496;
// (8, 9, 'lutff_4/lout')

wire n6497;
// (11, 30, 'lutff_0/lout')

wire n6498;
// (17, 8, 'lutff_3/lout')

wire n6499;
// (10, 18, 'lutff_1/out')

wire n6500;
// (10, 18, 'lutff_1/lout')

wire n6501;
// (9, 22, 'lutff_4/lout')

wire n6502;
// (23, 2, 'lutff_5/lout')

wire n6503;
// (4, 6, 'lutff_6/lout')

wire n6504;
// (14, 1, 'lutff_2/lout')

wire n6505;
// (8, 2, 'lutff_1/lout')

wire n6506;
// (16, 12, 'lutff_4/lout')

wire n6507;
// (16, 4, 'lutff_0/lout')

wire n6508;
// (13, 17, 'lutff_3/out')

wire n6509;
// (13, 17, 'lutff_3/lout')

wire n6510;
// (14, 4, 'lutff_7/lout')

wire n6511;
// (20, 16, 'lutff_3/lout')

wire n6512;
// (8, 1, 'lutff_5/lout')

wire n6513;
// (1, 19, 'lutff_7/lout')

wire n6514;
// (18, 21, 'lutff_1/lout')

wire n6515;
// (1, 11, 'lutff_3/lout')

wire n6516;
// (20, 15, 'lutff_7/lout')

wire n6517;
// (17, 4, 'lutff_5/lout')

wire n6518;
// (10, 10, 'lutff_2/lout')

wire n6519;
// (9, 6, 'lutff_1/lout')

wire n6520;
// (16, 5, 'lutff_1/lout')

wire n6521;
// (10, 13, 'lutff_7/lout')

wire n6522;
// (3, 20, 'lutff_1/lout')

wire n6523;
// (9, 9, 'lutff_6/lout')

wire n6524;
// (1, 12, 'lutff_4/lout')

wire n6525;
// (1, 4, 'lutff_0/lout')

wire n6526;
// (20, 8, 'lutff_4/lout')

wire n6527;
// (12, 22, 'lutff_5/lout')

wire n6528;
// (18, 13, 'lutff_2/lout')

wire n6529;
// (12, 14, 'lutff_1/lout')

wire n6530;
// (22, 17, 'lutff_1/lout')

wire n6531;
// (2, 17, 'lutff_0/out')

wire n6532;
// (2, 17, 'lutff_0/lout')

wire n6533;
// (2, 17, 'carry_in_mux')

// Carry-In for (2 17)
assign n6533 = 1;

wire n6534;
// (10, 6, 'lutff_4/lout')

wire n6535;
// (9, 10, 'lutff_7/lout')

wire n6536;
// (9, 2, 'lutff_3/lout')

wire n6537;
// (22, 20, 'lutff_6/lout')

wire n6538;
// (3, 16, 'lutff_3/lout')

wire n6539;
// (21, 16, 'lutff_5/lout')

wire n6540;
// (20, 1, 'lutff_1/out')

wire n6541;
// (20, 1, 'lutff_1/lout')

wire n6542;
// (3, 15, 'lutff_7/lout')

wire n6543;
// (10, 7, 'lutff_5/lout')

wire n6544;
// (18, 9, 'lutff_4/lout')

wire n6545;
// (22, 21, 'lutff_7/lout')

wire n6546;
// (22, 13, 'lutff_3/lout')

wire n6547;
// (4, 20, 'lutff_3/lout')

wire n6548;
// (2, 12, 'lutff_6/lout')

wire n6549;
// (13, 5, 'lutff_5/lout')

wire n6550;
// (3, 8, 'lutff_4/lout')

wire n6551;
// (18, 10, 'lutff_5/lout')

wire n6552;
// (18, 2, 'lutff_1/lout')

wire n6553;
// (15, 14, 'lutff_2/lout')

wire n6554;
// (5, 17, 'lutff_1/lout')

wire n6555;
// (4, 13, 'lutff_0/out')

wire n6556;
// (4, 13, 'lutff_0/lout')

wire n6557;
// (4, 13, 'carry_in_mux')

// Carry-In for (4 13)
assign n6557 = 1;

wire n6558;
// (2, 13, 'lutff_7/lout')

wire n6559;
// (12, 2, 'lutff_4/lout')

wire n6560;
// (13, 6, 'lutff_6/lout')

wire n6561;
// (2, 5, 'lutff_3/lout')

wire n6562;
// (3, 1, 'lutff_1/lout')

wire n6563;
// (4, 16, 'lutff_5/lout')

wire n6564;
// (11, 11, 'lutff_4/lout')

wire n6565;
// (14, 19, 'lutff_5/lout')

wire n6566;
// (11, 3, 'lutff_0/lout')

wire n6567;
// (14, 11, 'lutff_1/lout')

wire n6568;
// (15, 15, 'lutff_3/lout')

wire n6569;
// (3, 4, 'lutff_6/lout')

wire n6570;
// (7, 21, 'lutff_0/out')

wire n6571;
// (7, 21, 'lutff_0/lout')

wire n6572;
// (12, 3, 'lutff_5/out')

wire n6573;
// (12, 3, 'lutff_5/lout')

wire n6574;
// (22, 5, 'lutff_3/lout')

wire n6575;
// (5, 13, 'lutff_3/lout')

wire n6576;
// (4, 17, 'lutff_6/lout')

wire n6577;
// (4, 9, 'lutff_2/lout')

wire n6578;
// (17, 19, 'lutff_2/lout')

wire n6579;
// (11, 7, 'lutff_6/lout')

wire n6580;
// (17, 18, 'lutff_6/lout')

wire n6581;
// (7, 13, 'lutff_1/lout')

wire n6582;
// (14, 12, 'lutff_1/lout')

wire n6583;
// (5, 5, 'lutff_4/lout')

wire n6584;
// (4, 1, 'lutff_3/lout')

wire n6585;
// (8, 12, 'lutff_4/lout')

wire n6586;
// (8, 4, 'lutff_0/lout')

wire n6587;
// (16, 15, 'lutff_5/lout')

wire n6588;
// (23, 14, 'lutff_5/lout')

wire n6589;
// (20, 18, 'lutff_2/lout')

wire n6590;
// (15, 3, 'lutff_6/lout')

wire n6591;
// (9, 17, 'lutff_0/out')

wire n6592;
// (9, 17, 'lutff_0/lout')

wire n6593;
// (7, 17, 'lutff_7/lout')

wire n6594;
// (7, 9, 'lutff_3/lout')

wire n6595;
// (8, 13, 'lutff_5/lout')

wire n6596;
// (8, 5, 'lutff_1/lout')

wire n6597;
// (14, 7, 'lutff_7/lout')

wire n6598;
// (17, 7, 'lutff_5/lout')

wire n6599;
// (3, 18, 'lutff_3/lout')

wire n6600;
// (7, 2, 'lutff_0/lout')

wire n6601;
// (9, 21, 'lutff_6/lout')

wire n6602;
// (16, 8, 'lutff_1/lout')

wire n6603;
// (13, 13, 'lutff_0/lout')

wire n6604;
// (1, 7, 'lutff_0/out')

wire n6605;
// (1, 7, 'lutff_0/lout')

wire n6606;
// (1, 7, 'carry_in_mux')

// Carry-In for (1 7)
assign n6606 = 1;

wire n6607;
// (13, 16, 'lutff_5/lout')

wire n6608;
// (3, 19, 'lutff_4/lout')

wire n6609;
// (12, 17, 'lutff_1/lout')

wire n6610;
// (20, 6, 'lutff_5/lout')

wire n6611;
// (2, 20, 'lutff_0/lout')

wire n6612;
// (10, 9, 'lutff_4/lout')

wire n6613;
// (9, 13, 'lutff_7/lout')

wire n6614;
// (9, 5, 'lutff_3/lout')

wire n6615;
// (13, 17, 'lutff_6/lout')

wire n6616;
// (1, 8, 'lutff_1/out')

wire n6617;
// (1, 8, 'lutff_1/lout')

wire n6618;
// (22, 23, 'lutff_6/lout')

wire n6619;
// (1, 11, 'lutff_6/lout')

wire n6620;
// (12, 18, 'lutff_2/lout')

wire n6621;
// (20, 7, 'lutff_6/lout')

wire n6622;
// (10, 10, 'lutff_5/lout')

wire n6623;
// (10, 2, 'lutff_1/lout')

wire n6624;
// (12, 21, 'lutff_7/lout')

wire n6625;
// (9, 6, 'lutff_4/lout')

wire n6626;
// (18, 12, 'lutff_4/lout')

wire n6627;
// (18, 4, 'lutff_0/lout')

wire n6628;
// (22, 16, 'lutff_3/lout')

wire n6629;
// (13, 9, 'lutff_1/lout')

wire n6630;
// (21, 20, 'lutff_6/lout')

wire n6631;
// (21, 12, 'lutff_2/lout')

wire n6632;
// (3, 3, 'lutff_0/lout')

wire n6633;
// (18, 13, 'lutff_5/lout')

wire n6634;
// (1, 3, 'lutff_7/lout')

wire n6635;
// (18, 5, 'lutff_1/lout')

wire n6636;
// (5, 20, 'lutff_1/lout')

wire n6637;
// (17, 21, 'lutff_2/lout')

wire n6638;
// (12, 5, 'lutff_4/lout')

// RAM TILE 19 5
SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_19_5 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, n2470, n2469, n2468, n2467, n2466, n2465, n2481}),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, n2682, n2681, n2680, n2679, n2678, n2677, n2621}),
  .MASK({n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363, n2363}),
  .WDATA({n2190, n2335, n2337, n2336, n2338, n2334, n2458, n2443, n2339, n2444, n2617, n2460, n2464, n2446, n2445, n2171}),
  .RDATA({open_0, open_1, open_2, open_3, open_4, open_5, open_6, open_7, n2604, n2605, n2606, n2607, n2608, n2609, n2482, n2610}),
  .WE(n8),
  .WCLKE(n2683),
  .WCLK(io_13_31_1),
  .RE(n8),
  .RCLKE(n2623),
  .RCLK(io_13_31_1)
);

// RAM TILE 19 7
SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_19_7 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, n2470, n2469, n2468, n2467, n2466, n2465, n2481}),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, n2682, n2681, n2680, n2679, n2678, n2677, n2621}),
  .MASK({n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n2363, n2363, n2363, n2363}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n2463, n2462, n2461, n2459}),
  .RDATA({open_16, open_17, open_18, open_19, open_20, open_21, open_22, open_23, open_24, open_25, open_26, open_27, n2618, n2619, n2620, n2616}),
  .WE(n8),
  .WCLKE(n2683),
  .WCLK(io_13_31_1),
  .RE(n8),
  .RCLKE(n2623),
  .RCLK(io_13_31_1)
);

// RAM TILE 19 9
SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_19_9 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, n2388, n2256, n2255, n2387, n2385, n2386, n2257}),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, n2393, n2267, n2265, n2392, n2391, n2266, n2394}),
  .MASK({n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n2664, n2664, n2664, n2664}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n2249, n2398, n2264}),
  .RDATA({open_32, open_33, open_34, open_35, open_36, open_37, open_38, open_39, open_40, open_41, open_42, open_43, n2625, n2626, n2627, n2628}),
  .WE(n8),
  .WCLKE(n2133),
  .WCLK(io_13_31_1),
  .RE(n8),
  .RCLKE(n2275),
  .RCLK(io_13_31_1)
);

// RAM TILE 19 11
SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_19_11 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, n2388, n2256, n2255, n2387, n2385, n2386, n2257}),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, n2393, n2267, n2265, n2392, n2391, n2266, n2394}),
  .MASK({n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .RDATA({n2632, n2248, n2633, n2634, n2635, n2636, n2637, n2638, n2642, n2643, n2389, n2640, n2644, n2645, n2641, n2646}),
  .WE(n8),
  .WCLKE(n2133),
  .WCLK(io_13_31_1),
  .RE(n8),
  .RCLKE(n2275),
  .RCLK(io_13_31_1)
);

// RAM TILE 19 13
SB_RAM40_4K #(
  .READ_MODE(0),
  .WRITE_MODE(0),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_19_13 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, n2388, n2256, n2255, n2387, n2385, n2386, n2257}),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, n2393, n2267, n2265, n2392, n2391, n2266, n2394}),
  .MASK({n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664, n2664}),
  .WDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n2401, n2258, n2399, n2261, n2260, n2263, n2262, n2259}),
  .RDATA({n2648, n2649, n2647, n2650, n2651, n2652, n2653, n2654, n2657, n2659, n2660, n2655, n2661, n2662, n2656, n2658}),
  .WE(n8),
  .WCLKE(n2133),
  .WCLK(io_13_31_1),
  .RE(n8),
  .RCLKE(n2275),
  .RCLK(io_13_31_1)
);

// RAM TILE 19 15
SB_RAM40_4K #(
  .READ_MODE(1),
  .WRITE_MODE(1),
  .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) ram40_19_15 (
  .WADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n1651, n1650, n1780, n1812, n1978, n1980}),
  .RADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n1798, n1797, n1792, n1796, n1795, n1968}),
  .MASK({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .WDATA({1'b0, n1955, 1'b0, n1954, 1'b0, n1760, 1'b0, n1949, 1'b0, n1964, 1'b0, n1958, 1'b0, n1953, 1'b0, n1786}),
  .RDATA({open_64, n1625, open_65, n1616, open_66, n1782, open_67, n1615, open_68, n1791, open_70, n1626, open_72, n1627, open_74, n1204}),
  .WE(n8),
  .WCLKE(n1981),
  .WCLK(io_13_31_1),
  .RE(n8),
  .RCLKE(n8),
  .RCLK(io_13_31_1)
);

assign n3286 = /* LUT   13  1  2 */ 1'b0;
assign n3305 = /* LUT    8 15  5 */ 1'b0;
assign n3313 = /* LUT   16 19  1 */ 1'b0;
assign n3317 = /* LUT   16 18  5 */ 1'b0;
assign n3321 = /* LUT    9 20  0 */ 1'b0;
assign n3325 = /* LUT    7 20  7 */ 1'b0;
assign n3338 = /* LUT    9 16  2 */ 1'b0;
assign n3346 = /* LUT    3 14  0 */ 1'b0;
assign n3350 = /* LUT    1  6  3 */ 1'b0;
assign n3374 = /* LUT    8 18  0 */ 1'b0;
assign n3380 = /* LUT   12  1  1 */ 1'b0;
assign n3385 = /* LUT    8 19  1 */ 1'b0;
assign n3392 = /* LUT   15 17  5 */ 1'b0;
assign n3400 = /* LUT    1 21  0 */ 1'b0;
assign n3406 = /* LUT    7 15  3 */ 1'b0;
assign n3411 = /* LUT    8  7  4 */ 1'b0;
assign n3418 = /* LUT    7  8  0 */ 1'b0;
assign n3428 = /* LUT   17  6  2 */ 1'b0;
assign n3431 = /* LUT    3 17  0 */ 1'b0;
assign n3453 = /* LUT   12 12  0 */ 1'b0;
assign n3456 = /* LUT   22 15  0 */ 1'b0;
assign n3476 = /* LUT   11  1  0 */ 1'b0;
assign n3489 = /* LUT    8 17  7 */ 1'b0;
assign n3492 = /* LUT   10 18  0 */ 1'b0;
assign n3515 = /* LUT    7 15  6 */ 1'b0;
assign n3524 = /* LUT   20  1  0 */ 1'b0;
assign n3548 = /* LUT   15 15  2 */ 1'b0;
assign n3551 = /* LUT   15 18  7 */ 1'b0;
assign n3553 = /* LUT   12  3  4 */ 1'b0;
assign n3560 = /* LUT   17 19  1 */ 1'b0;
assign n3582 = /* LUT   11  1  3 */ 1'b0;
assign n3587 = /* LUT    9 18  0 */ 1'b0;
assign n3590 = /* LUT    7 18  7 */ 1'b0;
assign n3592 = /* LUT   17  7  4 */ 1'b0;
assign n3602 = /* LUT   10 18  3 */ 1'b0;
assign n3610 = /* LUT    1  8  0 */ 1'b0;
assign n3613 = /* LUT   13 17  5 */ 1'b0;
assign n3617 = /* LUT   20  7  5 */ 1'b0;
assign n3639 = /* LUT   14 23  0 */ 1'b0;
assign n3647 = /* LUT   21 13  1 */ 1'b0;
assign n3654 = /* LUT    4 12  1 */ 1'b0;
assign n3658 = /* LUT    8 16  0 */ 1'b0;
assign n3666 = /* LUT    4 13  2 */ 1'b0;
assign n3686 = /* LUT   17 11  0 */ 1'b0;
assign n3693 = /* LUT    9 16  1 */ 1'b0;
assign n3741 = /* LUT    8 19  0 */ 1'b0;
assign n3751 = /* LUT   13  1  4 */ 1'b0;
assign n3764 = /* LUT   17 14  0 */ 1'b0;
assign n3768 = /* LUT    8 15  7 */ 1'b0;
assign n3770 = /* LUT    8  7  3 */ 1'b0;
assign n3774 = /* LUT   13 23  0 */ 1'b0;
assign n3777 = /* LUT   16 18  7 */ 1'b0;
assign n3791 = /* LUT   20 14  1 */ 1'b0;
assign n3797 = /* LUT    9 16  4 */ 1'b0;
assign n3803 = /* LUT    3 14  2 */ 1'b0;
assign n3822 = /* LUT   21  7  0 */ 1'b0;
assign n3835 = /* LUT   18  1  0 */ 1'b0;
assign n3840 = /* LUT   12  1  3 */ 1'b0;
assign n3858 = /* LUT    7 15  5 */ 1'b0;
assign n3893 = /* LUT   22 15  2 */ 1'b0;
assign n3899 = /* LUT    2  6  1 */ 1'b0;
assign n3920 = /* LUT   11  1  2 */ 1'b0;
assign n3930 = /* LUT    7 18  6 */ 1'b0;
assign n3939 = /* LUT   10 18  2 */ 1'b0;
assign n3964 = /* LUT    2 17  1 */ 1'b0;
assign n3974 = /* LUT   21 13  0 */ 1'b0;
assign n3978 = /* LUT    4 21  0 */ 1'b0;
assign n4001 = /* LUT   12  3  6 */ 1'b0;
assign n4008 = /* LUT   17 19  3 */ 1'b0;
assign n4018 = /* LUT    5  6  0 */ 1'b0;
assign n4030 = /* LUT    9 18  2 */ 1'b0;
assign n4043 = /* LUT   10 18  5 */ 1'b0;
assign n4049 = /* LUT    1  8  2 */ 1'b0;
assign n4051 = /* LUT   13 17  7 */ 1'b0;
assign n4056 = /* LUT   20  7  7 */ 1'b0;
assign n4075 = /* LUT    2  9  0 */ 1'b0;
assign n4081 = /* LUT    8 20  0 */ 1'b0;
assign n4101 = /* LUT    4 13  4 */ 1'b0;
assign n4115 = /* LUT   20 14  0 */ 1'b0;
assign n4122 = /* LUT    9 16  3 */ 1'b0;
assign n4171 = /* LUT    8 19  2 */ 1'b0;
assign n4182 = /* LUT    4  8  0 */ 1'b0;
assign n4187 = /* LUT   13  1  6 */ 1'b0;
assign n4190 = /* LUT   17 18  0 */ 1'b0;
assign n4197 = /* LUT    7 16  0 */ 1'b0;
assign n4203 = /* LUT    8  7  5 */ 1'b0;
assign n4218 = /* LUT    9 12  0 */ 1'b0;
assign n4231 = /* LUT    9 16  6 */ 1'b0;
assign n4276 = /* LUT    7 19  0 */ 1'b0;
assign n4278 = /* LUT   12  1  5 */ 1'b0;
assign n4295 = /* LUT    1 13  0 */ 1'b0;
assign n4301 = /* LUT    7 15  7 */ 1'b0;
assign n4313 = /* LUT    3  9  0 */ 1'b0;
assign n4359 = /* LUT   11  1  4 */ 1'b0;
assign n4367 = /* LUT    9 18  1 */ 1'b0;
assign n4372 = /* LUT    1 16  0 */ 1'b0;
assign n4379 = /* LUT   10 18  4 */ 1'b0;
assign n4384 = /* LUT    1 17  1 */ 1'b0;
assign n4407 = /* LUT    3 13  1 */ 1'b0;
assign n4427 = /* LUT    4 13  3 */ 1'b0;
assign n4439 = /* LUT    8 17  1 */ 1'b0;
assign n4447 = /* LUT   17 19  5 */ 1'b0;
assign n4454 = /* LUT    1 19  0 */ 1'b0;
assign n4469 = /* LUT    9 18  4 */ 1'b0;
assign n4496 = /* LUT   15 18  1 */ 1'b0;
assign n4507 = /* LUT   13  1  5 */ 1'b0;
assign n4541 = /* LUT   23  2  1 */ 1'b0;
assign n4550 = /* LUT    9 16  5 */ 1'b0;
assign n4556 = /* LUT   12 21  0 */ 1'b0;
assign n4595 = /* LUT   12  1  4 */ 1'b0;
assign n4603 = /* LUT    8 19  4 */ 1'b0;
assign n4608 = /* LUT    7 20  0 */ 1'b0;
assign n4675 = /* LUT    4 18  5 */ 1'b0;
assign n4683 = /* LUT    8 15  1 */ 1'b0;
assign n4694 = /* LUT   12  1  7 */ 1'b0;
assign n4701 = /* LUT    1 17  0 */ 1'b0;
assign n4729 = /* LUT    3 13  0 */ 1'b0;
assign n4738 = /* LUT    4 21  1 */ 1'b0;
assign n4752 = /* LUT   15 16  1 */ 1'b0;
assign n4756 = /* LUT   22 14  5 */ 1'b0;
assign n4762 = /* LUT    8 17  0 */ 1'b0;
assign n4788 = /* LUT   11  1  6 */ 1'b0;
assign n4792 = /* LUT    9 18  3 */ 1'b0;
assign n4801 = /* LUT   10 18  6 */ 1'b0;
assign n4816 = /* LUT   15 18  0 */ 1'b0;
assign n4824 = /* LUT    3 13  3 */ 1'b0;
assign n4830 = /* LUT   15 19  1 */ 1'b0;
assign n4838 = /* LUT    4 21  4 */ 1'b0;
assign n4850 = /* LUT   16 19  3 */ 1'b0;
assign n4855 = /* LUT    7 18  0 */ 1'b0;
assign n4862 = /* LUT    8 17  3 */ 1'b0;
assign n4867 = /* LUT   17 19  7 */ 1'b0;
assign n4870 = /* LUT   23  2  0 */ 1'b0;
assign n4881 = /* LUT   23  3  1 */ 1'b0;
assign n4891 = /* LUT   12 22  0 */ 1'b0;
assign n4896 = /* LUT    9 18  6 */ 1'b0;
assign n4913 = /* LUT   21  8  1 */ 1'b0;
assign n4924 = /* LUT   14 19  0 */ 1'b0;
assign n4932 = /* LUT   15 18  3 */ 1'b0;
assign n4934 = /* LUT    8 19  3 */ 1'b0;
assign n4936 = /* LUT   12  3  0 */ 1'b0;
assign n4945 = /* LUT   13  1  7 */ 1'b0;
assign n4965 = /* LUT   17  7  0 */ 1'b0;
assign n4968 = /* LUT   17  6  4 */ 1'b0;
assign n4980 = /* LUT   20  6  0 */ 1'b0;
assign n4986 = /* LUT   13 17  1 */ 1'b0;
assign n4990 = /* LUT    9 16  7 */ 1'b0;
assign n4993 = /* LUT   20  7  1 */ 1'b0;
assign n5020 = /* LUT   21  7  3 */ 1'b0;
assign n5034 = /* LUT    8 15  0 */ 1'b0;
assign n5041 = /* LUT   12  1  6 */ 1'b0;
assign n5045 = /* LUT   16 18  0 */ 1'b0;
assign n5050 = /* LUT    8 19  6 */ 1'b0;
assign n5054 = /* LUT    7 20  2 */ 1'b0;
assign n5063 = /* LUT   17 10  0 */ 1'b0;
assign n5072 = /* LUT   13 19  0 */ 1'b0;
assign n5079 = /* LUT   13 20  1 */ 1'b0;
assign n5097 = /* LUT   15 16  0 */ 1'b0;
assign n5116 = /* LUT   21  3  0 */ 1'b0;
assign n5127 = /* LUT    4 18  7 */ 1'b0;
assign n5134 = /* LUT   11  1  5 */ 1'b0;
assign n5141 = /* LUT    8 15  3 */ 1'b0;
assign n5144 = /* LUT   17 13  0 */ 1'b0;
assign n5155 = /* LUT   16 18  3 */ 1'b0;
assign n5179 = /* LUT    3 13  2 */ 1'b0;
assign n5212 = /* LUT    8 17  2 */ 1'b0;
assign n5239 = /* LUT    9 18  5 */ 1'b0;
assign n5250 = /* LUT    2 21  0 */ 1'b0;
assign n5254 = /* LUT   20  5  1 */ 1'b0;
assign n5273 = /* LUT    3 13  5 */ 1'b0;
assign n5279 = /* LUT   15 19  3 */ 1'b0;
assign n5300 = /* LUT    7 18  2 */ 1'b0;
assign n5315 = /* LUT   13 17  0 */ 1'b0;
assign n5322 = /* LUT   23  3  3 */ 1'b0;
assign n5326 = /* LUT   20  7  0 */ 1'b0;
assign n5337 = /* LUT   20  8  1 */ 1'b0;
assign n5363 = /* LUT   21  8  3 */ 1'b0;
assign n5373 = /* LUT   11 11  1 */ 1'b0;
assign n5377 = /* LUT   15 15  0 */ 1'b0;
assign n5382 = /* LUT   15 18  5 */ 1'b0;
assign n5384 = /* LUT    8 19  5 */ 1'b0;
assign n5387 = /* LUT    7 20  1 */ 1'b0;
assign n5403 = /* LUT    7  9  0 */ 1'b0;
assign n5407 = /* LUT   13 20  0 */ 1'b0;
assign n5412 = /* LUT    3 18  0 */ 1'b0;
assign n5415 = /* LUT   17  6  6 */ 1'b0;
assign n5430 = /* LUT   20  7  3 */ 1'b0;
assign n5447 = /* LUT    2  8  0 */ 1'b0;
assign n5453 = /* LUT   21  7  5 */ 1'b0;
assign n5466 = /* LUT    8 15  2 */ 1'b0;
assign n5481 = /* LUT    7 20  4 */ 1'b0;
assign n5503 = /* LUT    1  6  0 */ 1'b0;
assign n5560 = /* LUT   11  1  7 */ 1'b0;
assign n5562 = /* LUT    7 15  0 */ 1'b0;
assign n5567 = /* LUT    9 19  0 */ 1'b0;
assign n5571 = /* LUT    8  7  1 */ 1'b0;
assign n5584 = /* LUT   10 18  7 */ 1'b0;
assign n5590 = /* LUT   20  5  0 */ 1'b0;
assign n5611 = /* LUT    3 13  4 */ 1'b0;
assign n5642 = /* LUT    7 18  1 */ 1'b0;
assign n5648 = /* LUT    8 17  4 */ 1'b0;
assign n5650 = /* LUT    8  9  0 */ 1'b0;
assign n5655 = /* LUT    9 22  0 */ 1'b0;
assign n5680 = /* LUT    9 18  7 */ 1'b0;
assign n5694 = /* LUT    3  8  0 */ 1'b0;
assign n5704 = /* LUT   11 11  0 */ 1'b0;
assign n5712 = /* LUT   12  3  1 */ 1'b0;
assign n5747 = /* LUT    7 18  4 */ 1'b0;
assign n5756 = /* LUT    3 19  0 */ 1'b0;
assign n5760 = /* LUT   23  2  4 */ 1'b0;
assign n5778 = /* LUT   20  8  3 */ 1'b0;
assign n5783 = /* LUT   12 14  0 */ 1'b0;
assign n5813 = /* LUT   11 11  3 */ 1'b0;
assign n5818 = /* LUT    8 19  7 */ 1'b0;
assign n5824 = /* LUT    7 20  3 */ 1'b0;
assign n5876 = /* LUT   21  3  1 */ 1'b0;
assign n5888 = /* LUT   13  1  1 */ 1'b0;
assign n5895 = /* LUT   21  7  7 */ 1'b0;
assign n5904 = /* LUT    8 15  4 */ 1'b0;
assign n5906 = /* LUT    8  7  0 */ 1'b0;
assign n5923 = /* LUT    7 20  6 */ 1'b0;
assign n5944 = /* LUT    1  6  2 */ 1'b0;
assign n5971 = /* LUT   12  1  0 */ 1'b0;
assign n5995 = /* LUT   23 12  0 */ 1'b0;
assign n5998 = /* LUT    7 15  2 */ 1'b0;
assign n6049 = /* LUT    4 18  1 */ 1'b0;
assign n6060 = /* LUT    7 18  3 */ 1'b0;
assign n6065 = /* LUT    8 17  6 */ 1'b0;
assign n6122 = /* LUT   15 15  1 */ 1'b0;
assign n6127 = /* LUT   12  3  3 */ 1'b0;
assign n6135 = /* LUT   17 19  0 */ 1'b0;
assign n6166 = /* LUT   23  2  6 */ 1'b0;
assign n6193 = /* LUT    2  8  1 */ 1'b0;
assign n6195 = /* LUT   13  1  0 */ 1'b0;
assign n6198 = /* LUT    4 19  3 */ 1'b0;
assign n6201 = /* LUT   18  6  0 */ 1'b0;
assign n6211 = /* LUT    4 12  0 */ 1'b0;
assign n6224 = /* LUT    4 13  1 */ 1'b0;
assign n6231 = /* LUT    7 20  5 */ 1'b0;
assign n6243 = /* LUT    9 16  0 */ 1'b0;
assign n6257 = /* LUT    1  6  1 */ 1'b0;
assign n6267 = /* LUT    2 19  0 */ 1'b0;
assign n6306 = /* LUT   13  1  3 */ 1'b0;
assign n6315 = /* LUT    7 15  1 */ 1'b0;
assign n6323 = /* LUT    8 15  6 */ 1'b0;
assign n6325 = /* LUT    8  7  2 */ 1'b0;
assign n6335 = /* LUT   17  6  0 */ 1'b0;
assign n6339 = /* LUT    9 20  1 */ 1'b0;
assign n6345 = /* LUT   13 15  0 */ 1'b0;
assign n6357 = /* LUT    3 14  1 */ 1'b0;
assign n6360 = /* LUT    1  6  4 */ 1'b0;
assign n6374 = /* LUT    4 18  0 */ 1'b0;
assign n6393 = /* LUT    8 17  5 */ 1'b0;
assign n6395 = /* LUT   12  1  2 */ 1'b0;
assign n6397 = /* LUT    5 11  0 */ 1'b0;
assign n6408 = /* LUT    1 20  0 */ 1'b0;
assign n6419 = /* LUT    7 15  4 */ 1'b0;
assign n6449 = /* LUT   22 14  0 */ 1'b0;
assign n6454 = /* LUT   12  3  2 */ 1'b0;
assign n6464 = /* LUT    2  6  0 */ 1'b0;
assign n6477 = /* LUT    4 18  3 */ 1'b0;
assign n6483 = /* LUT   11  1  1 */ 1'b0;
assign n6489 = /* LUT    7 18  5 */ 1'b0;
assign n6491 = /* LUT   17  7  2 */ 1'b0;
assign n6500 = /* LUT   10 18  1 */ 1'b0;
assign n6509 = /* LUT   13 17  3 */ 1'b0;
assign n6532 = /* LUT    2 17  0 */ 1'b0;
assign n6541 = /* LUT   20  1  1 */ 1'b0;
assign n6556 = /* LUT    4 13  0 */ 1'b0;
assign n6571 = /* LUT    7 21  0 */ 1'b0;
assign n6573 = /* LUT   12  3  5 */ 1'b0;
assign n6592 = /* LUT    9 17  0 */ 1'b0;
assign n6605 = /* LUT    1  7  0 */ 1'b0;
assign n6617 = /* LUT    1  8  1 */ 1'b0;
assign n3287 = /* LUT    2  8  3 */ (n412 ? (n227 ? 1'b0 : n240) : (n227 ? n240 : 1'b0));
assign n3288 = /* LUT    4 19  5 */ (n249 ? n783 : 1'b0);
assign n3289 = /* LUT   14 22  5 */ (n1846 ? 1'b0 : (n1528 ? 1'b0 : n2027));
assign n3290 = /* LUT   14 14  1 */ (n1963 ? (n1770 ? n1926 : 1'b1) : (n1770 ? n1926 : !n2118));
assign n3291 = /* LUT    3  7  6 */ n15;
assign n3292 = /* LUT   11 10  7 */ (n1459 ? n1349 : 1'b0);
assign n3293 = /* LUT   12  6  5 */ (n1570 ? (n1632 ? 1'b0 : !n1703) : (n1632 ? !n1703 : 1'b0));
assign n3294 = /* LUT   15 13  4 */ (n2251 ? n2121 : 1'b0);
assign n3295 = /* LUT    5 16  3 */ n766;
assign n3296 = /* LUT    4 20  6 */ (n785 ? (n623 ? 1'b1 : (n648 ? !n627 : 1'b1)) : 1'b0);
assign n3297 = /* LUT    4 12  2 */ (n740 ? (n579 ? 1'b0 : n274) : (n579 ? n274 : 1'b0));
assign n3298 = /* LUT   14 15  2 */ (n1795 ? (n1978 ? n1972 : 1'b0) : (n1978 ? 1'b0 : n1972));
assign n3299 = /* LUT    8 16  1 */ (n1198 ? (n912 ? (n1042 ? n212 : 1'b0) : 1'b0) : 1'b0);
assign n3300 = /* LUT    2  4  5 */ (n372 ? (n32 ? (n367 ? 1'b0 : n31) : 1'b0) : !n367);
assign n3301 = /* LUT   22  4  6 */ !n2770;
assign n3302 = /* LUT   14 18  7 */ !n1997;
assign n3303 = /* LUT   11  2  2 */ (n5 ? (n1249 ? 1'b0 : !n956) : (n1249 ? (n1398 ? 1'b0 : !n956) : !n956));
assign n3306 = /* LUT   15 14  5 */ (n2129 ? (n1790 ? 1'b0 : (n2252 ? !n1624 : 1'b0)) : 1'b0);
assign n3307 = /* LUT   15  6  1 */ (n1740 ? (n1903 ? !n2054 : (n1889 ? !n2054 : 1'b0)) : (n1903 ? !n2054 : (n1889 ? 1'b0 : !n2054)));
assign n3308 = /* LUT    5  9  0 */ (n545 ? (n564 ? 1'b0 : !n712) : (n5 ? (n564 ? 1'b0 : !n712) : !n712));
assign n3309 = /* LUT   24 13  4 */ n3018;
assign n3310 = /* LUT   12  2  7 */ !n1126;
assign n3311 = /* LUT    5  8  4 */ (n712 ? 1'b0 : (n213 ? !n564 : (n5 ? !n564 : 1'b1)));
assign n3314 = /* LUT    4  4  3 */ (n41 ? (n6 ? n666 : 1'b1) : (n6 ? n678 : 1'b0));
assign n3315 = /* LUT   11  3  3 */ (n852 ? n1412 : 1'b0);
assign n3318 = /* LUT    1 18  0 */ (n301 ? 1'b0 : n132);
assign n3319 = /* LUT   20 22  4 */ (n2156 ? (n2848 ? (n2293 ? n2297 : 1'b0) : 1'b0) : 1'b0);
assign n3323 = /* LUT    5  1  1 */ n177;
assign n3326 = /* LUT   17  9  4 */ (n2364 ? (n2355 ? !n2202 : 1'b1) : (n2355 ? !n2347 : 1'b0));
assign n3327 = /* LUT    7 12  3 */ n731;
assign n3328 = /* LUT    8  8  1 */ n15;
assign n3329 = /* LUT    5  4  6 */ (n665 ? (n6 ? (n381 ? n41 : 1'b1) : !n41) : (n6 ? (n381 ? n41 : 1'b1) : 1'b1));
assign n3330 = /* LUT   16 11  2 */ n1754;
assign n3331 = /* LUT   16 14  7 */ (n212 ? n1037 : 1'b0);
assign n3332 = /* LUT   17 10  5 */ (n2364 ? (n2230 ? !n2355 : 1'b1) : (n2355 ? !n2373 : 1'b0));
assign n3333 = /* LUT    7 13  4 */ (n895 ? (n899 ? 1'b0 : (n908 ? !n900 : 1'b1)) : (n899 ? 1'b0 : !n900));
assign n3334 = /* LUT   17  2  1 */ (n2182 ? (n2305 ? 1'b0 : n2311) : n2311);
assign n3335 = /* LUT    7  5  0 */ (n5 ? (n362 ? 1'b1 : n845) : (n362 ? n665 : n845));
assign n3336 = /* LUT    5  5  7 */ n15;
assign n3339 = /* LUT    4  1  6 */ (n6 ? (n657 ? (n659 ? 1'b0 : n41) : (n659 ? !n41 : 1'b1)) : 1'b1);
assign n3340 = /* LUT   14  3  4 */ (n1870 ? (n1727 ? (n1672 ? !n1875 : 1'b0) : n1672) : 1'b0);
assign n3341 = /* LUT    8  4  3 */ (n958 ? (n973 ? n861 : 1'b0) : 1'b0);
assign n3342 = /* LUT   16  7  4 */ (n2346 ? (n1893 ? 1'b0 : !n1883) : (n1893 ? !n1883 : 1'b0));
assign n3343 = /* LUT   13 19  5 */ (n2004 ? !n1648 : n1648);
assign n3344 = /* LUT   20 18  5 */ (n2156 ? (n2428 ? (n2293 ? 1'b0 : !n2297) : 1'b0) : 1'b0);
assign n3348 = /* LUT    1 14  7 */ (n45 ? n78 : !n78);
assign n3351 = /* LUT   10 12  4 */ (n1161 ? n1335 : (n1335 ? !n1303 : 1'b0));
assign n3352 = /* LUT    9  8  3 */ (n878 ? !n1267 : (n811 ? !n1267 : (n1267 ? 1'b0 : !n5)));
assign n3353 = /* LUT   13 20  6 */ (n2017 ? (n1647 ? n8 : !n8) : (n1647 ? !n8 : n8));
assign n3354 = /* LUT    2 18  1 */ (n300 ? 1'b1 : (n112 ? (n311 ? 1'b1 : n318) : 1'b1));
assign n3355 = /* LUT   21 22  5 */ (n2428 ? (n2297 ? (n2293 ? !n2156 : 1'b0) : 1'b0) : 1'b0);
assign n3356 = /* LUT   11 17  0 */ n233;
assign n3357 = /* LUT   18 16  0 */ n2413;
assign n3358 = /* LUT    3 18  6 */ (n461 ? (n309 ? n268 : 1'b0) : 1'b0);
assign n3359 = /* LUT   10  5  1 */ (n212 ? (n1424 ? !n861 : 1'b1) : !n975);
assign n3360 = /* LUT    9  1  0 */ (n1090 ? 1'b0 : !n1242);
assign n3361 = /* LUT    2 19  2 */ (n476 ? (n307 ? !n320 : 1'b0) : (n307 ? n320 : 1'b0));
assign n3362 = /* LUT    7  1  7 */ (n51 ? n52 : 1'b0);
assign n3363 = /* LUT    3 15  0 */ (n438 ? n287 : (n287 ? n597 : 1'b0));
assign n3364 = /* LUT   11 18  1 */ n1477;
assign n3365 = /* LUT   11 21  6 */ (n261 ? 1'b0 : (n1519 ? n1391 : 1'b0));
assign n3366 = /* LUT   12 17  4 */ (n1171 ? (n1505 ? 1'b1 : n1033) : n1505);
assign n3367 = /* LUT   12  9  0 */ (n1752 ? (n1270 ? 1'b0 : !n1577) : (n1270 ? 1'b0 : n1577));
assign n3368 = /* LUT    3 10  7 */ n233;
assign n3369 = /* LUT   22 12  0 */ n2650;
assign n3370 = /* LUT    3  2  3 */ n177;
assign n3371 = /* LUT   18 11  6 */ n2637;
assign n3372 = /* LUT   15 16  5 */ !n1624;
assign n3375 = /* LUT   11 13  7 */ n15;
assign n3376 = /* LUT   18 12  7 */ (n2521 ? (n2509 ? !n2500 : (n2381 ? 1'b1 : !n2500)) : (n2509 ? !n2500 : (n2381 ? n2500 : 1'b0)));
assign n3377 = /* LUT   11  5  3 */ n175;
assign n3378 = /* LUT   18  4  3 */ n2311;
assign n3381 = /* LUT    5 19  3 */ (n627 ? n765 : (n797 ? n765 : 1'b0));
assign n3382 = /* LUT    4 15  2 */ (n80 ? (n5 ? 1'b0 : (n134 ? !n132 : 1'b1)) : 1'b0);
assign n3383 = /* LUT   12  4  6 */ (n212 ? (n1538 ? n1397 : 1'b1) : !n1544);
assign n3386 = /* LUT    2  7  5 */ n233;
assign n3387 = /* LUT   22  7  6 */ (n2792 ? (n2692 ? (n2685 ? n2940 : 1'b0) : (n2685 ? !n2940 : 1'b1)) : (n2692 ? (n2685 ? 1'b1 : !n2940) : (n2685 ? 1'b0 : n2940)));
assign n3388 = /* LUT    3  3  3 */ (n362 ? (n5 ? 1'b1 : n355) : (n516 ? 1'b0 : !n5));
assign n3389 = /* LUT   21  3  5 */ (n2906 ? (n8 ? n2765 : !n2765) : (n8 ? !n2765 : n2765));
assign n3390 = /* LUT   14 21  7 */ (n2025 ? (n1665 ? 1'b0 : n1491) : n1491);
assign n3391 = /* LUT   11  6  4 */ (n212 ? 1'b0 : (n1563 ? !n852 : 1'b0));
assign n3393 = /* LUT   15  9  1 */ (n1882 ? !n1465 : (n1756 ? (n1465 ? 1'b0 : n1714) : (n1465 ? 1'b0 : !n1714)));
assign n3394 = /* LUT    5 12  0 */ (n698 ? (n450 ? !n564 : 1'b0) : !n564);
assign n3395 = /* LUT   17 21  5 */ (n2426 ? 1'b0 : (n2427 ? (n2292 ? 1'b0 : !n2022) : 1'b0));
assign n3396 = /* LUT   12  5  7 */ (n852 ? (n1564 ? (n816 ? n1001 : 1'b0) : 1'b0) : 1'b0);
assign n3397 = /* LUT   14 14  4 */ (n2126 ? (n1962 ? (n1494 ? n2124 : !n2124) : (n1494 ? n2124 : 1'b0)) : (n1962 ? (n1494 ? n2124 : 1'b1) : (n1494 ? n2124 : 1'b0)));
assign n3398 = /* LUT   14  6  0 */ (n1893 ? (n1434 ? 1'b0 : !n1883) : (n1434 ? !n1883 : 1'b0));
assign n3402 = /* LUT   23 12  1 */ (n2500 ? !n2809 : n2809);
assign n3403 = /* LUT    8 14  7 */ (n1041 ? (n1039 ? n932 : 1'b1) : 1'b1);
assign n3404 = /* LUT   20 17  0 */ (n2726 ? (n2408 ? n2843 : 1'b1) : (n2408 ? n2843 : n2560));
assign n3407 = /* LUT    5  7  6 */ (n552 ? (n6 ? 1'b1 : n212) : (n6 ? (n212 ? 1'b0 : n540) : n212));
assign n3408 = /* LUT    9 19  3 */ (n1019 ? 1'b0 : (n1061 ? 1'b0 : (n1044 ? 1'b0 : !n1043)));
assign n3409 = /* LUT    4  3  5 */ n189;
assign n3412 = /* LUT   16  9  3 */ (n2355 ? n2359 : (n2359 ? !n2356 : !n1597));
assign n3413 = /* LUT   20 21  6 */ (n2156 ? 1'b0 : (n2428 ? (n2293 ? !n2297 : 1'b0) : 1'b0));
assign n3414 = /* LUT   17 13  5 */ (n2540 ? !n2256 : n2256);
assign n3415 = /* LUT   17  5  1 */ n2329;
assign n3416 = /* LUT   20 13  2 */ (n2500 ? !n2703 : (n2529 ? (n2703 ? n2817 : 1'b1) : !n2703));
assign n3420 = /* LUT    5  8  7 */ (n5 ? (n712 ? 1'b0 : !n564) : (n712 ? 1'b0 : (n564 ? !n692 : 1'b1)));
assign n3421 = /* LUT   18 18  0 */ n2012;
assign n3422 = /* LUT    4  4  6 */ n189;
assign n3423 = /* LUT    7 11  5 */ (n711 ? 1'b1 : (n564 ? n889 : 1'b0));
assign n3424 = /* LUT   13 23  1 */ (n2030 ? (n2031 ? n1842 : !n1842) : n2031);
assign n3425 = /* LUT   16 10  4 */ (n2355 ? (n2226 ? !n2364 : 1'b0) : (n2374 ? !n2364 : 1'b0));
assign n3426 = /* LUT   13 22  5 */ (n1841 ? 1'b0 : !n5);
assign n3429 = /* LUT   14  2  7 */ (n1874 ? (n1263 ? 1'b0 : !n1822) : !n1263);
assign n3433 = /* LUT   10 16  0 */ n1362;
assign n3434 = /* LUT    1 17  7 */ (n307 ? !n126 : 1'b0);
assign n3435 = /* LUT   17  9  7 */ (n1928 ? (n2357 ? (n2355 ? n2215 : 1'b0) : n2215) : (n2357 ? (n2355 ? n2215 : !n2215) : (n2355 ? n2215 : 1'b1)));
assign n3436 = /* LUT    1  9  3 */ (n66 ? 1'b0 : n240);
assign n3437 = /* LUT    7  4  2 */ (n5 ? (n952 ? 1'b1 : n362) : (n952 ? (n381 ? 1'b1 : !n362) : (n381 ? n362 : 1'b0)));
assign n3438 = /* LUT    9 11  3 */ (n1170 ? (n1151 ? n1162 : 1'b0) : (n1151 ? (n1162 ? 1'b1 : n1160) : 1'b0));
assign n3439 = /* LUT   16  3  1 */ !n2315;
assign n3440 = /* LUT   13 15  2 */ (n1974 ? (n1788 ? n1806 : !n1806) : (n1788 ? !n1806 : n1806));
assign n3441 = /* LUT    7  3  6 */ (n942 ? 1'b0 : !n948);
assign n3442 = /* LUT   10 11  7 */ (n1171 ? 1'b0 : !n984);
assign n3443 = /* LUT   13 18  7 */ (n5 ? n1984 : (n1810 ? !n1650 : n1650));
assign n3444 = /* LUT    3 21  6 */ n277;
assign n3445 = /* LUT   10  8  1 */ (n1130 ? (n1442 ? (n708 ? !n1440 : 1'b1) : 1'b0) : (n1442 ? !n1440 : 1'b0));
assign n3446 = /* LUT   22 22  3 */ (n2296 ? (n2297 ? 1'b0 : (n2293 ? !n2156 : 1'b0)) : 1'b0);
assign n3447 = /* LUT    9  7  5 */ n175;
assign n3448 = /* LUT   13 11  4 */ n1718;
assign n3449 = /* LUT   21 21  7 */ (n2403 ? (n2878 ? 1'b0 : n2406) : (n3000 ? 1'b0 : n2406));
assign n3450 = /* LUT    3 14  3 */ n599;
assign n3451 = /* LUT   11 16  2 */ n1497;
assign n3457 = /* LUT    3 13  7 */ !n580;
assign n3458 = /* LUT   10 12  7 */ (n1312 ? 1'b0 : (n1296 ? 1'b0 : !n1350));
assign n3459 = /* LUT   10  4  3 */ (n956 ? 1'b0 : (n5 ? !n1410 : (n1410 ? !n1262 : 1'b1)));
assign n3460 = /* LUT    9  8  6 */ (n5 ? (n989 ? !n1267 : (n811 ? !n1267 : 1'b0)) : !n1267);
assign n3461 = /* LUT    2 18  4 */ (n306 ? !n142 : (n139 ? 1'b1 : (n151 ? !n142 : 1'b1)));
assign n3462 = /* LUT   21 14  4 */ (n2708 ? 1'b1 : n2706);
assign n3463 = /* LUT   11 17  3 */ n15;
assign n3464 = /* LUT    8 21  0 */ (n1069 ? (n1216 ? 1'b0 : !n924) : (n1216 ? 1'b0 : (n437 ? !n924 : 1'b0)));
assign n3465 = /* LUT   13  3  5 */ (n1420 ? n1106 : (n1543 ? (n816 ? n1106 : 1'b0) : 1'b0));
assign n3466 = /* LUT   18  7  3 */ n1757;
assign n3467 = /* LUT   15 20  6 */ (n1818 ? (n1827 ? !n5 : (n1646 ? 1'b0 : !n5)) : (n1827 ? (n1646 ? !n5 : 1'b0) : 1'b0));
assign n3468 = /* LUT   15 12  2 */ (n1891 ? (n2104 ? 1'b0 : !n2102) : !n2102);
assign n3469 = /* LUT    4 18  2 */ n778;
assign n3470 = /* LUT    2 10  5 */ (n243 ? (n423 ? 1'b0 : (n249 ? n199 : 1'b0)) : (n423 ? 1'b0 : n249));
assign n3471 = /* LUT    5 18  6 */ (n775 ? (n631 ? n189 : 1'b0) : (n787 ? 1'b1 : (n631 ? n189 : 1'b0)));
assign n3472 = /* LUT    2  2  1 */ (n163 ? (n167 ? !n200 : (n169 ? 1'b1 : !n200)) : (n169 ? 1'b1 : !n200));
assign n3473 = /* LUT   21  6  5 */ n2482;
assign n3474 = /* LUT   14 16  3 */ !n2128;
assign n3478 = /* LUT    5 15  0 */ (n756 ? 1'b0 : !n261);
assign n3479 = /* LUT    3  2  6 */ (n372 ? (n350 ? (n341 ? 1'b0 : n348) : 1'b0) : !n341);
assign n3480 = /* LUT   23 15  2 */ (n2975 ? (n3021 ? 1'b0 : (n2977 ? !n3023 : 1'b0)) : 1'b0);
assign n3481 = /* LUT   11  4  5 */ (n1414 ? (n1549 ? 1'b1 : n1410) : (n1549 ? (n5 ? 1'b1 : !n1410) : (n5 ? n1410 : 1'b0)));
assign n3482 = /* LUT   12  8  7 */ (n1575 ? (n1571 ? (n1598 ? 1'b1 : n1428) : 1'b0) : (n1571 ? (n1598 ? n1428 : 1'b1) : 1'b0));
assign n3483 = /* LUT    2  3  2 */ (n195 ? (n184 ? (n192 ? n187 : !n187) : 1'b0) : (n184 ? 1'b0 : (n192 ? n187 : !n187)));
assign n3484 = /* LUT   24 14  5 */ (n2818 ? 1'b0 : !n2827);
assign n3485 = /* LUT    4 14  4 */ !n582;
assign n3486 = /* LUT   14  9  0 */ (n1936 ? (n1702 ? 1'b0 : !n1595) : (n1702 ? !n1595 : 1'b0));
assign n3487 = /* LUT   11  5  6 */ (n1422 ? n816 : 1'b0);
assign n3490 = /* LUT   17  8  2 */ (n2072 ? (n2360 ? n2355 : (n1923 ? 1'b0 : !n2355)) : (n2360 ? 1'b1 : (n1923 ? 1'b0 : !n2355)));
assign n3494 = /* LUT    9 22  3 */ (n1393 ? !n931 : n931);
assign n3495 = /* LUT   17 11  7 */ (n2515 ? (n2366 ? 1'b1 : (n2514 ? 1'b1 : n2223)) : (n2366 ? 1'b0 : (n2514 ? 1'b1 : n2223)));
assign n3496 = /* LUT    4  6  5 */ (n547 ? (n51 ? 1'b0 : (n399 ? !n232 : 1'b1)) : (n51 ? 1'b0 : !n232));
assign n3497 = /* LUT    7 14  6 */ (n304 ? (n905 ? !n903 : 1'b0) : !n903);
assign n3498 = /* LUT    8 10  4 */ (n698 ? 1'b0 : (n1023 ? !n362 : 1'b1));
assign n3499 = /* LUT    8  2  0 */ (n200 ? (n1085 ? 1'b0 : !n1092) : n1076);
assign n3500 = /* LUT    1 20  2 */ (n332 ? !n148 : n148);
assign n3501 = /* LUT   14  4  6 */ (n1878 ? (n1249 ? (n1873 ? !n1700 : 1'b0) : n1873) : 1'b0);
assign n3502 = /* LUT   10 19  1 */ (n932 ? (n1373 ? 1'b1 : !n1031) : (n1374 ? (n1373 ? 1'b1 : !n1031) : 1'b0));
assign n3503 = /* LUT    5  3  3 */ n177;
assign n3504 = /* LUT   23  3  5 */ (n3050 ? (n3010 ? n8 : !n8) : (n3010 ? !n8 : n8));
assign n3505 = /* LUT    9 15  0 */ (n1193 ? (n1196 ? (n1036 ? n1038 : 1'b0) : 1'b0) : 1'b0);
assign n3506 = /* LUT   17  4  4 */ n2449;
assign n3507 = /* LUT    8  3  1 */ (n1099 ? (n176 ? 1'b0 : n1100) : 1'b0);
assign n3508 = /* LUT   16 13  4 */ n1965;
assign n3509 = /* LUT    4  2  7 */ (n353 ? (n518 ? (n212 ? !n52 : 1'b0) : 1'b0) : n212);
assign n3510 = /* LUT   16  5  0 */ n188;
assign n3511 = /* LUT   14  5  7 */ n189;
assign n3512 = /* LUT   18 22  1 */ (n2404 ? (n2403 ? n2586 : n2302) : n2403);
assign n3513 = /* LUT    1 12  3 */ (io_4_31_0 ? (n253 ? !n93 : 1'b1) : (n5 ? (n253 ? !n93 : 1'b1) : (n253 ? 1'b0 : n93)));
assign n3516 = /* LUT    7  7  2 */ !n868;
assign n3517 = /* LUT   16  6  1 */ (n2184 ? 1'b0 : (n2186 ? 1'b0 : (n2189 ? 1'b0 : !n2187)));
assign n3518 = /* LUT   10 14  7 */ (n1487 ? !n984 : 1'b0);
assign n3519 = /* LUT    9 10  6 */ (n1144 ? (n1146 ? n984 : 1'b0) : n984);
assign n3520 = /* LUT   16  9  6 */ (n2364 ? (n2080 ? (n2355 ? n1748 : 1'b1) : (n2355 ? n1748 : 1'b0)) : 1'b0);
assign n3521 = /* LUT    1  5  0 */ (n37 ? !n35 : n35);
assign n3522 = /* LUT    3 16  2 */ (n609 ? (io_4_31_0 ? 1'b0 : n45) : (n303 ? (io_4_31_0 ? 1'b0 : n45) : (io_4_31_0 ? !n45 : n45)));
assign n3526 = /* LUT   12 15  1 */ (n1634 ? !n1181 : (n1181 ? 1'b0 : n1476));
assign n3527 = /* LUT   20  4  5 */ (n7 ? (n2673 ? 1'b0 : (n2675 ? 1'b0 : !n2674)) : 1'b0);
assign n3528 = /* LUT   13 14  4 */ (n1785 ? (n1772 ? 1'b1 : n1960) : (n1772 ? 1'b0 : n1474));
assign n3529 = /* LUT   22 13  2 */ (n2720 ? (n2808 ? 1'b1 : (n2530 ? n2814 : 1'b0)) : (n2530 ? n2814 : 1'b0));
assign n3530 = /* LUT    3 17  3 */ (n313 ? (n300 ? !n295 : (n457 ? 1'b0 : !n295)) : 1'b0);
assign n3531 = /* LUT    1  9  6 */ (n72 ? 1'b0 : !n65);
assign n3532 = /* LUT   15 23  1 */ n2012;
assign n3533 = /* LUT   20  5  6 */ !n2683;
assign n3534 = /* LUT    9 11  6 */ (n5 ? 1'b1 : (n423 ? 1'b1 : (n258 ? !n249 : 1'b1)));
assign n3535 = /* LUT   12 19  7 */ (n1826 ? (n1820 ? !n5 : (n5 ? 1'b0 : n1646)) : (n1820 ? (n5 ? 1'b0 : !n1646) : 1'b0));
assign n3536 = /* LUT   18 10  4 */ n2067;
assign n3537 = /* LUT    9  3  2 */ n233;
assign n3538 = /* LUT   12 11  3 */ (n1608 ? (n1609 ? 1'b0 : (n1637 ? n5 : 1'b0)) : 1'b0);
assign n3539 = /* LUT   18  2  0 */ n2327;
assign n3540 = /* LUT   13  7  1 */ (n1910 ? (n1738 ? (n1579 ? n841 : 1'b0) : (n1579 ? 1'b1 : !n841)) : (n1579 ? 1'b1 : !n841));
assign n3541 = /* LUT   21 17  4 */ (n2984 ? (n2403 ? 1'b0 : (n2404 ? !n2853 : 1'b0)) : (n2403 ? 1'b0 : (n2404 ? !n2853 : 1'b1)));
assign n3542 = /* LUT   11 20  3 */ (n5 ? 1'b0 : (n188 ? (n1520 ? !n80 : 1'b1) : 1'b0));
assign n3543 = /* LUT    2 13  6 */ (n276 ? (n97 ? n435 : 1'b0) : 1'b0);
assign n3544 = /* LUT   13  6  5 */ (n1871 ? 1'b0 : (n1694 ? !n1891 : n1891));
assign n3545 = /* LUT    3  1  0 */ (n343 ? (n342 ? n6 : (n41 ? 1'b1 : n6)) : (n342 ? (n41 ? n6 : 1'b1) : 1'b1));
assign n3546 = /* LUT   22 14  2 */ (n3026 ? (n2966 ? n8 : !n8) : (n2966 ? !n8 : n8));
assign n3549 = /* LUT    3  4  5 */ (n6 ? (n41 ? 1'b1 : n192) : (n195 ? 1'b1 : !n41));
assign n3554 = /* LUT    5 13  2 */ (n754 ? n45 : 1'b0);
assign n3555 = /* LUT    4 17  5 */ (n111 ? (n612 ? 1'b1 : (n448 ? !n316 : 1'b1)) : 1'b1);
assign n3556 = /* LUT    4  9  1 */ (n398 ? !n711 : (n559 ? 1'b0 : !n711));
assign n3557 = /* LUT    3  5  6 */ (n6 ? (n390 ? (n41 ? !n365 : 1'b0) : (n41 ? !n365 : 1'b1)) : 1'b1);
assign n3558 = /* LUT   16 23  3 */ n2012;
assign n3561 = /* LUT   11  7  5 */ (n1122 ? n1419 : 1'b0);
assign n3562 = /* LUT   15 11  4 */ (n1330 ? 1'b0 : (n1473 ? 1'b0 : !n1329));
assign n3563 = /* LUT    2  6  2 */ (n392 ? (n176 ? 1'b0 : n222) : (n176 ? n222 : 1'b0));
assign n3564 = /* LUT    5 14  3 */ (n752 ? n128 : 1'b0);
assign n3565 = /* LUT   14 20  4 */ n1831;
assign n3566 = /* LUT    8 21  3 */ (n1064 ? (n771 ? 1'b1 : n925) : 1'b1);
assign n3567 = /* LUT   14 12  0 */ (n1770 ? 1'b0 : (n1593 ? 1'b1 : !n2102));
assign n3568 = /* LUT   21  5  7 */ (n2780 ? 1'b0 : (n2776 ? 1'b0 : (n2777 ? 1'b0 : !n2782)));
assign n3569 = /* LUT   17 20  2 */ (n2421 ? (n2411 ? (n2022 ? 1'b1 : !n2156) : (n2022 ? 1'b0 : !n2156)) : (n2411 ? (n2022 ? 1'b1 : n2156) : (n2022 ? 1'b0 : n2156)));
assign n3570 = /* LUT   11  8  6 */ (n1267 ? (n1428 ? 1'b0 : (n5 ? n1146 : 1'b0)) : n1146);
assign n3571 = /* LUT   15 12  5 */ (n2096 ? (n2238 ? 1'b1 : !n1452) : (n2238 ? 1'b0 : !n1452));
assign n3572 = /* LUT   15  4  1 */ n177;
assign n3573 = /* LUT   23 14  4 */ (n2972 ? (n3022 ? (n3020 ? 1'b1 : !n3025) : n3020) : (n3022 ? n3020 : (n3020 ? 1'b1 : !n3025)));
assign n3574 = /* LUT    4 10  1 */ n175;
assign n3575 = /* LUT   14 13  1 */ (n2107 ? 1'b0 : (n1772 ? (n1732 ? !n1494 : 1'b0) : !n1494));
assign n3576 = /* LUT   22  2  5 */ (n2888 ? !n2886 : (n2886 ? (n3007 ? n2891 : !n2891) : 1'b1));
assign n3577 = /* LUT    2  2  4 */ n177;
assign n3578 = /* LUT   16 24  3 */ (n2297 ? 1'b0 : (n2156 ? (n2298 ? n2293 : 1'b0) : 1'b0));
assign n3579 = /* LUT    7 17  6 */ !n477;
assign n3580 = /* LUT   14 16  6 */ (n1621 ? (n1980 ? !n1968 : n1968) : 1'b1);
assign n3583 = /* LUT    8 13  4 */ (n897 ? (n896 ? n1013 : (n1013 ? !n1030 : 1'b0)) : (n896 ? n1013 : 1'b0));
assign n3584 = /* LUT    8  5  0 */ n175;
assign n3585 = /* LUT   23  7  1 */ !n2621;
assign n3593 = /* LUT    7 10  3 */ n726;
assign n3594 = /* LUT    9 21  5 */ (n1031 ? !n175 : 1'b0);
assign n3595 = /* LUT    8  6  1 */ (n1106 ? (n816 ? n956 : 1'b0) : 1'b0);
assign n3596 = /* LUT   16  8  0 */ (n2053 ? !n2200 : (n1914 ? (n2200 ? 1'b0 : n2357) : (n2200 ? 1'b0 : !n2357)));
assign n3597 = /* LUT   20 20  3 */ (n2406 ? (n2863 ? 1'b1 : n2408) : (n2583 ? 1'b1 : n2408));
assign n3598 = /* LUT   14  8  7 */ (n1556 ? (n1700 ? 1'b0 : !n1931) : (n1700 ? !n1931 : 1'b0));
assign n3599 = /* LUT    8  9  6 */ n233;
assign n3600 = /* LUT   17  8  5 */ n2067;
assign n3603 = /* LUT    9 22  6 */ (n1069 ? (n924 ? n1231 : 1'b0) : (n437 ? (n924 ? n1231 : 1'b0) : n1231));
assign n3604 = /* LUT    5  2  5 */ (n493 ? 1'b0 : (n52 ? 1'b0 : (n805 ? 1'b0 : n51)));
assign n3605 = /* LUT   23  2  7 */ (n3046 ? (n8 ? n2892 : !n2892) : (n8 ? !n2892 : n2892));
assign n3606 = /* LUT    9 14  2 */ n175;
assign n3607 = /* LUT   16 12  6 */ (n2245 ? (n1624 ? 1'b0 : n1790) : 1'b0);
assign n3608 = /* LUT   16  4  2 */ (io_19_0_1 ? (n2303 ? n2333 : 1'b0) : 1'b0);
assign n3614 = /* LUT    8  1  7 */ (n1081 ? 1'b0 : !n1083);
assign n3615 = /* LUT   12 18  1 */ n1609;
assign n3618 = /* LUT   10 10  4 */ (n334 ? (n1308 ? 1'b1 : (n1318 ? 1'b1 : n679)) : (n1308 ? !n679 : (n1318 ? !n679 : 1'b0)));
assign n3619 = /* LUT   10  2  0 */ (n1241 ? (n1249 ? 1'b0 : n1256) : (n1249 ? (n1256 ? !n5 : 1'b0) : n1256));
assign n3620 = /* LUT    9  6  3 */ (n1121 ? (n697 ? (n1117 ? 1'b0 : !n1269) : !n1269) : (n1117 ? 1'b0 : !n1269));
assign n3621 = /* LUT   22 16  2 */ (n2406 ? (n3033 ? !n2404 : 1'b0) : (n3034 ? !n2404 : 1'b0));
assign n3622 = /* LUT   13  9  0 */ (n1585 ? (n1594 ? !n212 : (n1711 ? 1'b1 : !n212)) : 1'b0);
assign n3623 = /* LUT    2 16  1 */ (n120 ? n119 : 1'b0);
assign n3624 = /* LUT    3 20  3 */ (n644 ? (n628 ? 1'b0 : (n627 ? 1'b0 : !n469)) : (n628 ? !n627 : (n627 ? 1'b0 : !n469)));
assign n3625 = /* LUT   21 20  5 */ (n2156 ? 1'b0 : (n2855 ? (n2293 ? !n2297 : 1'b0) : 1'b0));
assign n3626 = /* LUT   21 12  1 */ (n2809 ? (n2390 ? !n2509 : 1'b0) : (n2390 ? (n2525 ? n2509 : 1'b0) : 1'b0));
assign n3627 = /* LUT    1 12  6 */ (n113 ? (n102 ? n271 : 1'b0) : 1'b0);
assign n3628 = /* LUT    1  4  2 */ n27;
assign n3629 = /* LUT   20  8  6 */ n2197;
assign n3630 = /* LUT   12 22  7 */ (n1835 ? (n5 ? 1'b0 : n1664) : (n5 ? 1'b0 : n1849));
assign n3631 = /* LUT   18 13  4 */ n2648;
assign n3632 = /* LUT   12 14  3 */ (n1794 ? (n1619 ? 1'b0 : n1623) : (n1619 ? n1623 : 1'b0));
assign n3633 = /* LUT   18  5  0 */ (n2452 ? (n2451 ? (n2453 ? n2450 : 1'b0) : 1'b0) : 1'b0);
assign n3634 = /* LUT   22 17  3 */ (n2293 ? 1'b0 : (n2986 ? (n2156 ? !n2297 : 1'b0) : 1'b0));
assign n3635 = /* LUT    2 17  2 */ (n458 ? !n315 : n315);
assign n3636 = /* LUT   13 10  1 */ n1556;
assign n3637 = /* LUT    9  2  5 */ (n41 ? (n6 ? !n1078 : 1'b1) : (n6 ? !n1082 : 1'b1));
assign n3641 = /* LUT   21 16  7 */ n2012;
assign n3642 = /* LUT   20  1  3 */ (n2760 ? !n2448 : n2448);
assign n3643 = /* LUT   10  3  0 */ n15;
assign n3644 = /* LUT   18  6  1 */ (n2481 ? !n2465 : n2465);
assign n3645 = /* LUT   12  7  0 */ (n1581 ? (n1713 ? 1'b0 : (n1562 ? !n1710 : 1'b0)) : 1'b0);
assign n3648 = /* LUT   18  9  6 */ (n2495 ? (n2355 ? 1'b1 : !n2069) : (n2355 ? 1'b0 : !n1596));
assign n3649 = /* LUT   12  6  4 */ (n1555 ? !n1717 : (n1698 ? (n1556 ? !n1717 : 1'b0) : (n1556 ? 1'b0 : !n1717)));
assign n3650 = /* LUT    5 16  2 */ (n611 ? (n767 ? 1'b0 : (n249 ? 1'b0 : !n449)) : (n767 ? 1'b0 : !n249));
assign n3651 = /* LUT   11 19  5 */ (n426 ? (n5 ? n1519 : (n1519 ? n1477 : 1'b0)) : n1519);
assign n3652 = /* LUT    4 20  5 */ (n175 ? n631 : 1'b0);
assign n3655 = /* LUT   13  5  7 */ n15;
assign n3656 = /* LUT   14 15  1 */ (n1541 ? 1'b1 : n1966);
assign n3659 = /* LUT    2  4  4 */ (n33 ? !n37 : n37);
assign n3660 = /* LUT    3  8  6 */ (n416 ? (n230 ? (n417 ? n227 : 1'b0) : (n417 ? 1'b0 : n227)) : (n230 ? (n417 ? !n227 : 1'b0) : (n417 ? 1'b0 : !n227)));
assign n3661 = /* LUT   17 22  1 */ n2012;
assign n3662 = /* LUT   18  2  3 */ n2321;
assign n3663 = /* LUT    5 17  3 */ (n772 ? 1'b0 : (n773 ? n268 : 1'b0));
assign n3664 = /* LUT   15  6  0 */ (n1416 ? (n1726 ? (n2194 ? n2066 : 1'b0) : (n2194 ? 1'b1 : !n2066)) : (n1726 ? (n2194 ? 1'b1 : !n2066) : (n2194 ? n2066 : 1'b0)));
assign n3667 = /* LUT   12  2  6 */ !n1125;
assign n3668 = /* LUT    2  5  5 */ (n191 ? (n41 ? 1'b1 : (n35 ? 1'b1 : !n6)) : (n41 ? n6 : (n35 ? 1'b1 : !n6)));
assign n3669 = /* LUT   16 19  0 */ n2419;
assign n3670 = /* LUT    4 16  7 */ (n605 ? (n448 ? 1'b1 : (n249 ? n117 : 1'b0)) : (n249 ? n117 : 1'b0));
assign n3671 = /* LUT    3  1  3 */ (n338 ? (n232 ? !n340 : 1'b0) : n232);
assign n3672 = /* LUT   11 11  6 */ (n1564 ? n816 : 1'b0);
assign n3673 = /* LUT   11  3  2 */ (n1417 ? (n1410 ? (n5 ? 1'b1 : n1409) : 1'b1) : (n1410 ? (n5 ? 1'b1 : n1409) : 1'b0));
assign n3674 = /* LUT   15 15  5 */ (n1037 ? (n212 ? 1'b1 : n1790) : (n212 ? !n1790 : n1790));
assign n3675 = /* LUT   14 11  3 */ n1892;
assign n3676 = /* LUT   14 19  7 */ (n2007 ? !n1966 : n1966);
assign n3677 = /* LUT   15  7  1 */ (n1749 ? (n1702 ? 1'b0 : !n1595) : (n1702 ? !n1595 : 1'b0));
assign n3678 = /* LUT    5 10  0 */ (n726 ? (n711 ? n5 : 1'b1) : 1'b0);
assign n3679 = /* LUT    7 21  2 */ (n1071 ? 1'b0 : (n437 ? 1'b1 : n1069));
assign n3680 = /* LUT   12  3  7 */ (n1680 ? 1'b0 : (n807 ? !n1539 : 1'b1));
assign n3681 = /* LUT   22  5  5 */ n2170;
assign n3682 = /* LUT    5 13  5 */ (n630 ? !n362 : (n362 ? 1'b0 : !n679));
assign n3683 = /* LUT    4  9  4 */ (n559 ? (n401 ? !n711 : 1'b0) : !n711);
assign n3684 = /* LUT    8  8  0 */ !n867;
assign n3688 = /* LUT   17 10  4 */ (n2490 ? (n2355 ? n2504 : (n2365 ? 1'b0 : n2504)) : (n2355 ? n2504 : (n2365 ? !n2504 : 1'b1)));
assign n3689 = /* LUT    7 13  3 */ (n759 ? !n564 : (n698 ? 1'b0 : !n564));
assign n3690 = /* LUT   15  2  7 */ (n1863 ? (n1408 ? 1'b0 : !n2169) : !n1408);
assign n3691 = /* LUT    5  5  6 */ n189;
assign n3694 = /* LUT    4  1  5 */ (n371 ? 1'b0 : !n51);
assign n3695 = /* LUT   14  3  3 */ n354;
assign n3696 = /* LUT    8  4  2 */ (n971 ? (n1101 ? 1'b0 : n964) : !n1101);
assign n3697 = /* LUT   16 15  7 */ n2132;
assign n3698 = /* LUT   20 18  4 */ (n2403 ? (n2728 ? !n2404 : 1'b0) : (n2725 ? !n2404 : 1'b0));
assign n3699 = /* LUT   17  3  1 */ (n2319 ? 1'b1 : n2323);
assign n3700 = /* LUT    7  6  0 */ (n861 ? (n967 ? (n976 ? 1'b1 : n977) : n977) : n977);
assign n3701 = /* LUT    9 17  2 */ n1201;
assign n3702 = /* LUT    7  9  5 */ n1005;
assign n3703 = /* LUT    8  5  3 */ (n976 ? (n958 ? (n1115 ? 1'b1 : n1116) : n1116) : (n958 ? n1115 : 1'b0));
assign n3704 = /* LUT   13 20  5 */ (n2016 ? (n8 ? n1648 : !n1648) : (n8 ? !n1648 : n1648));
assign n3705 = /* LUT   20 11  1 */ n2632;
assign n3706 = /* LUT   10 14  0 */ (n212 ? (n819 ? 1'b1 : n1459) : 1'b0);
assign n3707 = /* LUT   18 24  3 */ n2012;
assign n3708 = /* LUT   17  7  7 */ (n2341 ? 1'b0 : (n2375 ? n2345 : 1'b0));
assign n3709 = /* LUT    3 18  5 */ (n463 ? (n312 ? 1'b0 : !n464) : !n464);
assign n3710 = /* LUT   16  8  3 */ (n2169 ? 1'b0 : (n2179 ? !n2356 : n2356));
assign n3711 = /* LUT    2 19  1 */ (n323 ? (n319 ? 1'b0 : n307) : (n319 ? n307 : 1'b0));
assign n3712 = /* LUT    7  1  6 */ (n679 ? (n658 ? 1'b1 : n5) : (n834 ? 1'b0 : !n5));
assign n3713 = /* LUT   13 13  2 */ (n1624 ? 1'b0 : (n1957 ? n1790 : 1'b0));
assign n3714 = /* LUT   18 17  0 */ n2012;
assign n3715 = /* LUT    1  7  2 */ (n229 ? (n48 ? n64 : !n64) : (n48 ? !n64 : n64));
assign n3716 = /* LUT   13 16  7 */ (n1982 ? (n212 ? 1'b1 : n1125) : (n212 ? n1125 : 1'b0));
assign n3717 = /* LUT    3 19  6 */ (n321 ? 1'b0 : n462);
assign n3718 = /* LUT   20  3  2 */ n2601;
assign n3719 = /* LUT   11 21  5 */ (n1521 ? (n5 ? 1'b0 : (n1525 ? 1'b0 : !n1511)) : (n5 ? 1'b0 : !n1525));
assign n3720 = /* LUT   12 17  3 */ (n1033 ? (n1507 ? 1'b1 : n1495) : n1507);
assign n3721 = /* LUT   20  6  7 */ (n2693 ? 1'b1 : n1);
assign n3722 = /* LUT    2 20  2 */ (n142 ? (n475 ? (n45 ? 1'b0 : !n318) : !n318) : !n318);
assign n3723 = /* LUT   10  9  6 */ (n1267 ? 1'b0 : (n1000 ? 1'b1 : (n811 ? 1'b1 : !n5)));
assign n3724 = /* LUT    9  5  5 */ (n5 ? 1'b0 : n841);
assign n3725 = /* LUT    1  8  3 */ n236;
assign n3726 = /* LUT   21 19  7 */ (n2293 ? (n2297 ? 1'b0 : (n2855 ? n2156 : 1'b0)) : 1'b0);
assign n3727 = /* LUT    3 11  1 */ !n579;
assign n3728 = /* LUT   11 14  2 */ (n1478 ? (n212 ? !n1146 : 1'b0) : 1'b0);
assign n3729 = /* LUT   12 18  4 */ n1644;
assign n3730 = /* LUT   12 10  0 */ n177;
assign n3731 = /* LUT   10 10  7 */ n1459;
assign n3732 = /* LUT   10  2  3 */ (n1249 ? (n1396 ? 1'b0 : (n5 ? 1'b0 : !n956)) : !n956);
assign n3733 = /* LUT   18 12  6 */ n2636;
assign n3734 = /* LUT    9  6  6 */ n1123;
assign n3735 = /* LUT   18  4  2 */ n2310;
assign n3736 = /* LUT   22 16  5 */ (n2156 ? (n2293 ? 1'b0 : (n2992 ? !n2297 : 1'b0)) : 1'b0);
assign n3737 = /* LUT   22  8  1 */ (n3014 ? 1'b0 : (n1 ? 1'b0 : (n1645 ? 1'b0 : !n2946)));
assign n3738 = /* LUT   21 12  4 */ (n2698 ? n2704 : 1'b0);
assign n3739 = /* LUT   21  4  0 */ (n2909 ? (n8 ? !n2672 : n2672) : (n8 ? n2672 : !n2672));
assign n3743 = /* LUT    3  3  2 */ n179;
assign n3744 = /* LUT   18 13  7 */ n2652;
assign n3745 = /* LUT   18  5  3 */ n2318;
assign n3746 = /* LUT    5 20  3 */ (n645 ? (n627 ? n785 : (n628 ? n785 : 1'b0)) : (n627 ? n785 : 1'b0));
assign n3747 = /* LUT   17 21  4 */ (n2428 ? (n2293 ? (n2156 ? n2297 : 1'b0) : 1'b0) : 1'b0);
assign n3748 = /* LUT   12  5  6 */ (n1694 ? 1'b0 : n956);
assign n3749 = /* LUT    8 20  1 */ (n1220 ? (n797 ? !n1211 : 1'b0) : 1'b0);
assign n3752 = /* LUT    2  8  5 */ !n66;
assign n3753 = /* LUT    4 19  7 */ (n784 ? (n472 ? (n785 ? !n786 : 1'b1) : 1'b1) : !n785);
assign n3754 = /* LUT   14 14  3 */ (n2128 ? 1'b0 : (n1766 ? n2129 : 1'b0));
assign n3755 = /* LUT   15 10  1 */ (n1888 ? (n1756 ? n2077 : (n2077 ? n2049 : 1'b0)) : (n1756 ? (n2077 ? n2049 : 1'b0) : n2077));
assign n3756 = /* LUT   12  6  7 */ (n1564 ? (n816 ? n956 : 1'b0) : 1'b0);
assign n3757 = /* LUT   15 13  6 */ (n2109 ? (n1494 ? n2127 : n1943) : (n1494 ? n2127 : (n1943 ? !n2127 : 1'b0)));
assign n3758 = /* LUT    5 16  5 */ (n455 ? 1'b1 : (n266 ? 1'b1 : !n758));
assign n3759 = /* LUT    4 12  4 */ (n742 ? (n581 ? 1'b0 : n274) : (n581 ? n274 : 1'b0));
assign n3760 = /* LUT   14 15  4 */ (n1517 ? (n1 ? 1'b1 : n1645) : n1);
assign n3761 = /* LUT    2  4  7 */ (n6 ? (n41 ? n33 : 1'b1) : (n193 ? 1'b1 : n41));
assign n3762 = /* LUT   23 13  1 */ (n3052 ? n2841 : 1'b0);
assign n3766 = /* LUT   11  2  4 */ n188;
assign n3771 = /* LUT   15  6  3 */ (n2193 ? (n2066 ? n2197 : !n1126) : (n2066 ? n2197 : n1126));
assign n3772 = /* LUT    5  8  6 */ (n719 ? (n551 ? (n703 ? !n701 : 1'b0) : 1'b1) : 1'b0);
assign n3778 = /* LUT   16 10  3 */ (n2217 ? (n2219 ? n2366 : (n2366 ? n2225 : 1'b0)) : (n2219 ? 1'b1 : (n2366 ? n2225 : 1'b1)));
assign n3779 = /* LUT   17  6  1 */ n2473;
assign n3780 = /* LUT   14  2  6 */ (n1550 ? n1864 : 1'b0);
assign n3781 = /* LUT    9 20  2 */ (n1382 ? (n1061 ? (n8 ? n1064 : 1'b0) : (n8 ? 1'b0 : n1064)) : (n1061 ? (n8 ? 1'b0 : n1064) : (n8 ? n1064 : 1'b0)));
assign n3782 = /* LUT    5  1  3 */ (n501 ? (n5 ? n362 : (n359 ? n362 : 1'b0)) : (n5 ? n362 : (n359 ? 1'b1 : !n362)));
assign n3783 = /* LUT   17  9  6 */ n1754;
assign n3784 = /* LUT   18 19  0 */ n2012;
assign n3785 = /* LUT    7 12  5 */ n732;
assign n3786 = /* LUT    7  4  1 */ (n847 ? (n356 ? 1'b1 : (n362 ? n5 : 1'b1)) : (n356 ? n362 : (n362 ? n5 : 1'b0)));
assign n3787 = /* LUT    8  8  3 */ !n870;
assign n3788 = /* LUT   16 11  4 */ (n2376 ? !n2222 : (n2366 ? (n2235 ? !n2222 : 1'b0) : !n2222));
assign n3789 = /* LUT   16  3  0 */ n15;
assign n3792 = /* LUT   17 10  7 */ n2204;
assign n3793 = /* LUT   17  2  3 */ (n2182 ? (n2313 ? io_19_0_1 : 1'b0) : 1'b0);
assign n3794 = /* LUT    3 21  5 */ n5;
assign n3795 = /* LUT    7  5  2 */ (n698 ? (n5 ? 1'b1 : n678) : n842);
assign n3798 = /* LUT   12 20  4 */ (n1652 ? 1'b0 : (n1653 ? 1'b0 : (n15 ? !n5 : 1'b0)));
assign n3799 = /* LUT   14  3  6 */ n175;
assign n3800 = /* LUT   16  7  6 */ n2204;
assign n3801 = /* LUT   13 19  7 */ (n1828 ? (n1646 ? !n5 : (n5 ? 1'b0 : n1819)) : (n1646 ? 1'b0 : (n5 ? 1'b0 : n1819)));
assign n3804 = /* LUT    1  6  5 */ n216;
assign n3805 = /* LUT   10 12  6 */ (n1319 ? 1'b0 : (n1327 ? (n1462 ? !n1168 : 1'b1) : !n1462));
assign n3806 = /* LUT   10  4  2 */ (n5 ? (n956 ? 1'b0 : !n1249) : (n1236 ? (n956 ? 1'b0 : !n1249) : !n956));
assign n3807 = /* LUT    9  8  5 */ (n1276 ? (n1133 ? n707 : 1'b1) : 1'b0);
assign n3808 = /* LUT    2 18  3 */ (n318 ? 1'b0 : (n112 ? (n300 ? 1'b0 : n459) : 1'b0));
assign n3809 = /* LUT   13 12  4 */ (n1763 ? (n1494 ? 1'b1 : n1718) : (n1494 ? 1'b0 : n1718));
assign n3810 = /* LUT   13  4  0 */ (n1715 ? (n1543 ? (n1699 ? 1'b0 : !n1874) : !n1874) : (n1543 ? !n1699 : 1'b1));
assign n3811 = /* LUT   21 14  3 */ (n2958 ? 1'b1 : n2812);
assign n3812 = /* LUT   11 17  2 */ (n151 ? (n1512 ? 1'b0 : n1469) : (n1512 ? (n1469 ? !n277 : 1'b0) : 1'b0));
assign n3813 = /* LUT   12 13  0 */ (n1622 ? (n1617 ? (n1604 ? n1612 : 1'b0) : (n1604 ? 1'b0 : n1612)) : (n1617 ? (n1604 ? !n1612 : 1'b0) : (n1604 ? 1'b0 : !n1612)));
assign n3814 = /* LUT   20  2  4 */ (n2668 ? 1'b1 : n2669);
assign n3815 = /* LUT   18  7  2 */ n2204;
assign n3816 = /* LUT   22 19  5 */ (n2426 ? (n2427 ? (n2022 ? 1'b0 : n2292) : 1'b0) : 1'b0);
assign n3817 = /* LUT    2 19  4 */ (n45 ? 1'b0 : (n475 ? (n139 ? !n327 : 1'b0) : 1'b0));
assign n3818 = /* LUT    2 11  0 */ (n243 ? (n251 ? 1'b1 : n42) : 1'b0);
assign n3819 = /* LUT   21 15  4 */ (n2820 ? 1'b0 : (n2824 ? 1'b0 : !n2821));
assign n3820 = /* LUT   11 18  3 */ (n1509 ? 1'b0 : n1518);
assign n3824 = /* LUT    8 22  0 */ (n924 ? !n1228 : (n1069 ? 1'b0 : (n437 ? 1'b0 : !n1228)));
assign n3825 = /* LUT   18  8  3 */ (n2341 ? (n2345 ? !n2375 : 1'b0) : 1'b0);
assign n3826 = /* LUT   12  9  2 */ (n1590 ? 1'b0 : (n1735 ? 1'b0 : n1584));
assign n3827 = /* LUT    3  2  5 */ n354;
assign n3828 = /* LUT   12  8  6 */ n354;
assign n3829 = /* LUT   15 16  7 */ (n1624 ? (n1623 ? !n1790 : 1'b0) : (n1623 ? n1790 : 1'b0));
assign n3830 = /* LUT    2  3  1 */ n180;
assign n3831 = /* LUT    4 14  3 */ (n455 ? (n132 ? 1'b0 : (n436 ? !n594 : 1'b0)) : (n132 ? 1'b0 : !n594));
assign n3832 = /* LUT   14 17  3 */ (n1636 ? 1'b0 : !n1986);
assign n3833 = /* LUT    8 18  2 */ !n630;
assign n3837 = /* LUT   17 17  1 */ (n2011 ? n2412 : n2554);
assign n3838 = /* LUT   11  5  5 */ (n1539 ? (n1425 ? !n212 : 1'b0) : 1'b0);
assign n3841 = /* LUT    5 19  5 */ (n785 ? (n784 ? !n786 : 1'b0) : 1'b1);
assign n3842 = /* LUT    5 11  1 */ (n733 ? (n731 ? 1'b0 : n764) : (n731 ? n764 : 1'b0));
assign n3843 = /* LUT    4 15  4 */ (n593 ? (n756 ? 1'b0 : (n286 ? !n758 : 1'b1)) : !n756);
assign n3844 = /* LUT    4  7  0 */ n179;
assign n3845 = /* LUT    2  7  7 */ (n363 ? (n391 ? 1'b0 : !n114) : !n391);
assign n3846 = /* LUT   14 10  0 */ n1925;
assign n3847 = /* LUT    3  3  5 */ (n366 ? (n223 ? n363 : 1'b0) : (n223 ? (n514 ? n363 : 1'b1) : 1'b0));
assign n3848 = /* LUT   21  3  7 */ (n2908 ? (n2767 ? n8 : !n8) : (n2767 ? !n8 : n8));
assign n3849 = /* LUT   11  6  6 */ n188;
assign n3850 = /* LUT   15  9  3 */ n2067;
assign n3851 = /* LUT    5 12  2 */ (n103 ? (n212 ? !n483 : 1'b1) : (n212 ? (n261 ? !n483 : 1'b0) : (n261 ? 1'b1 : n483)));
assign n3852 = /* LUT    4  8  1 */ (n398 ? (n8 ? n401 : !n401) : (n8 ? !n401 : n401));
assign n3853 = /* LUT   14  6  2 */ (n1727 ? 1'b0 : (n1901 ? !n1934 : n1934));
assign n3854 = /* LUT    8  3  0 */ (n1086 ? (n1089 ? !n176 : 1'b0) : 1'b0);
assign n3855 = /* LUT    1 21  2 */ (n336 ? (n153 ? 1'b0 : n157) : (n153 ? n157 : 1'b0));
assign n3856 = /* LUT   15  1  4 */ (n1875 ? n1704 : 1'b0);
assign n3859 = /* LUT    7  7  1 */ (n863 ? (n859 ? n868 : 1'b0) : (n859 ? !n868 : 1'b0));
assign n3860 = /* LUT    9 19  5 */ (n1189 ? 1'b0 : (n1210 ? (n1209 ? !n1050 : 1'b0) : 1'b0));
assign n3861 = /* LUT    4  3  7 */ (n389 ? (n41 ? (n658 ? !n6 : 1'b1) : n6) : (n41 ? (n658 ? !n6 : 1'b1) : 1'b1));
assign n3862 = /* LUT   16  6  0 */ (n1884 ? 1'b0 : (n1891 ? !n1542 : n1542));
assign n3863 = /* LUT    8  7  6 */ (n1127 ? !n854 : 1'b0);
assign n3864 = /* LUT   16  9  5 */ (n2346 ? (n2364 ? 1'b1 : n1930) : (n2364 ? 1'b0 : n1930));
assign n3865 = /* LUT   17 13  7 */ !n2257;
assign n3866 = /* LUT   17  5  3 */ n2326;
assign n3867 = /* LUT   20 13  4 */ (n2720 ? (n2528 ? (n2814 ? 1'b1 : n2524) : n2524) : (n2528 ? n2814 : 1'b0));
assign n3868 = /* LUT    7  8  2 */ (n991 ? (n866 ? 1'b0 : n981) : (n866 ? n981 : 1'b0));
assign n3869 = /* LUT   18 18  2 */ (n2156 ? (n2293 ? (n2432 ? n2297 : 1'b0) : 1'b0) : 1'b0);
assign n3870 = /* LUT   16 10  6 */ (n2361 ? (n2368 ? 1'b1 : !n2366) : (n2368 ? (n2214 ? 1'b1 : n2366) : (n2214 ? !n2366 : 1'b0)));
assign n3871 = /* LUT   13 22  7 */ (n1844 ? n1842 : 1'b1);
assign n3872 = /* LUT   13 14  3 */ (n1494 ? 1'b0 : (n1772 ? n1598 : 1'b1));
assign n3873 = /* LUT    3 17  2 */ (n616 ? !n615 : n615);
assign n3874 = /* LUT   18 19  3 */ !n2397;
assign n3875 = /* LUT    1  9  5 */ n72;
assign n3876 = /* LUT   20  5  5 */ !n2675;
assign n3877 = /* LUT    9 11  5 */ (n898 ? (n1165 ? !n1156 : 1'b0) : (n1165 ? (n1159 ? 1'b1 : !n1156) : 1'b0));
assign n3878 = /* LUT   13 15  4 */ (n1976 ? (n1804 ? n1803 : !n1803) : (n1804 ? !n1803 : n1803));
assign n3879 = /* LUT   13  7  0 */ (n1749 ? (n1887 ? 1'b0 : !n1689) : (n1887 ? !n1689 : 1'b0));
assign n3880 = /* LUT    1  2  2 */ n22;
assign n3881 = /* LUT   10  8  3 */ n1146;
assign n3882 = /* LUT   12 20  7 */ (n5 ? 1'b0 : (n1652 ? 1'b0 : (n179 ? !n1653 : 1'b0)));
assign n3883 = /* LUT    9  4  2 */ (n1112 ? (n806 ? 1'b0 : (n1105 ? n1097 : 1'b1)) : (n806 ? 1'b0 : n1097));
assign n3884 = /* LUT   22 14  1 */ (n2976 ? (n3019 ? n8 : !n8) : (n3019 ? !n8 : n8));
assign n3885 = /* LUT    2 14  0 */ (n45 ? n80 : 1'b0);
assign n3886 = /* LUT   13  8  1 */ (n1037 ? (n1465 ? (n1736 ? 1'b1 : n1724) : n1736) : (n1465 ? 1'b1 : !n1724));
assign n3887 = /* LUT    9  7  7 */ (n477 ? (n852 ? n679 : (n1116 ? 1'b1 : n679)) : (n852 ? 1'b0 : (n1116 ? !n679 : 1'b0)));
assign n3888 = /* LUT   13 11  6 */ n1452;
assign n3889 = /* LUT   10  1  0 */ (n1236 ? (n1396 ? (n6 ? !n41 : n41) : (n6 ? 1'b1 : n41)) : (n1396 ? (n6 ? !n41 : 1'b1) : 1'b1));
assign n3890 = /* LUT   11 16  4 */ (n212 ? (n422 ? 1'b1 : n1459) : 1'b0);
assign n3891 = /* LUT   12 12  2 */ (n1768 ? (n1600 ? n1766 : !n1766) : (n1600 ? !n1766 : n1766));
assign n3894 = /* LUT    3  5  5 */ (n536 ? (n535 ? (n377 ? 1'b1 : n51) : 1'b1) : (n535 ? (n377 ? !n51 : 1'b0) : !n51));
assign n3895 = /* LUT   10  4  5 */ (n1413 ? (n1253 ? 1'b1 : !n1107) : (n1253 ? !n1259 : (n1259 ? 1'b0 : !n1107)));
assign n3896 = /* LUT   15 19  7 */ (n1998 ? 1'b0 : n1652);
assign n3897 = /* LUT   22 18  7 */ (n2990 ? (n2403 ? (n2404 ? n3038 : 1'b0) : n2404) : (n2403 ? (n2404 ? n3038 : 1'b0) : 1'b0));
assign n3900 = /* LUT    5 14  2 */ (n748 ? 1'b0 : (n249 ? (n266 ? 1'b1 : n578) : 1'b0));
assign n3901 = /* LUT   21 14  6 */ (n2961 ? n2824 : (n2824 ? n2830 : 1'b0));
assign n3902 = /* LUT   11  9  1 */ (n5 ? (n1548 ? !n1146 : 1'b0) : !n1146);
assign n3903 = /* LUT    8 21  2 */ (n1215 ? 1'b0 : (n437 ? !n924 : (n1069 ? !n924 : 1'b0)));
assign n3904 = /* LUT   13  3  7 */ (n1675 ? (n1554 ? 1'b1 : !n1875) : (n1554 ? n1875 : 1'b0));
assign n3905 = /* LUT    3  6  6 */ (n51 ? 1'b0 : !n52);
assign n3906 = /* LUT   17 20  1 */ (n2292 ? (n2022 ? n2409 : !n2427) : (n2022 ? n2409 : n2427));
assign n3907 = /* LUT   11  8  5 */ (n1146 ? (n1267 ? (n1270 ? 1'b0 : n5) : 1'b1) : 1'b0);
assign n3908 = /* LUT   18  7  5 */ n1789;
assign n3909 = /* LUT   15 12  4 */ (n2243 ? (n1945 ? !n1941 : 1'b0) : (n1778 ? n1945 : (n1945 ? !n1941 : 1'b0)));
assign n3910 = /* LUT   15  4  0 */ (n1249 ? n1179 : 1'b0);
assign n3911 = /* LUT    4 18  4 */ n779;
assign n3912 = /* LUT    4 10  0 */ n188;
assign n3913 = /* LUT    8 22  3 */ (n1069 ? (n1019 ? n924 : 1'b0) : (n437 ? (n1019 ? n924 : 1'b0) : n1019));
assign n3914 = /* LUT    2 10  7 */ (n304 ? 1'b0 : (n258 ? (n5 ? 1'b0 : !n142) : 1'b0));
assign n3915 = /* LUT   14 13  0 */ n45;
assign n3916 = /* LUT   22  2  4 */ (n2888 ? n2886 : (n2886 ? (n2890 ? n3011 : !n3011) : 1'b0));
assign n3917 = /* LUT    2  2  3 */ n188;
assign n3918 = /* LUT   21  6  7 */ n2610;
assign n3921 = /* LUT    5 15  2 */ (n601 ? 1'b0 : !n756);
assign n3922 = /* LUT   17 24  7 */ (n2297 ? (n2293 ? (n2298 ? !n2156 : 1'b0) : 1'b0) : 1'b0);
assign n3923 = /* LUT   17 16  3 */ n1325;
assign n3924 = /* LUT   11  4  7 */ (n1001 ? (n212 ? !n1539 : (n1539 ? !n1412 : 1'b1)) : (n212 ? 1'b1 : (n1539 ? !n1412 : 1'b1)));
assign n3925 = /* LUT    4 11  1 */ (n243 ? n249 : 1'b0);
assign n3926 = /* LUT   22  3  5 */ (n2762 ? 1'b0 : (n2765 ? 1'b0 : (n2763 ? 1'b0 : n2901)));
assign n3927 = /* LUT    2  3  4 */ n25;
assign n3928 = /* LUT    4 14  6 */ (n45 ? (n594 ? n128 : 1'b0) : (n594 ? n128 : (n128 ? n752 : 1'b0)));
assign n3931 = /* LUT   14 17  6 */ !n1636;
assign n3932 = /* LUT   14  9  2 */ n1789;
assign n3933 = /* LUT   15  5  0 */ n175;
assign n3934 = /* LUT    8  6  0 */ (n852 ? 1'b0 : n960);
assign n3935 = /* LUT   20 20  2 */ n2012;
assign n3936 = /* LUT    8  9  5 */ (n1150 ? (n1000 ? !n874 : n874) : (n1000 ? n874 : !n874));
assign n3937 = /* LUT   17  8  4 */ (n2350 ? (n2483 ? 1'b1 : !n2364) : (n2483 ? n2364 : 1'b0));
assign n3940 = /* LUT    9 22  5 */ (n1395 ? !n932 : n932);
assign n3941 = /* LUT    5  2  4 */ n177;
assign n3942 = /* LUT    9 14  1 */ (n1142 ? (n1351 ? 1'b0 : (n1017 ? !n1192 : 1'b1)) : (n1351 ? 1'b0 : !n1192));
assign n3943 = /* LUT    4  6  7 */ (n386 ? 1'b0 : !n538);
assign n3944 = /* LUT    8 10  6 */ (n1006 ? (n879 ? (n1134 ? 1'b0 : n1009) : 1'b0) : n879);
assign n3945 = /* LUT    8  2  2 */ (n823 ? (n176 ? n934 : 1'b0) : 1'b0);
assign n3946 = /* LUT    1 20  4 */ (n329 ? 1'b0 : (n143 ? (n150 ? n137 : 1'b0) : 1'b0));
assign n3947 = /* LUT   16 12  5 */ (n2103 ? (n1454 ? (n2382 ? 1'b1 : !n2238) : (n2382 ? n2238 : 1'b0)) : 1'b0);
assign n3948 = /* LUT   10 19  3 */ (n1381 ? (n1376 ? 1'b0 : (n277 ? 1'b1 : n930)) : (n1376 ? 1'b0 : n277));
assign n3949 = /* LUT    5  3  5 */ (n6 ? (n665 ? (n357 ? 1'b0 : !n41) : (n357 ? n41 : 1'b1)) : 1'b1);
assign n3950 = /* LUT    9 15  2 */ (n886 ? (n1353 ? 1'b0 : !n1194) : (n1353 ? 1'b0 : (n1194 ? n1137 : 1'b1)));
assign n3951 = /* LUT   18 21  2 */ (n2297 ? 1'b0 : (n2428 ? (n2156 ? n2293 : 1'b0) : 1'b0));
assign n3952 = /* LUT   17  4  6 */ n2310;
assign n3953 = /* LUT   23  3  7 */ !n3011;
assign n3954 = /* LUT   16 13  6 */ n1789;
assign n3955 = /* LUT   16  5  2 */ n189;
assign n3956 = /* LUT    3 20  2 */ (n628 ? (n643 ? 1'b0 : !n627) : (n468 ? 1'b0 : !n627));
assign n3957 = /* LUT   20  9  1 */ n1938;
assign n3958 = /* LUT   18 22  3 */ n2012;
assign n3959 = /* LUT    1 12  5 */ (n87 ? (n270 ? !n81 : 1'b0) : (n104 ? (n270 ? !n81 : 1'b0) : 1'b0));
assign n3960 = /* LUT    7  7  4 */ (n812 ? (n867 ? (n862 ? n865 : 1'b0) : (n862 ? 1'b0 : n865)) : (n867 ? (n862 ? !n865 : 1'b0) : (n862 ? 1'b0 : !n865)));
assign n3961 = /* LUT   12 22  6 */ (n1854 ? !n1665 : n1665);
assign n3962 = /* LUT   22 17  2 */ n2012;
assign n3965 = /* LUT   13 10  0 */ n1706;
assign n3966 = /* LUT   10  6  5 */ (n852 ? 1'b1 : !n980);
assign n3967 = /* LUT    9  2  4 */ (n956 ? 1'b0 : (n1239 ? !n1249 : (n1249 ? !n5 : 1'b1)));
assign n3968 = /* LUT    3 16  4 */ (n91 ? (n128 ? 1'b0 : n112) : n112);
assign n3969 = /* LUT   20  1  2 */ (n2759 ? !n2447 : n2447);
assign n3970 = /* LUT   12 15  3 */ (n1517 ? (n1645 ? n1608 : 1'b1) : 1'b1);
assign n3971 = /* LUT   20  4  7 */ !n2768;
assign n3972 = /* LUT   10  7  6 */ (n1271 ? n984 : (n5 ? (n1146 ? n984 : 1'b0) : n984));
assign n3976 = /* LUT   24 21  1 */ n2012;
assign n3980 = /* LUT   13 14  6 */ n45;
assign n3981 = /* LUT    2 21  7 */ (n112 ? !n159 : 1'b0);
assign n3982 = /* LUT   22 13  4 */ (n2395 ? 1'b0 : n3018);
assign n3983 = /* LUT    3 17  5 */ (n249 ? !n257 : 1'b0);
assign n3984 = /* LUT    3  9  1 */ (n569 ? (n566 ? n407 : !n407) : (n566 ? !n407 : n407));
assign n3985 = /* LUT   11 19  4 */ (n5 ? n1510 : (n1510 ? 1'b1 : (n1653 ? 1'b0 : n1508)));
assign n3986 = /* LUT   18 10  6 */ !n212;
assign n3987 = /* LUT    9  3  4 */ n189;
assign n3988 = /* LUT   18  2  2 */ (n2440 ? !n2441 : 1'b0);
assign n3989 = /* LUT   21 17  6 */ (n2156 ? (n2848 ? (n2293 ? 1'b0 : n2297) : 1'b0) : 1'b0);
assign n3990 = /* LUT   21  9  2 */ n2484;
assign n3991 = /* LUT   11 12  1 */ (n1474 ? 1'b0 : (n45 ? 1'b0 : (n1473 ? 1'b0 : !n1329)));
assign n3992 = /* LUT   13  6  7 */ n175;
assign n3993 = /* LUT    2  5  4 */ (n202 ? (n176 ? (n62 ? 1'b0 : !n375) : 1'b0) : !n62);
assign n3994 = /* LUT    3  1  2 */ (n345 ? (n6 ? (n41 ? !n339 : 1'b0) : 1'b1) : (n6 ? (n41 ? !n339 : 1'b1) : 1'b1));
assign n3995 = /* LUT   14 19  6 */ (n1647 ? n1813 : 1'b0);
assign n3996 = /* LUT   15 15  4 */ (n1624 ? (n212 ? (n2128 ? 1'b0 : n1790) : 1'b0) : 1'b0);
assign n3997 = /* LUT    3  4  7 */ (n41 ? (n6 ? !n356 : 1'b1) : (n6 ? 1'b1 : !n380));
assign n3998 = /* LUT   15  7  0 */ (n2064 ? (n2063 ? 1'b0 : (n2185 ? n2055 : 1'b0)) : 1'b0);
assign n3999 = /* LUT    7 21  1 */ n1070;
assign n4002 = /* LUT   22  5  4 */ !n2781;
assign n4003 = /* LUT    5 13  4 */ (n579 ? 1'b0 : (n580 ? (n113 ? !n271 : 1'b0) : 1'b0));
assign n4004 = /* LUT    4 17  7 */ (n448 ? (n612 ? 1'b0 : (n111 ? n299 : 1'b0)) : 1'b0);
assign n4005 = /* LUT    4  9  3 */ (n5 ? 1'b0 : n712);
assign n4006 = /* LUT   15  8  1 */ n1965;
assign n4009 = /* LUT   11  7  7 */ (n1576 ? (n841 ? 1'b1 : n1557) : (n841 ? 1'b0 : n1557));
assign n4010 = /* LUT   15 11  6 */ (n2238 ? (n2103 ? !n2110 : 1'b0) : (n2103 ? n1749 : 1'b0));
assign n4011 = /* LUT    2  6  4 */ (n394 ? (n51 ? 1'b0 : n222) : (n51 ? n222 : 1'b0));
assign n4012 = /* LUT    5 14  5 */ (n748 ? (n296 ? (n249 ? !n128 : 1'b0) : n249) : (n296 ? (n249 ? !n128 : 1'b0) : 1'b0));
assign n4013 = /* LUT   14 12  2 */ (n1770 ? 1'b0 : (n1452 ? !n2102 : 1'b1));
assign n4014 = /* LUT   17 12  0 */ n2248;
assign n4015 = /* LUT   15  4  3 */ n189;
assign n4016 = /* LUT   23 14  6 */ (n2970 ? (n3025 ? n3020 : (n3020 ? 1'b1 : n3024)) : (n3025 ? n3020 : (n3020 ? 1'b1 : !n3024)));
assign n4020 = /* LUT   15  3  7 */ n233;
assign n4021 = /* LUT   22  2  7 */ (n2887 ? 1'b0 : (n2892 ? 1'b0 : (n3011 ? 1'b0 : !n3010)));
assign n4022 = /* LUT   16 16  1 */ (n2272 ? !n1 : (n2274 ? (n2278 ? !n1 : 1'b0) : !n1));
assign n4023 = /* LUT    9 17  1 */ n1371;
assign n4024 = /* LUT   13 21  0 */ (n2021 ? (n1967 ? 1'b1 : !n1491) : n1967);
assign n4025 = /* LUT    7  9  4 */ (n1004 ? (n8 ? n999 : !n999) : (n8 ? !n999 : n999));
assign n4026 = /* LUT    8 13  6 */ (n1020 ? (n1019 ? (n1021 ? n907 : !n907) : 1'b0) : (n1019 ? 1'b0 : (n1021 ? n907 : !n907)));
assign n4027 = /* LUT    8  5  2 */ (n816 ? (n852 ? n1106 : 1'b0) : 1'b0);
assign n4028 = /* LUT   20 11  0 */ n2646;
assign n4031 = /* LUT   17  7  6 */ (n2345 ? (n2375 ? 1'b0 : !n2341) : 1'b0);
assign n4032 = /* LUT    7 10  5 */ (n1001 ? n892 : 1'b0);
assign n4033 = /* LUT    7  2  1 */ (n52 ? (n940 ? 1'b0 : !n200) : (n200 ? 1'b0 : !n838));
assign n4034 = /* LUT    9 21  7 */ (n233 ? n1031 : 1'b0);
assign n4035 = /* LUT    8  6  3 */ (n1122 ? (n973 ? n861 : 1'b0) : 1'b0);
assign n4036 = /* LUT    1 16  1 */ (n294 ? (n119 ? 1'b0 : n129) : (n119 ? n129 : 1'b0));
assign n4037 = /* LUT   16  8  2 */ n1789;
assign n4038 = /* LUT   20 20  5 */ (n2742 ? (n2290 ? n2404 : (n2404 ? n2403 : 1'b0)) : (n2290 ? (n2404 ? !n2403 : 1'b0) : 1'b0));
assign n4039 = /* LUT   20 12  1 */ (n2500 ? (n2809 ? !n2509 : 1'b0) : 1'b0);
assign n4040 = /* LUT   10 15  0 */ (n1459 ? n212 : (n1465 ? n212 : 1'b0));
assign n4041 = /* LUT   17  8  7 */ n1757;
assign n4044 = /* LUT    3 19  5 */ (n635 ? !n490 : n490);
assign n4045 = /* LUT    5  2  7 */ (n654 ? (n52 ? (n518 ? n497 : 1'b0) : 1'b0) : (n52 ? (n518 ? n497 : 1'b0) : n497));
assign n4046 = /* LUT    9 14  4 */ n177;
assign n4047 = /* LUT    2 20  1 */ (n150 ? (n93 ? n318 : 1'b0) : 1'b1);
assign n4052 = /* LUT    3 11  0 */ (n199 ? n128 : 1'b0);
assign n4053 = /* LUT    1 11  7 */ n45;
assign n4054 = /* LUT   12 18  3 */ n1640;
assign n4057 = /* LUT   10 10  6 */ (n931 ? n806 : 1'b0);
assign n4058 = /* LUT   10  2  2 */ (n1401 ? (n1398 ? (n6 ? !n41 : n41) : (n6 ? 1'b1 : n41)) : (n1398 ? (n6 ? !n41 : 1'b1) : 1'b1));
assign n4059 = /* LUT    9  6  5 */ (n967 ? (n1126 ? n1125 : 1'b0) : 1'b0);
assign n4060 = /* LUT   22 16  4 */ (n2293 ? 1'b0 : (n2156 ? 1'b0 : (n2297 ? 1'b0 : n2992)));
assign n4061 = /* LUT    2 16  3 */ (n294 ? 1'b0 : n129);
assign n4062 = /* LUT    3 20  5 */ (n631 ? (n479 ? n177 : (n177 ? 1'b1 : n637)) : (n479 ? 1'b0 : n637));
assign n4063 = /* LUT   13  9  2 */ n1592;
assign n4064 = /* LUT    3 12  1 */ (n258 ? (n283 ? (n434 ? 1'b0 : !n578) : 1'b0) : 1'b0);
assign n4065 = /* LUT   22  8  0 */ (n3015 ? !n1645 : 1'b0);
assign n4066 = /* LUT   21 20  7 */ (n2406 ? (n2864 ? (n2877 ? 1'b0 : n2403) : (n2877 ? !n2403 : 1'b1)) : 1'b0);
assign n4067 = /* LUT   21 12  3 */ (n2500 ? n2817 : 1'b0);
assign n4068 = /* LUT    1  4  4 */ (n41 ? (n6 ? n34 : 1'b1) : (n30 ? 1'b1 : n6));
assign n4069 = /* LUT   18 13  6 */ n2657;
assign n4070 = /* LUT   12 14  5 */ (n1781 ? 1'b0 : (n1792 ? (n1780 ? n1779 : 1'b0) : (n1780 ? 1'b0 : n1779)));
assign n4071 = /* LUT   18  5  2 */ n2453;
assign n4072 = /* LUT    2 17  4 */ (n257 ? (n249 ? !n158 : 1'b0) : (n132 ? (n249 ? !n158 : 1'b0) : 1'b0));
assign n4073 = /* LUT   13 10  3 */ n1730;
assign n4077 = /* LUT    9  2  7 */ (n176 ? 1'b0 : (n1088 ? n1096 : 1'b0));
assign n4078 = /* LUT   11 15  1 */ (n1483 ? n1364 : (n1488 ? 1'b1 : n1364));
assign n4079 = /* LUT   14 23  2 */ (n2162 ? (n2028 ? n1843 : !n1843) : (n2028 ? !n1843 : n1843));
assign n4082 = /* LUT   10  3  2 */ (n5 ? (n1410 ? 1'b1 : n1263) : (n1403 ? (n1410 ? 1'b1 : n1263) : (n1410 ? 1'b0 : n1263)));
assign n4083 = /* LUT   18  6  3 */ (n2612 ? !n2467 : n2467);
assign n4084 = /* LUT    3  7  7 */ n189;
assign n4085 = /* LUT   21 13  3 */ (n2964 ? !n2821 : n2821);
assign n4086 = /* LUT   12  6  6 */ (n1558 ? 1'b0 : (n1554 ? 1'b1 : (n1434 ? n1418 : !n1418)));
assign n4087 = /* LUT    5 16  4 */ (n212 ? (n252 ? (n304 ? !n422 : 1'b0) : !n422) : (n252 ? n304 : 1'b1));
assign n4088 = /* LUT    4 20  7 */ (n467 ? (n628 ? n647 : 1'b1) : (n628 ? n647 : n627));
assign n4089 = /* LUT   23 22  0 */ n2012;
assign n4090 = /* LUT    4 12  3 */ (n741 ? (n580 ? 1'b0 : n274) : (n580 ? n274 : 1'b0));
assign n4091 = /* LUT   14 15  3 */ (n1608 ? (n1563 ? (n1637 ? !n1609 : 1'b0) : 1'b0) : 1'b0);
assign n4092 = /* LUT    8 16  2 */ !n1043;
assign n4093 = /* LUT    2  4  6 */ (n37 ? !n194 : n194);
assign n4094 = /* LUT   22  4  7 */ !n2769;
assign n4095 = /* LUT   15 14  6 */ (n2117 ? (n1330 ? 1'b0 : n2116) : n2116);
assign n4096 = /* LUT    5 17  5 */ (n249 ? (n139 ? 1'b0 : n770) : 1'b0);
assign n4097 = /* LUT   15  6  2 */ (n2049 ? 1'b0 : (n1888 ? !n1463 : n1463));
assign n4098 = /* LUT    2  1  0 */ n175;
assign n4099 = /* LUT    5  9  1 */ (n5 ? (n564 ? 1'b0 : !n712) : (n564 ? (n712 ? 1'b0 : !n537) : !n712));
assign n4102 = /* LUT    4  5  0 */ (n371 ? (n529 ? 1'b1 : !n372) : (n388 ? !n372 : 1'b1));
assign n4103 = /* LUT    2  5  7 */ (n6 ? (n44 ? !n41 : 1'b1) : (n382 ? n41 : 1'b1));
assign n4104 = /* LUT   16 19  2 */ n2424;
assign n4105 = /* LUT   11  3  4 */ !n1416;
assign n4106 = /* LUT   14 11  5 */ (n2104 ? (n1705 ? 1'b0 : !n2102) : !n2102);
assign n4107 = /* LUT   15  7  3 */ (n1454 ? (n1885 ? 1'b0 : !n1699) : (n1885 ? !n1699 : 1'b0));
assign n4108 = /* LUT   20 22  5 */ (n2436 ? (n2404 ? 1'b1 : n2755) : (n2404 ? 1'b0 : n2755));
assign n4109 = /* LUT   22  5  7 */ (n2925 ? (n7 ? 1'b1 : n2911) : n7);
assign n4110 = /* LUT    5  1  2 */ (n494 ? (n498 ? n176 : 1'b0) : 1'b0);
assign n4111 = /* LUT    8  8  2 */ n188;
assign n4112 = /* LUT    5  4  7 */ (n680 ? (n41 ? (n6 ? 1'b0 : !n527) : 1'b0) : (n41 ? (n6 ? 1'b1 : !n527) : 1'b0));
assign n4113 = /* LUT   16 11  3 */ (n2366 ? (n2111 ? 1'b0 : !n2234) : 1'b0);
assign n4117 = /* LUT   17 10  6 */ (n1622 ? (n2507 ? n8 : !n8) : (n2507 ? !n8 : n8));
assign n4118 = /* LUT    7 13  5 */ (n711 ? 1'b1 : (n888 ? n564 : 1'b0));
assign n4119 = /* LUT   17  2  2 */ (n2304 ? (n2170 ? !n2333 : 1'b0) : n2170);
assign n4120 = /* LUT    7  5  1 */ (n362 ? n358 : (n358 ? (n679 ? 1'b0 : n808) : (n679 ? 1'b1 : n808)));
assign n4123 = /* LUT    1 19  1 */ (n141 ? (n135 ? 1'b0 : n150) : (n135 ? n150 : 1'b0));
assign n4124 = /* LUT    4  1  7 */ (n176 ? 1'b0 : (n649 ? n655 : 1'b0));
assign n4125 = /* LUT   20 15  1 */ n2012;
assign n4126 = /* LUT   14  3  5 */ (n1422 ? (n1290 ? 1'b0 : n2046) : n2046);
assign n4127 = /* LUT    8  4  4 */ n177;
assign n4128 = /* LUT   16  7  5 */ (n1542 ? (n1884 ? 1'b0 : !n2072) : (n1884 ? 1'b0 : n2072));
assign n4129 = /* LUT   20 18  6 */ (n2414 ? (n2406 ? n2849 : 1'b0) : (n2406 ? n2849 : (n2730 ? 1'b0 : n2849)));
assign n4130 = /* LUT   17  3  3 */ (n2318 ? (n2305 ? !n2333 : 1'b1) : 1'b0);
assign n4131 = /* LUT    7  6  2 */ (n698 ? 1'b0 : n970);
assign n4132 = /* LUT   10 13  1 */ (n1294 ? (n1340 ? (n1324 ? 1'b0 : n1336) : n1336) : (n1340 ? 1'b0 : n1336));
assign n4133 = /* LUT    9 17  4 */ n277;
assign n4134 = /* LUT    9  9  0 */ (n679 ? 1'b0 : (n907 ? !n806 : 1'b1));
assign n4135 = /* LUT    7  9  7 */ n854;
assign n4136 = /* LUT   13 20  7 */ n2012;
assign n4137 = /* LUT   13 12  3 */ (n1759 ? (n1494 ? 1'b0 : (n1762 ? n1939 : 1'b1)) : (n1494 ? 1'b0 : (n1762 ? n1939 : 1'b0)));
assign n4138 = /* LUT   20 11  3 */ n2642;
assign n4139 = /* LUT   18 16  1 */ n2411;
assign n4140 = /* LUT   20 10  7 */ n1789;
assign n4141 = /* LUT    3 18  7 */ (n142 ? (n130 ? n443 : (n443 ? n473 : 1'b0)) : (n130 ? n443 : 1'b0));
assign n4142 = /* LUT   22 20  0 */ 1'b1;
assign n4143 = /* LUT    9  1  1 */ (n1091 ? (n6 ? (n176 ? n41 : 1'b0) : n176) : n176);
assign n4144 = /* LUT    2 19  3 */ (n325 ? (n324 ? n331 : 1'b0) : 1'b0);
assign n4145 = /* LUT   13 13  4 */ n1953;
assign n4146 = /* LUT   22 19  4 */ (n2297 ? 1'b0 : (n2293 ? (n2992 ? !n2156 : 1'b0) : 1'b0));
assign n4147 = /* LUT    3 15  1 */ (n249 ? !n595 : 1'b0);
assign n4148 = /* LUT   21 15  3 */ n2012;
assign n4149 = /* LUT   11 18  2 */ n1518;
assign n4150 = /* LUT    1  7  4 */ !n226;
assign n4151 = /* LUT   12 17  5 */ n1635;
assign n4152 = /* LUT   18  8  2 */ (n2375 ? 1'b0 : (n2341 ? 1'b0 : (n577 ? n2377 : 1'b0)));
assign n4153 = /* LUT    2 20  4 */ (n134 ? n93 : 1'b0);
assign n4154 = /* LUT   12  9  1 */ (n1586 ? 1'b0 : (n1578 ? (n1580 ? 1'b0 : n1587) : 1'b0));
assign n4155 = /* LUT   22 12  1 */ (n2137 ? 1'b1 : n2663);
assign n4156 = /* LUT    2 12  0 */ n90;
assign n4157 = /* LUT   18 11  7 */ n2640;
assign n4158 = /* LUT   21  8  0 */ n2944;
assign n4159 = /* LUT    9  5  7 */ (n362 ? n841 : (n841 ? (n1113 ? 1'b1 : !n1111) : n1111));
assign n4160 = /* LUT    3 11  3 */ (n128 ? n87 : 1'b0);
assign n4161 = /* LUT   11 14  4 */ (n1484 ? (n1614 ? (n1343 ? !n1181 : 1'b0) : 1'b0) : (n1614 ? !n1181 : 1'b0));
assign n4162 = /* LUT   12 10  2 */ n179;
assign n4163 = /* LUT   10  2  5 */ n233;
assign n4164 = /* LUT   22 16  7 */ (n2156 ? (n2293 ? 1'b0 : (n2992 ? n2297 : 1'b0)) : 1'b0);
assign n4165 = /* LUT    5 19  4 */ (n466 ? 1'b0 : !n631);
assign n4166 = /* LUT   22  8  3 */ n2947;
assign n4167 = /* LUT   21 12  6 */ (n2509 ? !n2809 : 1'b0);
assign n4168 = /* LUT   21  4  2 */ (n2918 ? (n2914 ? !n8 : n8) : (n2914 ? n8 : !n8));
assign n4169 = /* LUT    4 15  3 */ (n756 ? 1'b0 : !n443);
assign n4172 = /* LUT    2  7  6 */ (n219 ? (n61 ? (n59 ? 1'b0 : n272) : 1'b0) : (n61 ? n272 : 1'b0));
assign n4173 = /* LUT    3  3  4 */ n233;
assign n4174 = /* LUT   11  6  5 */ (n1424 ? (n1125 ? 1'b0 : !n1126) : 1'b0);
assign n4175 = /* LUT   18  5  5 */ n2452;
assign n4176 = /* LUT    5 20  5 */ (n354 ? n631 : 1'b0);
assign n4177 = /* LUT   15  9  2 */ (n1595 ? n1465 : (n1465 ? (n1702 ? n1930 : !n1930) : 1'b0));
assign n4178 = /* LUT   23 20  7 */ n2012;
assign n4179 = /* LUT    5 12  1 */ (n62 ? n128 : 1'b0);
assign n4180 = /* LUT   17 21  6 */ (n2406 ? 1'b0 : (n2435 ? (n2433 ? 1'b0 : n2403) : (n2433 ? !n2403 : 1'b1)));
assign n4184 = /* LUT    8 20  3 */ (n925 ? 1'b1 : !n1064);
assign n4185 = /* LUT    2  8  7 */ !n238;
assign n4188 = /* LUT   16 22  2 */ (n2293 ? 1'b0 : (n2297 ? (n2428 ? !n2156 : 1'b0) : 1'b0));
assign n4192 = /* LUT   14 14  5 */ (n1454 ? (n2102 ? 1'b0 : !n1770) : !n1770);
assign n4193 = /* LUT   14  6  1 */ (n1877 ? (n1730 ? 1'b0 : !n1716) : (n1730 ? !n1716 : 1'b0));
assign n4194 = /* LUT   15 10  3 */ n1938;
assign n4195 = /* LUT   23 12  2 */ (n3051 ? !n2509 : n2509);
assign n4198 = /* LUT    5 16  7 */ (n252 ? (n151 ? n598 : 1'b0) : 1'b0);
assign n4199 = /* LUT    4 12  6 */ (n271 ? 1'b0 : n274);
assign n4200 = /* LUT   14 15  6 */ (n1650 ? !n1797 : n1797);
assign n4201 = /* LUT   17 14  2 */ (n2545 ? !n2391 : n2391);
assign n4204 = /* LUT   17 13  6 */ (n2541 ? !n2388 : n2388);
assign n4205 = /* LUT   20 21  7 */ (n2406 ? 1'b0 : (n2753 ? (n2749 ? 1'b0 : !n2403) : (n2749 ? n2403 : 1'b1)));
assign n4206 = /* LUT   20 13  3 */ (n2696 ? (n2707 ? n2705 : 1'b1) : !n2707);
assign n4207 = /* LUT    7  8  1 */ (n871 ? (n865 ? 1'b0 : n981) : (n865 ? n981 : 1'b0));
assign n4208 = /* LUT   14  7  1 */ (n1692 ? (n1904 ? 1'b0 : !n1718) : (n1904 ? 1'b0 : n1718));
assign n4209 = /* LUT    4  4  7 */ (n232 ? (n670 ? !n370 : 1'b1) : 1'b0);
assign n4210 = /* LUT    7 11  6 */ (n892 ? (n891 ? (n212 ? !n277 : 1'b0) : 1'b0) : 1'b0);
assign n4211 = /* LUT   13 23  2 */ (n2039 ? (n2032 ? n1842 : !n1842) : n2032);
assign n4212 = /* LUT   16 10  5 */ n2067;
assign n4213 = /* LUT   17  6  3 */ n2474;
assign n4214 = /* LUT   16  2  1 */ n177;
assign n4215 = /* LUT    9 20  4 */ (n1384 ? (n8 ? n1050 : !n1050) : (n8 ? !n1050 : n1050));
assign n4216 = /* LUT    5  1  5 */ (n502 ? (n503 ? n200 : 1'b1) : (n503 ? (n651 ? n200 : 1'b0) : (n651 ? 1'b1 : !n200)));
assign n4220 = /* LUT   18 19  2 */ (n2298 ? (n2297 ? (n2156 ? !n2293 : 1'b0) : 1'b0) : 1'b0);
assign n4221 = /* LUT    7 12  7 */ (n893 ? (n881 ? !n901 : 1'b0) : (n881 ? (n894 ? 1'b1 : !n901) : 1'b0));
assign n4222 = /* LUT    8  8  5 */ n179;
assign n4223 = /* LUT    7  4  3 */ (n679 ? (n652 ? n362 : !n362) : (n652 ? (n362 ? 1'b1 : n965) : (n362 ? 1'b0 : n965)));
assign n4224 = /* LUT   16 11  6 */ (n2364 ? (n2236 ? 1'b0 : n2355) : (n2355 ? !n2099 : 1'b0));
assign n4225 = /* LUT   16  3  2 */ n188;
assign n4226 = /* LUT   20 14  3 */ (n2838 ? (n2835 ? 1'b0 : (n2719 ? 1'b0 : !n2714)) : 1'b0);
assign n4227 = /* LUT   17  2  5 */ (n2309 ? 1'b1 : n2308);
assign n4228 = /* LUT    3 21  7 */ (n5 ? 1'b1 : (n485 ? 1'b0 : !n486));
assign n4229 = /* LUT    1  2  1 */ n12;
assign n4232 = /* LUT   13  8  0 */ n175;
assign n4233 = /* LUT   13 11  5 */ n1891;
assign n4234 = /* LUT    3 14  4 */ (n103 ? 1'b0 : !n288);
assign n4235 = /* LUT    1  6  7 */ n45;
assign n4236 = /* LUT   12 12  1 */ (n1767 ? (n1606 ? n1765 : !n1765) : (n1606 ? !n1765 : n1765));
assign n4237 = /* LUT   22 15  1 */ n3035;
assign n4238 = /* LUT    2 15  0 */ (n266 ? 1'b0 : (n151 ? !n142 : 1'b1));
assign n4239 = /* LUT   10  4  4 */ (n6 ? 1'b1 : (n41 ? !n1257 : !n1414));
assign n4240 = /* LUT    9  8  7 */ (n1124 ? (n1189 ? 1'b1 : n679) : (n1274 ? !n679 : 1'b0));
assign n4241 = /* LUT   21 11  0 */ n1757;
assign n4242 = /* LUT   22 18  6 */ n2012;
assign n4243 = /* LUT    1  3  1 */ (n24 ? (n23 ? (n190 ? n21 : 1'b0) : 1'b0) : 1'b0);
assign n4244 = /* LUT    2 18  5 */ (n158 ? 1'b0 : n112);
assign n4245 = /* LUT   13 12  6 */ (n1763 ? (n1632 ? 1'b0 : !n1037) : (n1632 ? n1037 : 1'b1));
assign n4246 = /* LUT   13  4  2 */ (n852 ? (n980 ? n1876 : n1674) : n1674);
assign n4247 = /* LUT   21 14  5 */ (n2836 ? (n2831 ? 1'b0 : !n2825) : (n2831 ? n2825 : 1'b1));
assign n4248 = /* LUT   11  9  0 */ (n212 ? 1'b0 : n1268);
assign n4249 = /* LUT   12 13  2 */ (n212 ? !n1607 : n1607);
assign n4250 = /* LUT   20  2  6 */ (io_19_0_1 ? (n2333 ? n2313 : 1'b0) : 1'b0);
assign n4251 = /* LUT   10  5  5 */ (n1248 ? (n1411 ? n1410 : 1'b1) : (n1411 ? (n5 ? n1410 : 1'b0) : (n5 ? 1'b1 : !n1410)));
assign n4252 = /* LUT    3  6  5 */ (n528 ? (n371 ? 1'b0 : (n207 ? 1'b0 : n176)) : (n371 ? 1'b1 : (n207 ? !n176 : 1'b1)));
assign n4253 = /* LUT   24 19  0 */ n2012;
assign n4254 = /* LUT    9  1  4 */ (n41 ? (n6 ? 1'b1 : !n951) : (n6 ? !n954 : 1'b1));
assign n4255 = /* LUT   15 20  7 */ (n2154 ? (n1652 ? !n2152 : 1'b1) : !n2152);
assign n4256 = /* LUT   22 19  7 */ (n2022 ? 1'b0 : (n2427 ? (n2426 ? 1'b0 : n2292) : 1'b0));
assign n4257 = /* LUT   22 11  3 */ (n2954 ? (n2952 ? !n2950 : 1'b0) : 1'b0);
assign n4258 = /* LUT    2 11  2 */ (n428 ? (n427 ? (n360 ? 1'b0 : n429) : 1'b0) : n427);
assign n4259 = /* LUT   21  7  2 */ n2941;
assign n4260 = /* LUT   11 10  1 */ (n1599 ? (n1458 ? 1'b0 : !n1451) : 1'b0);
assign n4261 = /* LUT    8 22  2 */ n1069;
assign n4262 = /* LUT   18  8  5 */ n1965;
assign n4263 = /* LUT    3  2  7 */ (n346 ? (n52 ? (n352 ? n168 : 1'b0) : 1'b1) : 1'b0);
assign n4264 = /* LUT    5 15  1 */ (n608 ? 1'b0 : (n752 ? 1'b0 : !n296));
assign n4265 = /* LUT   17 16  2 */ n1628;
assign n4266 = /* LUT    4 11  0 */ n737;
assign n4267 = /* LUT   22  3  4 */ (n3013 ? (n2889 ? !n2756 : n2897) : (n2889 ? !n2756 : !n2897));
assign n4268 = /* LUT    2  3  3 */ (n28 ? (n20 ? (n185 ? n19 : 1'b0) : 1'b0) : 1'b0);
assign n4269 = /* LUT    4 14  5 */ (n439 ? (n594 ? 1'b1 : n755) : 1'b0);
assign n4270 = /* LUT   14 17  5 */ (n5 ? 1'b1 : n1981);
assign n4271 = /* LUT    8 18  4 */ (n1057 ? (n334 ? (n648 ? !n620 : 1'b0) : 1'b0) : 1'b0);
assign n4272 = /* LUT   14  9  1 */ n1757;
assign n4273 = /* LUT   17 17  3 */ (n2011 ? n2410 : n2556);
assign n4274 = /* LUT   11  5  7 */ (n1126 ? (n212 ? (n1125 ? 1'b0 : !n1416) : 1'b0) : (n212 ? 1'b0 : (n1125 ? 1'b0 : n1416)));
assign n4279 = /* LUT    5 19  7 */ (n785 ? (n628 ? (n627 ? 1'b1 : n782) : n627) : 1'b0);
assign n4280 = /* LUT    5 11  3 */ (n814 ? (n732 ? 1'b0 : n764) : (n732 ? n764 : 1'b0));
assign n4281 = /* LUT    4 15  6 */ (n275 ? (n756 ? 1'b0 : (n594 ? 1'b1 : n132)) : !n756);
assign n4282 = /* LUT    4  7  2 */ n177;
assign n4283 = /* LUT   14 10  2 */ n1926;
assign n4284 = /* LUT    8 11  1 */ (n566 ? n811 : (n811 ? !n711 : 1'b0));
assign n4285 = /* LUT   15  9  5 */ (n1928 ? (n1731 ? 1'b0 : !n1890) : (n1731 ? !n1890 : 1'b0));
assign n4286 = /* LUT    1 20  3 */ (n146 ? (n148 ? 1'b0 : n80) : n80);
assign n4287 = /* LUT    5  4  0 */ (n531 ? (n681 ? 1'b0 : !n176) : !n176);
assign n4288 = /* LUT   10 19  2 */ (n188 ? n1031 : 1'b0);
assign n4289 = /* LUT    5  3  4 */ (n359 ? (n6 ? (n41 ? 1'b1 : !n380) : !n41) : (n6 ? (n41 ? 1'b1 : !n380) : 1'b1));
assign n4290 = /* LUT   16 14  1 */ (n1645 ? 1'b1 : (n1807 ? 1'b1 : n1));
assign n4291 = /* LUT   14  6  4 */ (n1882 ? 1'b0 : (n1714 ? !n1934 : n1934));
assign n4292 = /* LUT    8  3  2 */ (n679 ? (n5 ? 1'b1 : n659) : (n5 ? 1'b0 : !n836));
assign n4293 = /* LUT   16 13  5 */ n1938;
assign n4297 = /* LUT   20 17  4 */ n2012;
assign n4298 = /* LUT   20  9  0 */ (n2375 ? (n577 ? (n2341 ? 1'b0 : n2377) : 1'b0) : 1'b0);
assign n4299 = /* LUT   18 22  2 */ (n2403 ? (n2404 ? n2158 : 1'b0) : (n2404 ? n2592 : 1'b0));
assign n4302 = /* LUT    7  7  3 */ (n564 ? (n693 ? 1'b0 : (n5 ? 1'b0 : !n712)) : !n712);
assign n4303 = /* LUT    9 19  7 */ (n1189 ? (n1050 ? 1'b0 : (n931 ? !n932 : 1'b0)) : 1'b0);
assign n4304 = /* LUT   16  6  2 */ (n1453 ? (n1731 ? 1'b0 : !n1890) : (n1731 ? !n1890 : 1'b0));
assign n4305 = /* LUT   16  9  7 */ (n2366 ? 1'b0 : (n2351 ? (n2218 ? 1'b0 : !n2355) : (n2218 ? n2355 : 1'b1)));
assign n4306 = /* LUT   20 13  6 */ (n2500 ? !n2700 : (n2817 ? (n2544 ? 1'b1 : !n2700) : !n2700));
assign n4307 = /* LUT    7  8  4 */ (n993 ? (n868 ? 1'b0 : n981) : (n868 ? n981 : 1'b0));
assign n4308 = /* LUT   20 10  0 */ (n2375 ? 1'b0 : (n577 ? (n2377 ? n2341 : 1'b0) : 1'b0));
assign n4309 = /* LUT    2 21  6 */ (n155 ? n267 : 1'b0);
assign n4310 = /* LUT   13 14  5 */ (n1416 ? n1956 : !n1956);
assign n4311 = /* LUT    3 17  4 */ (n615 ? (n614 ? 1'b0 : n465) : 1'b0);
assign n4315 = /* LUT   18 19  5 */ (n2667 ? (n2430 ? !n2404 : (n2404 ? 1'b0 : n2403)) : (n2430 ? (n2404 ? 1'b0 : !n2403) : 1'b0));
assign n4316 = /* LUT   20  5  7 */ (n7 ? (n2673 ? (n2675 ? 1'b0 : !n2674) : 1'b0) : 1'b1);
assign n4317 = /* LUT    9 11  7 */ (n1320 ? (n1185 ? n984 : (n1146 ? n984 : 1'b0)) : 1'b0);
assign n4318 = /* LUT    4 22  0 */ (n803 ? !n488 : n488);
assign n4319 = /* LUT    9  3  3 */ (n1090 ? 1'b0 : (n200 ? !n1242 : 1'b0));
assign n4320 = /* LUT   13 15  6 */ n1786;
assign n4321 = /* LUT   13  7  2 */ (n1699 ? 1'b0 : (n1885 ? !n1593 : n1593));
assign n4322 = /* LUT   21 17  5 */ (n2404 ? (n2857 ? 1'b0 : n2403) : (n2403 ? !n2979 : 1'b0));
assign n4323 = /* LUT    3 10  1 */ n354;
assign n4324 = /* LUT   11 20  4 */ (n1520 ? (n5 ? 1'b1 : (n80 ? 1'b1 : n1501)) : (n5 ? 1'b1 : n1501));
assign n4325 = /* LUT   11 12  0 */ n1473;
assign n4326 = /* LUT    1  2  4 */ n13;
assign n4327 = /* LUT   18 11  0 */ n2634;
assign n4328 = /* LUT   10  8  5 */ (n1278 ? (n1436 ? 1'b0 : !n1132) : 1'b0);
assign n4329 = /* LUT    9  4  4 */ n177;
assign n4330 = /* LUT   22 22  7 */ (n2293 ? 1'b0 : (n2156 ? (n2297 ? 1'b0 : n2848) : 1'b0));
assign n4331 = /* LUT   22 14  3 */ (n3027 ? (n8 ? n3023 : !n3023) : (n8 ? !n3023 : n3023));
assign n4332 = /* LUT    2 14  2 */ (n271 ? 1'b0 : (n288 ? n113 : 1'b0));
assign n4333 = /* LUT   21 18  6 */ (n2156 ? 1'b0 : (n2986 ? (n2293 ? 1'b0 : !n2297) : 1'b0));
assign n4334 = /* LUT   21 10  2 */ n2625;
assign n4335 = /* LUT   11 16  6 */ (n1457 ? n1478 : 1'b0);
assign n4336 = /* LUT   12 12  4 */ (n1330 ? 1'b1 : (n1475 ? (n1473 ? n1474 : !n1474) : 1'b1));
assign n4337 = /* LUT   18  3  1 */ (n2066 ? n2601 : (n2342 ? !n1868 : n1868));
assign n4338 = /* LUT   12  4  0 */ (n852 ? n1419 : 1'b0);
assign n4339 = /* LUT    3  5  7 */ n188;
assign n4340 = /* LUT   15  8  0 */ (n1889 ? (n1597 ? 1'b0 : !n1903) : (n1597 ? !n1903 : 1'b0));
assign n4341 = /* LUT   22  7  0 */ !n2794;
assign n4342 = /* LUT   15 11  5 */ n1938;
assign n4343 = /* LUT    2  6  3 */ (n393 ? (n200 ? 1'b0 : n222) : (n200 ? n222 : 1'b0));
assign n4344 = /* LUT    5 14  4 */ (n128 ? n296 : 1'b0);
assign n4345 = /* LUT    8 21  4 */ (n158 ? 1'b0 : (n768 ? n249 : 1'b0));
assign n4346 = /* LUT   17 20  3 */ (n2410 ? (n2420 ? (n2426 ? n2022 : 1'b1) : (n2426 ? 1'b1 : n2022)) : (n2420 ? (n2426 ? 1'b0 : !n2022) : (n2426 ? !n2022 : 1'b0)));
assign n4347 = /* LUT   11  8  7 */ (n984 ? (n1577 ? 1'b1 : (n1146 ? 1'b1 : !n5)) : 1'b0);
assign n4348 = /* LUT   15 12  6 */ n2204;
assign n4349 = /* LUT   15  4  2 */ n354;
assign n4350 = /* LUT    4 18  6 */ n780;
assign n4351 = /* LUT    4 10  2 */ n179;
assign n4352 = /* LUT   14 13  2 */ (n2114 ? (n2123 ? (n2122 ? 1'b0 : !n2108) : 1'b1) : 1'b0);
assign n4353 = /* LUT    8 14  1 */ (n620 ? (n1025 ? (n910 ? n630 : !n630) : 1'b0) : (n1025 ? 1'b0 : (n910 ? n630 : !n630)));
assign n4354 = /* LUT    2  2  5 */ (n41 ? (n173 ? !n6 : 1'b1) : (n171 ? !n6 : 1'b1));
assign n4355 = /* LUT   22  2  6 */ (n2889 ? (n2757 ? !io_19_0_1 : 1'b0) : (n2757 ? !io_19_0_1 : n3008));
assign n4356 = /* LUT   16 16  0 */ (n2400 ? (n2272 ? (n1985 ? 1'b1 : n2270) : (n1985 ? !n2270 : 1'b0)) : (n1985 ? 1'b1 : n2270));
assign n4357 = /* LUT   14 16  7 */ (n1966 ? (n5 ? 1'b1 : !n1980) : (n5 ? 1'b0 : !n1980));
assign n4360 = /* LUT    5 15  4 */ (n441 ? 1'b0 : !n756);
assign n4361 = /* LUT   23 15  6 */ n2012;
assign n4362 = /* LUT    5  7  0 */ n175;
assign n4363 = /* LUT   23  7  2 */ (n1 ? 1'b1 : n3014);
assign n4364 = /* LUT   24  3  0 */ (n8 ? (n2901 ? n2894 : !n2894) : (n2901 ? !n2894 : n2894));
assign n4365 = /* LUT   22  3  7 */ (n2779 ? 1'b0 : (n2767 ? 1'b0 : (n2894 ? 1'b0 : !n2766)));
assign n4368 = /* LUT   16 17  1 */ (n1517 ? n2250 : (n1645 ? 1'b1 : n2250));
assign n4369 = /* LUT   14  9  4 */ n2067;
assign n4370 = /* LUT    8  6  2 */ (n1122 ? n1106 : 1'b0);
assign n4374 = /* LUT   20 20  4 */ (n2432 ? (n2156 ? 1'b0 : (n2297 ? !n2293 : 1'b0)) : 1'b0);
assign n4375 = /* LUT    8  9  7 */ n189;
assign n4376 = /* LUT   20 12  0 */ (n2697 ? (n2380 ? (n2704 ? 1'b0 : !n2705) : !n2704) : (n2380 ? !n2705 : 1'b1));
assign n4377 = /* LUT   17  8  6 */ n1755;
assign n4380 = /* LUT    9 22  7 */ (n437 ? (n1229 ? 1'b0 : n924) : (n1229 ? 1'b0 : (n924 ? 1'b1 : !n1069)));
assign n4381 = /* LUT    5  2  6 */ n15;
assign n4382 = /* LUT    9 14  3 */ n179;
assign n4385 = /* LUT    8  2  4 */ n15;
assign n4386 = /* LUT    1 20  6 */ (n150 ? (n137 ? (n144 ? !n329 : 1'b0) : 1'b0) : 1'b0);
assign n4387 = /* LUT   16 12  7 */ n1938;
assign n4388 = /* LUT   16  4  3 */ (n2173 ? (n2303 ? !n2182 : 1'b1) : 1'b0);
assign n4389 = /* LUT   10 19  5 */ (n1377 ? (n1210 ? (n1054 ? !n907 : 1'b0) : 1'b0) : 1'b0);
assign n4390 = /* LUT    7  3  0 */ n15;
assign n4391 = /* LUT   10 11  1 */ n1320;
assign n4392 = /* LUT    5  3  7 */ (n6 ? (n41 ? 1'b1 : !n359) : (n41 ? !n355 : 1'b1));
assign n4393 = /* LUT    9 15  4 */ (n477 ? (n1023 ? (n1021 ? n488 : !n488) : 1'b0) : (n1023 ? 1'b0 : (n1021 ? n488 : !n488)));
assign n4394 = /* LUT   16  5  4 */ (n2178 ? 1'b0 : (n2315 ? 1'b0 : !n1868));
assign n4395 = /* LUT   17  1  2 */ (n2439 ? 1'b0 : (n2314 ? 1'b0 : n2442));
assign n4396 = /* LUT    3 20  4 */ (n277 ? !n486 : 1'b0);
assign n4397 = /* LUT    3 12  0 */ !n113;
assign n4398 = /* LUT    1 12  7 */ (n247 ? (n267 ? n92 : 1'b1) : 1'b0);
assign n4399 = /* LUT   18 14  1 */ n2662;
assign n4400 = /* LUT    1  4  3 */ (n37 ? !n29 : n29);
assign n4401 = /* LUT   21 21  1 */ (n2403 ? (n2406 ? 1'b0 : !n2885) : (n2880 ? 1'b0 : !n2406));
assign n4402 = /* LUT   12 14  4 */ (n1605 ? (n1467 ? (n1619 ? n1618 : 1'b0) : (n1619 ? 1'b0 : n1618)) : (n1467 ? (n1619 ? !n1618 : 1'b0) : (n1619 ? 1'b0 : !n1618)));
assign n4403 = /* LUT   22 17  4 */ (n2297 ? (n2156 ? 1'b0 : (n2986 ? !n2293 : 1'b0)) : 1'b0);
assign n4404 = /* LUT    2 17  3 */ (n307 ? (n300 ? 1'b1 : (n267 ? n457 : 1'b0)) : 1'b0);
assign n4405 = /* LUT   13 10  2 */ n1750;
assign n4408 = /* LUT    9  2  6 */ (n6 ? (n969 ? !n41 : 1'b1) : (n968 ? n41 : 1'b1));
assign n4409 = /* LUT    1  5  4 */ n38;
assign n4410 = /* LUT   11 15  0 */ (n1504 ? (n1033 ? n1487 : 1'b0) : (n1033 ? (n1487 ? 1'b1 : n1355) : 1'b0));
assign n4411 = /* LUT   14 23  1 */ (n2161 ? (n2029 ? n1528 : !n1528) : (n2029 ? !n1528 : n1528));
assign n4412 = /* LUT    3 16  6 */ (n282 ? (n304 ? !n159 : (n159 ? 1'b0 : n611)) : 1'b0);
assign n4413 = /* LUT   20  1  4 */ (n2314 ? !n2595 : n2595);
assign n4414 = /* LUT   10  3  1 */ (n41 ? (n1407 ? !n6 : 1'b1) : (n1262 ? !n6 : 1'b1));
assign n4415 = /* LUT   12 15  5 */ (n1637 ? (n1608 ? 1'b0 : !n1609) : 1'b0);
assign n4416 = /* LUT   18  6  2 */ (n2611 ? !n2466 : n2466);
assign n4417 = /* LUT   12  7  1 */ (n1592 ? (n1429 ? 1'b0 : !n1135) : (n1429 ? 1'b0 : n1135));
assign n4418 = /* LUT   21 13  2 */ (n2963 ? !n2820 : n2820);
assign n4419 = /* LUT    4 21  2 */ (n798 ? !n777 : n777);
assign n4420 = /* LUT   18  9  7 */ (n2478 ? (n2364 ? n2355 : (n2355 ? n2221 : 1'b0)) : (n2364 ? 1'b0 : (n2355 ? n2221 : 1'b0)));
assign n4421 = /* LUT   15 20  0 */ (n1646 ? (n2021 ? (n1491 ? 1'b0 : !n5) : 1'b0) : !n5);
assign n4422 = /* LUT    3  9  3 */ (n571 ? (n567 ? n405 : !n405) : (n567 ? !n405 : n405));
assign n4423 = /* LUT    3  8  7 */ (n404 ? (n83 ? (n43 ? 1'b1 : n239) : 1'b0) : (n83 ? (n43 ? 1'b0 : n239) : 1'b0));
assign n4424 = /* LUT    9  3  6 */ (n1092 ? 1'b0 : (n200 ? 1'b0 : !n1085));
assign n4425 = /* LUT    5 17  4 */ (n252 ? (n763 ? !n304 : (n613 ? 1'b0 : !n304)) : 1'b0);
assign n4428 = /* LUT   11 12  3 */ n1474;
assign n4429 = /* LUT    2  5  6 */ n191;
assign n4430 = /* LUT    3  1  4 */ n189;
assign n4431 = /* LUT   11 11  7 */ (n1563 ? (n852 ? 1'b0 : n1564) : 1'b0);
assign n4432 = /* LUT   23 18  1 */ n2012;
assign n4433 = /* LUT   14 11  4 */ n1749;
assign n4434 = /* LUT   15 15  6 */ n2134;
assign n4435 = /* LUT   15  7  2 */ (n1678 ? !n2058 : (n1596 ? (n1573 ? !n2058 : 1'b0) : (n1573 ? 1'b0 : !n2058)));
assign n4436 = /* LUT    5 10  1 */ (n5 ? n728 : (n728 ? !n711 : 1'b0));
assign n4437 = /* LUT    7 21  3 */ (n177 ? n1031 : 1'b0);
assign n4440 = /* LUT   22  5  6 */ (n2457 ? 1'b1 : n2927);
assign n4441 = /* LUT    5 13  6 */ (n266 ? (n580 ? 1'b0 : (n579 ? 1'b0 : n581)) : 1'b0);
assign n4442 = /* LUT   21  1  5 */ (n2448 ? 1'b0 : (n2314 ? 1'b0 : (n2595 ? 1'b0 : !n2447)));
assign n4443 = /* LUT    4  9  5 */ (n711 ? 1'b0 : (n382 ? 1'b1 : !n559));
assign n4444 = /* LUT   15  8  3 */ (n1555 ? !n2074 : (n2074 ? 1'b0 : (n1930 ? n1698 : !n1698)));
assign n4445 = /* LUT   16 23  7 */ (n2156 ? 1'b0 : (n2293 ? 1'b0 : (n2297 ? n2296 : 1'b0)));
assign n4448 = /* LUT   17 11  1 */ (n2377 ? (n2375 ? 1'b0 : n577) : (n2375 ? n577 : 1'b0));
assign n4449 = /* LUT    7 14  0 */ (n304 ? (n905 ? 1'b0 : !n903) : 1'b0);
assign n4450 = /* LUT    2  6  6 */ (n39 ? (n200 ? (n26 ? !n374 : 1'b1) : 1'b0) : 1'b0);
assign n4451 = /* LUT   14 12  4 */ (n1772 ? 1'b0 : (n1730 ? !n1770 : 1'b1));
assign n4452 = /* LUT   14  4  0 */ (n1115 ? n852 : 1'b0);
assign n4456 = /* LUT    8 12  7 */ n177;
assign n4457 = /* LUT   10 21  4 */ (n1391 ? !n1519 : (n1367 ? !n1519 : 1'b1));
assign n4458 = /* LUT   10 13  0 */ (n1339 ? (n1304 ? (n1027 ? 1'b0 : !n1348) : 1'b0) : !n1348);
assign n4459 = /* LUT    9 17  3 */ (n490 ? (n1049 ? 1'b0 : !n1056) : (n1190 ? !n1056 : (n1049 ? 1'b0 : !n1056)));
assign n4460 = /* LUT   13 21  2 */ (n1657 ? (n2021 ? (n5 ? 1'b0 : n1491) : !n5) : 1'b0);
assign n4461 = /* LUT    7  9  6 */ !n812;
assign n4462 = /* LUT    8  5  4 */ (n5 ? (n1108 ? !n956 : 1'b0) : (n1108 ? n674 : 1'b1));
assign n4463 = /* LUT   21 23  1 */ n2012;
assign n4464 = /* LUT   20 19  6 */ n2012;
assign n4465 = /* LUT   20 11  2 */ n2643;
assign n4466 = /* LUT   10 14  1 */ (n1477 ? (n1459 ? n1268 : 1'b0) : n1459);
assign n4467 = /* LUT   18 24  4 */ (n2156 ? (n2297 ? (n2293 ? n2298 : 1'b0) : 1'b0) : 1'b0);
assign n4470 = /* LUT    9 10  0 */ (n811 ? (n565 ? 1'b1 : !n711) : 1'b0);
assign n4471 = /* LUT   16  8  4 */ (n2053 ? 1'b0 : (n1928 ? !n1914 : n1914));
assign n4472 = /* LUT   13 13  3 */ n1958;
assign n4473 = /* LUT   20 12  3 */ !n2133;
assign n4474 = /* LUT    3 19  7 */ (n139 ? 1'b0 : !n151);
assign n4475 = /* LUT   16  1  1 */ n2167;
assign n4476 = /* LUT    2 20  3 */ (n150 ? !n328 : 1'b0);
assign n4477 = /* LUT   10  9  7 */ (n721 ? (n1285 ? n1293 : 1'b0) : (n1285 ? (n1293 ? 1'b1 : n1131) : 1'b0));
assign n4478 = /* LUT    9  5  6 */ n175;
assign n4479 = /* LUT    1  8  4 */ (n237 ? 1'b0 : (n69 ? (n235 ? 1'b1 : n56) : n56));
assign n4480 = /* LUT    3 11  2 */ n74;
assign n4481 = /* LUT   11 14  3 */ (n1486 ? (n1356 ? (n1445 ? 1'b0 : !n1348) : 1'b1) : 1'b0);
assign n4482 = /* LUT   12 18  5 */ n1642;
assign n4483 = /* LUT   12 10  1 */ (n212 ? n1563 : 1'b0);
assign n4484 = /* LUT    2 13  0 */ (n117 ? n100 : 1'b0);
assign n4485 = /* LUT   10  2  4 */ (n1237 ? (n956 ? 1'b0 : !n1249) : (n5 ? (n956 ? 1'b0 : !n1249) : !n956));
assign n4486 = /* LUT    9  6  7 */ (n1126 ? (n1125 ? n973 : 1'b0) : 1'b0);
assign n4487 = /* LUT   22 16  6 */ (n2293 ? 1'b0 : (n2156 ? (n2986 ? n2297 : 1'b0) : 1'b0));
assign n4488 = /* LUT    2 16  5 */ (n452 ? n80 : (n129 ? 1'b0 : n80));
assign n4489 = /* LUT   13  9  4 */ (n1743 ? 1'b0 : (n1747 ? 1'b0 : (n1734 ? 1'b0 : !n1744)));
assign n4490 = /* LUT   22  8  2 */ (n1 ? 1'b0 : n3014);
assign n4491 = /* LUT    3 12  3 */ (n573 ? (n74 ? (n79 ? 1'b1 : n425) : (n79 ? n425 : 1'b0)) : n79);
assign n4492 = /* LUT   21 12  5 */ (n2720 ? (n2807 ? 1'b1 : (n2814 ? n2717 : 1'b0)) : (n2814 ? n2717 : 1'b0));
assign n4493 = /* LUT   21  4  1 */ (n2917 ? (n2915 ? !n8 : n8) : (n2915 ? n8 : !n8));
assign n4494 = /* LUT    1  4  6 */ (n37 ? !n40 : n40);
assign n4497 = /* LUT   12 14  7 */ (n5 ? 1'b0 : (n1620 ? !n1610 : 1'b1));
assign n4498 = /* LUT   18  5  4 */ n2451;
assign n4499 = /* LUT    5 20  4 */ (n631 ? n15 : 1'b0);
assign n4500 = /* LUT    2  9  2 */ n420;
assign n4501 = /* LUT   13  2  1 */ !n1868;
assign n4502 = /* LUT   11 15  3 */ (n264 ? !n5 : 1'b0);
assign n4503 = /* LUT   14 23  4 */ (n2164 ? (n8 ? n1848 : !n1848) : (n8 ? !n1848 : n1848));
assign n4504 = /* LUT    8 20  2 */ (n925 ? (n179 ? (n1206 ? 1'b1 : n1031) : n1206) : (n179 ? n1031 : 1'b0));
assign n4505 = /* LUT    2  8  6 */ (n83 ? 1'b1 : !n68);
assign n4508 = /* LUT   18  6  5 */ (n2614 ? !n2469 : n2469);
assign n4509 = /* LUT   15 10  2 */ (n2086 ? (n2089 ? (n1632 ? 1'b0 : n2088) : 1'b0) : (n2089 ? !n1632 : 1'b0));
assign n4510 = /* LUT   21  5  1 */ (n2930 ? (n8 ? n2777 : !n2777) : (n8 ? !n2777 : n2777));
assign n4511 = /* LUT   15 13  7 */ n1757;
assign n4512 = /* LUT    5 16  6 */ (n268 ? (io_4_31_0 ? (n766 ? n252 : 1'b0) : 1'b0) : 1'b0);
assign n4513 = /* LUT    4 12  5 */ (n743 ? (n582 ? 1'b0 : n274) : (n582 ? n274 : 1'b0));
assign n4514 = /* LUT   14 15  5 */ !n1968;
assign n4515 = /* LUT    8 16  4 */ !n1044;
assign n4516 = /* LUT   17 22  5 */ (n2404 ? 1'b0 : (n2403 ? n2299 : n2295));
assign n4517 = /* LUT   23 13  2 */ (n2960 ? 1'b1 : n2811);
assign n4518 = /* LUT   17 14  1 */ (n2394 ? !n2266 : n2266);
assign n4519 = /* LUT   11  2  5 */ n175;
assign n4520 = /* LUT    7 17  0 */ !n777;
assign n4521 = /* LUT    5 17  7 */ (n475 ? 1'b0 : (n767 ? !n772 : (n773 ? !n772 : 1'b0)));
assign n4522 = /* LUT   15  6  4 */ (n2065 ? (n2066 ? n2195 : !n1125) : (n2066 ? n2195 : n1125));
assign n4523 = /* LUT    2  1  2 */ n179;
assign n4524 = /* LUT    5  9  3 */ (n712 ? 1'b0 : (n410 ? !n564 : (n5 ? !n564 : 1'b1)));
assign n4525 = /* LUT    4 13  6 */ (n592 ? (n142 ? 1'b0 : (n434 ? !n280 : 1'b1)) : 1'b0);
assign n4526 = /* LUT    4  5  2 */ (n677 ? (n682 ? (n176 ? 1'b1 : n673) : n176) : (n682 ? (n176 ? 1'b0 : n673) : 1'b0));
assign n4527 = /* LUT   14  7  0 */ (n1692 ? (n1933 ? 1'b0 : !n1904) : (n1933 ? !n1904 : 1'b0));
assign n4528 = /* LUT   16 19  4 */ (n2425 ? (n2279 ? (n1823 ? n2146 : 1'b0) : (n1823 ? !n2146 : 1'b1)) : (n2279 ? (n1823 ? n2146 : 1'b1) : (n1823 ? !n2146 : 1'b0)));
assign n4529 = /* LUT   17 15  2 */ (n1 ? 1'b1 : n2272);
assign n4530 = /* LUT   11  3  6 */ (n5 ? n1249 : (n1401 ? n1249 : 1'b0));
assign n4531 = /* LUT   14 11  7 */ n1705;
assign n4532 = /* LUT   15  7  5 */ n2204;
assign n4533 = /* LUT   20 22  7 */ (n2752 ? (n2404 ? n2883 : 1'b1) : (n2404 ? n2883 : 1'b0));
assign n4534 = /* LUT   14  8  1 */ (n1926 ? (n1914 ? 1'b0 : !n2053) : (n1914 ? !n2053 : 1'b0));
assign n4535 = /* LUT    9 20  3 */ (n1383 ? (n1019 ? n8 : !n8) : (n1019 ? !n8 : n8));
assign n4536 = /* LUT    5  1  4 */ n175;
assign n4537 = /* LUT    7 12  6 */ (n582 ? (n1024 ? (n902 ? n581 : 1'b0) : (n902 ? !n581 : 1'b0)) : (n1024 ? (n902 ? 1'b0 : n581) : (n902 ? 1'b0 : !n581)));
assign n4538 = /* LUT    8  8  4 */ n354;
assign n4539 = /* LUT   16 11  5 */ (n2231 ? (n2355 ? (n2101 ? 1'b1 : n2364) : 1'b0) : (n2355 ? (n2101 ? !n2364 : 1'b0) : 1'b0));
assign n4542 = /* LUT   20 14  2 */ (n2837 ? (n8 ? n2821 : !n2821) : (n8 ? !n2821 : n2821));
assign n4543 = /* LUT   10 17  1 */ n189;
assign n4544 = /* LUT    9 13  0 */ (n698 ? 1'b0 : (n362 ? !n910 : 1'b1));
assign n4545 = /* LUT    7 13  7 */ (n679 ? (n621 ? !n362 : 1'b0) : !n362);
assign n4546 = /* LUT   17  2  4 */ (n2182 ? (n2313 ? 1'b0 : n2310) : n2310);
assign n4547 = /* LUT    7  5  3 */ (n843 ? (n698 ? (n680 ? 1'b1 : n5) : 1'b1) : (n698 ? (n680 ? 1'b1 : n5) : 1'b0));
assign n4548 = /* LUT    8  1  1 */ (n834 ? (n41 ? (n6 ? 1'b1 : !n825) : n6) : (n41 ? (n6 ? 1'b1 : !n825) : 1'b1));
assign n4551 = /* LUT    1 19  3 */ (n142 ? (n318 ? 1'b0 : n111) : 1'b0);
assign n4552 = /* LUT   14  3  7 */ (n807 ? n852 : 1'b0);
assign n4553 = /* LUT    8  4  6 */ (n971 ? (n961 ? !n1102 : 1'b0) : !n1102);
assign n4554 = /* LUT   16  7  7 */ (n1692 ? (n1923 ? 1'b0 : !n1904) : (n1923 ? !n1904 : 1'b0));
assign n4558 = /* LUT   17  3  5 */ (n2317 ? 1'b1 : n2322);
assign n4559 = /* LUT   10 21  7 */ (n1073 ? !n1389 : (n1389 ? n1069 : 1'b1));
assign n4560 = /* LUT   10 13  3 */ (n1459 ? (n1471 ? 1'b0 : (n1188 ? n1268 : 1'b1)) : 1'b0);
assign n4561 = /* LUT    9 17  6 */ !n932;
assign n4562 = /* LUT    9  9  2 */ (n1153 ? n1285 : (n1140 ? n1285 : (n1139 ? 1'b0 : n1285)));
assign n4563 = /* LUT   21 23  4 */ (n2293 ? (n2156 ? 1'b0 : (n2986 ? n2297 : 1'b0)) : 1'b0);
assign n4564 = /* LUT    1  3  0 */ n186;
assign n4565 = /* LUT   13 12  5 */ (n1770 ? 1'b0 : !n1772);
assign n4566 = /* LUT   13  4  1 */ n15;
assign n4567 = /* LUT   18 16  3 */ n2409;
assign n4568 = /* LUT   12 13  1 */ (n1783 ? (n1349 ? 1'b0 : n1776) : (n1625 ? !n1349 : 1'b0));
assign n4569 = /* LUT   10  5  4 */ n189;
assign n4570 = /* LUT    9  1  3 */ n354;
assign n4571 = /* LUT    2 19  5 */ (n307 ? (n93 ? n300 : 1'b0) : 1'b1);
assign n4572 = /* LUT   13 13  6 */ n1955;
assign n4573 = /* LUT   22 11  2 */ !n1645;
assign n4574 = /* LUT    2 11  1 */ (n82 ? 1'b1 : n260);
assign n4575 = /* LUT    3 15  3 */ (n435 ? (n142 ? 1'b0 : (n132 ? 1'b0 : !n288)) : 1'b0);
assign n4576 = /* LUT   22 19  6 */ (n2297 ? (n2156 ? (n2992 ? n2293 : 1'b0) : 1'b0) : 1'b0);
assign n4577 = /* LUT   21 15  5 */ (n2840 ? !n2818 : 1'b0);
assign n4578 = /* LUT   21  7  1 */ (n2794 ? (n2790 ? n2940 : !n2940) : (n2790 ? !n2940 : n2940));
assign n4579 = /* LUT    1  7  6 */ !n227;
assign n4580 = /* LUT   11 10  0 */ (n1146 ? 1'b0 : n1469);
assign n4581 = /* LUT   12 17  7 */ (n1636 ? (n1488 ? 1'b0 : (n1358 ? 1'b0 : !n1495)) : 1'b0);
assign n4582 = /* LUT   18  8  4 */ (n2375 ? (n2341 ? (n577 ? n2377 : 1'b0) : 1'b0) : 1'b0);
assign n4583 = /* LUT    2 20  6 */ (n249 ? (n329 ? !n80 : 1'b0) : 1'b1);
assign n4584 = /* LUT   12  9  3 */ (n1435 ? 1'b0 : (n1548 ? !n1593 : n1593));
assign n4585 = /* LUT    2 12  2 */ (n225 ? n100 : (n103 ? n100 : 1'b0));
assign n4586 = /* LUT   13  5  1 */ n177;
assign n4587 = /* LUT   21  8  2 */ n2948;
assign n4588 = /* LUT   14 18  0 */ (n1992 ? (n1999 ? (n2139 ? n1823 : 1'b0) : (n2139 ? 1'b1 : !n1823)) : (n1999 ? (n2139 ? !n1823 : 1'b1) : (n2139 ? 1'b0 : n1823)));
assign n4589 = /* LUT   11 14  6 */ (n1346 ? n1599 : (n1436 ? n1599 : (n1599 ? n1347 : 1'b0)));
assign n4590 = /* LUT   18  1  1 */ (n2314 ? (n8 ? n2595 : !n2595) : (n8 ? !n2595 : n2595));
assign n4591 = /* LUT    8 18  3 */ (n477 ? 1'b0 : (n620 ? 1'b0 : n1057));
assign n4592 = /* LUT   12  2  0 */ n1667;
assign n4593 = /* LUT   17 17  2 */ (n2555 ? (n2011 ? n2415 : 1'b1) : (n2011 ? n2415 : 1'b0));
assign n4596 = /* LUT    5 19  6 */ (n628 ? 1'b0 : !n627);
assign n4597 = /* LUT   22  8  5 */ (n2937 ? (n2801 ? n2803 : 1'b1) : 1'b1);
assign n4598 = /* LUT    5 11  2 */ (n813 ? (n730 ? 1'b0 : n764) : (n730 ? n764 : 1'b0));
assign n4599 = /* LUT   21  4  4 */ (n2920 ? (n8 ? !n2670 : n2670) : (n8 ? n2670 : !n2670));
assign n4600 = /* LUT    4 15  5 */ (n591 ? (n600 ? (n756 ? 1'b0 : n585) : !n756) : !n756);
assign n4601 = /* LUT    4  7  1 */ (n6 ? n696 : (n696 ? (n371 ? n52 : !n52) : !n52));
assign n4604 = /* LUT   14 10  1 */ n45;
assign n4605 = /* LUT    8 11  0 */ (n698 ? (n586 ? !n564 : 1'b0) : !n564);
assign n4606 = /* LUT   11  6  7 */ n233;
assign n4610 = /* LUT    5 20  7 */ (n627 ? (n621 ? (n628 ? !n646 : 1'b1) : (n628 ? n646 : 1'b1)) : (n621 ? (n628 ? !n646 : 1'b0) : (n628 ? n646 : 1'b1)));
assign n4611 = /* LUT   15  9  4 */ (n2084 ? (n2078 ? (n2071 ? !n2209 : 1'b0) : 1'b0) : 1'b0);
assign n4612 = /* LUT    5 12  3 */ (n817 ? (n749 ? !n580 : 1'b0) : (n749 ? n580 : 1'b0));
assign n4613 = /* LUT    4  8  2 */ (n713 ? (n396 ? n8 : !n8) : (n396 ? !n8 : n8));
assign n4614 = /* LUT   16 14  0 */ (n1766 ? n2128 : 1'b0);
assign n4615 = /* LUT   17 18  2 */ (n2569 ? !n2410 : n2410);
assign n4616 = /* LUT   14 14  7 */ (n1772 ? n1784 : (n1494 ? n1784 : n1959));
assign n4617 = /* LUT   15 10  5 */ (n2081 ? (n2098 ? (n1474 ? !n2060 : 1'b0) : !n2060) : (n2098 ? n1474 : 1'b1));
assign n4618 = /* LUT   14  6  3 */ (n1884 ? 1'b0 : (n1753 ? !n1542 : n1542));
assign n4619 = /* LUT   15  2  1 */ (n1649 ? (n1931 ? (n1874 ? 1'b0 : !n1863) : !n1874) : (n1931 ? !n1863 : 1'b1));
assign n4620 = /* LUT    1 21  3 */ (n337 ? (n157 ? !n154 : 1'b0) : (n157 ? n154 : 1'b0));
assign n4621 = /* LUT    5  5  0 */ (n6 ? (n41 ? !n527 : !n541) : 1'b1);
assign n4622 = /* LUT    7 16  2 */ !n334;
assign n4623 = /* LUT   16 15  1 */ n1629;
assign n4624 = /* LUT    9 19  6 */ (n1054 ? (n488 ? (n334 ? 1'b0 : !n490) : 1'b0) : 1'b0);
assign n4625 = /* LUT    1 14  0 */ (n107 ? (n80 ? 1'b1 : !n99) : !n99);
assign n4626 = /* LUT   10 20  1 */ (n179 ? (n354 ? (n15 ? n233 : 1'b0) : 1'b0) : 1'b0);
assign n4627 = /* LUT    8  7  7 */ !n865;
assign n4628 = /* LUT   17  5  4 */ n2325;
assign n4629 = /* LUT   20 13  5 */ (n2523 ? (n2814 ? (n2542 ? 1'b1 : n2720) : n2720) : (n2814 ? n2542 : 1'b0));
assign n4630 = /* LUT    7  8  3 */ (n992 ? (n867 ? 1'b0 : n981) : (n867 ? n981 : 1'b0));
assign n4631 = /* LUT   13 23  4 */ (n2041 ? (n2034 ? n1842 : !n1842) : n2034);
assign n4632 = /* LUT   16 10  7 */ (n1929 ? (n2364 ? n2087 : 1'b1) : (n2364 ? n2087 : 1'b0));
assign n4633 = /* LUT   17  6  5 */ n2475;
assign n4634 = /* LUT   16  2  3 */ n188;
assign n4635 = /* LUT   10 16  3 */ (n1370 ? 1'b0 : !n1459);
assign n4636 = /* LUT    9 20  6 */ (n1386 ? (n931 ? n8 : !n8) : (n931 ? !n8 : n8));
assign n4637 = /* LUT    5  1  7 */ (n6 ? (n41 ? !n492 : 1'b1) : (n41 ? !n496 : 1'b1));
assign n4638 = /* LUT    9 12  2 */ (n1332 ? (n1330 ? !n8 : (n8 ? n1329 : !n1329)) : (n1330 ? n8 : (n8 ? !n1329 : n1329)));
assign n4639 = /* LUT    7  4  5 */ (n950 ? (n955 ? (n679 ? 1'b1 : !n806) : n679) : (n955 ? !n679 : (n679 ? 1'b0 : n806)));
assign n4640 = /* LUT   13 15  5 */ (n1977 ? (n1805 ? (n1868 ? n1503 : !n1503) : (n1868 ? !n1503 : n1503)) : (n1805 ? (n1868 ? !n1503 : n1503) : (n1868 ? n1503 : !n1503)));
assign n4641 = /* LUT   20 14  5 */ n2661;
assign n4642 = /* LUT   20  6  1 */ (n2621 ? !n2677 : n2677);
assign n4643 = /* LUT   10  9  0 */ (n5 ? (n1267 ? n1435 : 1'b0) : n1267);
assign n4644 = /* LUT    1 10  7 */ n79;
assign n4645 = /* LUT   17  2  7 */ (n2182 ? (io_19_0_1 ? n2305 : 1'b0) : 1'b0);
assign n4646 = /* LUT    1  2  3 */ n16;
assign n4647 = /* LUT   10  8  4 */ (n5 ? (n1146 ? 1'b0 : n1291) : !n1146);
assign n4648 = /* LUT    9  4  3 */ (n1107 ? (n841 ? 1'b0 : (n1082 ? n1250 : 1'b1)) : (n841 ? 1'b0 : n1250));
assign n4649 = /* LUT    2 14  1 */ (n183 ? 1'b0 : (n5 ? 1'b0 : !n159));
assign n4650 = /* LUT   13  8  2 */ (n1567 ? (n1560 ? (n1721 ? n1582 : 1'b0) : 1'b0) : 1'b0);
assign n4651 = /* LUT   18 12  0 */ n2633;
assign n4652 = /* LUT   13 11  7 */ n1728;
assign n4653 = /* LUT   11 16  5 */ (n264 ? (n1514 ? (n1589 ? !n159 : 1'b0) : 1'b0) : (n1589 ? !n159 : 1'b0));
assign n4654 = /* LUT   10  1  1 */ n177;
assign n4655 = /* LUT   12 12  3 */ n1769;
assign n4656 = /* LUT   22 15  3 */ (n3036 ? (n8 ? n2973 : !n2973) : (n8 ? !n2973 : n2973));
assign n4657 = /* LUT    2 15  2 */ (n297 ? 1'b0 : (n199 ? 1'b0 : !n296));
assign n4658 = /* LUT   10  4  6 */ (n1078 ? (n1405 ? !n841 : 1'b0) : (n1405 ? !n841 : (n841 ? 1'b0 : n1107)));
assign n4659 = /* LUT    1  3  3 */ (n26 ? (n13 ? (n11 ? n27 : 1'b0) : (n11 ? !n27 : 1'b0)) : (n13 ? (n11 ? 1'b0 : n27) : (n11 ? 1'b0 : !n27)));
assign n4660 = /* LUT    2 18  7 */ (n264 ? 1'b0 : (n132 ? 1'b0 : (n142 ? 1'b0 : !n303)));
assign n4661 = /* LUT   14 21  0 */ !n2007;
assign n4662 = /* LUT   13  4  4 */ (n1872 ? (n1270 ? !n1422 : 1'b1) : 1'b0);
assign n4663 = /* LUT   21 14  7 */ (n2709 ? 1'b1 : n2815);
assign n4664 = /* LUT   11 17  6 */ (n1479 ? (n1639 ? 1'b0 : (n1369 ? 1'b1 : n212)) : (n1639 ? 1'b0 : (n1369 ? !n212 : 1'b0)));
assign n4665 = /* LUT   11  9  2 */ (n1446 ? !n1282 : 1'b0);
assign n4666 = /* LUT   12 13  4 */ (n1775 ? (n1783 ? !n1349 : (n1616 ? !n1349 : 1'b0)) : (n1783 ? 1'b0 : (n1616 ? !n1349 : 1'b0)));
assign n4667 = /* LUT   12  5  0 */ n177;
assign n4668 = /* LUT    3  6  7 */ (n6 ? (n530 ? 1'b0 : !n41) : (n530 ? (n41 ? n398 : 1'b0) : (n41 ? n398 : 1'b1)));
assign n4669 = /* LUT   10  5  7 */ (n1255 ? (n1265 ? 1'b1 : n956) : (n1265 ? !n956 : 1'b0));
assign n4670 = /* LUT    4 19  1 */ (n788 ? (n8 ? n334 : !n334) : (n8 ? !n334 : n334));
assign n4671 = /* LUT    9  1  6 */ (n1243 ? (n176 ? 1'b0 : n1240) : 1'b0);
assign n4672 = /* LUT   14 22  1 */ (n1848 ? 1'b0 : (n1843 ? 1'b0 : (n1847 ? 1'b0 : !n1845)));
assign n4673 = /* LUT    2 11  4 */ (n91 ? (n93 ? 1'b0 : (n132 ? 1'b0 : !n142)) : (n132 ? 1'b0 : !n142));
assign n4676 = /* LUT   21  7  4 */ n2942;
assign n4677 = /* LUT    8 14  0 */ (n1028 ? (n1043 ? (n1026 ? n1061 : !n1061) : 1'b0) : (n1043 ? 1'b0 : (n1026 ? n1061 : !n1061)));
assign n4678 = /* LUT   18  8  7 */ n2204;
assign n4679 = /* LUT    5 15  3 */ (n303 ? (n212 ? (n819 ? 1'b0 : n264) : n264) : 1'b0);
assign n4680 = /* LUT   17 16  4 */ (n2397 ? 1'b0 : n2395);
assign n4681 = /* LUT    4 11  2 */ (n391 ? 1'b0 : n248);
assign n4684 = /* LUT    2  3  5 */ (n193 ? (n180 ? n182 : 1'b0) : (n180 ? 1'b0 : n182));
assign n4685 = /* LUT   22  3  6 */ (n2899 ? (n2889 ? n2756 : n3006) : (n2889 ? n2756 : !n3006));
assign n4686 = /* LUT    4 14  7 */ (n151 ? 1'b0 : (n142 ? !n277 : 1'b0));
assign n4687 = /* LUT   16 17  0 */ (n2279 ? 1'b1 : (n2280 ? 1'b1 : !n1994));
assign n4688 = /* LUT    8 18  6 */ !n642;
assign n4689 = /* LUT   14  9  3 */ n1938;
assign n4690 = /* LUT   15  5  1 */ (n1701 ? 1'b0 : (n1679 ? !n1728 : n1728));
assign n4691 = /* LUT    5  8  0 */ (n559 ? (n711 ? 1'b0 : n371) : !n711);
assign n4692 = /* LUT   17 17  5 */ (n2011 ? n2411 : n2552);
assign n4695 = /* LUT   16 18  1 */ (n1997 ? (n2142 ? n1823 : !n1823) : (n2142 ? !n1823 : n1823));
assign n4696 = /* LUT    4  7  4 */ (n200 ? 1'b0 : n176);
assign n4697 = /* LUT   14 10  4 */ n1936;
assign n4698 = /* LUT   14  2  0 */ (n1125 ? (n967 ? (n1126 ? n852 : 1'b0) : 1'b0) : 1'b0);
assign n4699 = /* LUT   16 21  6 */ n2012;
assign n4703 = /* LUT   23  8  1 */ n2686;
assign n4704 = /* LUT   17  9  0 */ n2067;
assign n4705 = /* LUT    8 10  7 */ (n811 ? (n568 ? 1'b1 : !n711) : 1'b0);
assign n4706 = /* LUT    8  2  3 */ (n1079 ? (n945 ? n176 : 1'b0) : 1'b0);
assign n4707 = /* LUT    1 20  5 */ (n145 ? 1'b1 : (n329 ? 1'b1 : !n150));
assign n4708 = /* LUT   10 19  4 */ (n334 ? 1'b0 : (n5 ? 1'b0 : !n931));
assign n4709 = /* LUT   10 11  0 */ (n1471 ? 1'b0 : (n1459 ? (n1268 ? 1'b1 : n739) : 1'b0));
assign n4710 = /* LUT    5  3  6 */ (n510 ? (n200 ? 1'b1 : !n672) : (n513 ? (n200 ? 1'b1 : !n672) : (n200 ? 1'b0 : !n672)));
assign n4711 = /* LUT    9 15  3 */ (n984 ? (n1184 ? 1'b1 : n1146) : 1'b0);
assign n4712 = /* LUT   17  4  7 */ n2321;
assign n4713 = /* LUT   13 18  0 */ (n1991 ? (n1651 ? (n1503 ? n5 : 1'b0) : (n1503 ? 1'b1 : !n5)) : (n1651 ? (n1503 ? 1'b1 : !n5) : (n1503 ? n5 : 1'b0)));
assign n4714 = /* LUT    8  3  4 */ (n946 ? (n806 ? (n679 ? n826 : !n826) : (n679 ? n826 : 1'b1)) : (n806 ? (n679 ? n826 : !n826) : (n679 ? n826 : 1'b0)));
assign n4715 = /* LUT    1 21  6 */ (n157 ? !n156 : 1'b0);
assign n4716 = /* LUT   16 13  7 */ (n1790 ? 1'b0 : (n2254 ? n2251 : 1'b0));
assign n4717 = /* LUT   16  5  3 */ n15;
assign n4718 = /* LUT    1 13  2 */ (n279 ? (n99 ? !n95 : 1'b0) : (n99 ? n95 : 1'b0));
assign n4719 = /* LUT   17  1  1 */ (n2314 ? 1'b0 : (n2442 ? n2439 : 1'b0));
assign n4720 = /* LUT   20  9  2 */ n1757;
assign n4721 = /* LUT   18 22  4 */ (n2293 ? 1'b0 : (n2156 ? (n2296 ? !n2297 : 1'b0) : 1'b0));
assign n4722 = /* LUT   18 14  0 */ (n2274 ? !n1 : 1'b0);
assign n4723 = /* LUT   13 19  1 */ (n1822 ? !n1836 : n1836);
assign n4724 = /* LUT    7  7  5 */ (n550 ? (n849 ? 1'b0 : (n872 ? n856 : 1'b0)) : n872);
assign n4725 = /* LUT   21 21  0 */ n2012;
assign n4726 = /* LUT   16  6  4 */ (n1701 ? 1'b0 : (n1452 ? !n1679 : n1679));
assign n4727 = /* LUT   10 12  0 */ (n1268 ? n212 : 1'b0);
assign n4731 = /* LUT   17  5  7 */ n2328;
assign n4732 = /* LUT    1  5  3 */ (n30 ? !n45 : n45);
assign n4733 = /* LUT    3 16  5 */ (n607 ? (n249 ? (n80 ? !n303 : n303) : 1'b0) : (n249 ? (n80 ? 1'b0 : n303) : 1'b0));
assign n4734 = /* LUT   18 18  6 */ (n2576 ? (n2573 ? 1'b1 : !n2404) : (n2573 ? n2404 : 1'b0));
assign n4735 = /* LUT   12 15  4 */ (n1491 ? 1'b1 : !n1623);
assign n4736 = /* LUT   10  7  7 */ (n1431 ? n1268 : 1'b0);
assign n4739 = /* LUT   16  2  6 */ n15;
assign n4740 = /* LUT   13 14  7 */ (n1956 ? 1'b1 : n1416);
assign n4741 = /* LUT    3 17  6 */ (n316 ? !n456 : n456);
assign n4742 = /* LUT    3  9  2 */ (n570 ? (n409 ? n568 : !n568) : (n409 ? !n568 : n568));
assign n4743 = /* LUT   18 10  7 */ n1755;
assign n4744 = /* LUT    9  3  5 */ (n41 ? (n1095 ? n6 : 1'b1) : (n1255 ? n6 : 1'b1));
assign n4745 = /* LUT   12 11  6 */ n1434;
assign n4746 = /* LUT   13  7  4 */ (n1037 ? (n1716 ? !n1720 : (n1720 ? 1'b0 : !n1708)) : (n1716 ? 1'b1 : !n1708));
assign n4747 = /* LUT   21 17  7 */ n2012;
assign n4748 = /* LUT   11 20  6 */ (n1380 ? (n5 ? 1'b1 : (n80 ? 1'b1 : n1501)) : (n5 ? 1'b1 : n1501));
assign n4749 = /* LUT    1  2  6 */ n10;
assign n4750 = /* LUT   12  8  0 */ n15;
assign n4753 = /* LUT   10  8  7 */ (n1439 ? (n1284 ? (n705 ? !n1441 : 1'b1) : !n1441) : 1'b0);
assign n4754 = /* LUT    9  4  6 */ n233;
assign n4757 = /* LUT    2 14  4 */ (n128 ? (n5 ? 1'b1 : (n159 ? 1'b1 : n91)) : (n5 ? 1'b1 : n159));
assign n4758 = /* LUT   22  6  1 */ n2455;
assign n4759 = /* LUT   11 13  3 */ n179;
assign n4760 = /* LUT   21  2  0 */ (n2756 ? !n2889 : 1'b1);
assign n4764 = /* LUT   23 19  1 */ (n3040 ? (n3055 ? 1'b1 : !n2404) : (n3055 ? n2404 : 1'b0));
assign n4765 = /* LUT   12  4  2 */ (n852 ? n1563 : 1'b0);
assign n4766 = /* LUT   15  8  2 */ (n1925 ? (n2179 ? 1'b0 : !n2169) : (n2179 ? !n2169 : 1'b0));
assign n4767 = /* LUT   22  7  2 */ (n2684 ? (n2940 ? n2690 : (n2791 ? !n2690 : n2690)) : (n2940 ? !n2690 : (n2791 ? !n2690 : n2690)));
assign n4768 = /* LUT   17 19  4 */ n2578;
assign n4769 = /* LUT   15 11  7 */ n1754;
assign n4770 = /* LUT    2  6  5 */ (n395 ? (n52 ? 1'b0 : n222) : (n52 ? n222 : 1'b0));
assign n4771 = /* LUT    5 14  6 */ (n128 ? n608 : 1'b0);
assign n4772 = /* LUT    8 21  6 */ (n1221 ? (n1227 ? n1064 : (n1064 ? n925 : 1'b0)) : (n1227 ? (n1064 ? !n925 : 1'b0) : 1'b0));
assign n4773 = /* LUT   14 12  3 */ (n1750 ? (n1772 ? 1'b1 : (n1925 ? 1'b0 : n1770)) : (n1772 ? 1'b0 : (n1925 ? 1'b0 : n1770)));
assign n4774 = /* LUT   17 20  5 */ (n2427 ? (n2415 ? n2022 : 1'b0) : (n2415 ? 1'b1 : !n2022));
assign n4775 = /* LUT   17 12  1 */ (n2113 ? 1'b1 : (n2066 ? 1'b0 : n1807));
assign n4776 = /* LUT   15  4  4 */ (n1932 ? (n1875 ? 1'b0 : (n2051 ? n2048 : 1'b0)) : (n2051 ? n2048 : 1'b0));
assign n4777 = /* LUT   23 14  7 */ (n3018 ? 1'b0 : n3025);
assign n4778 = /* LUT    5  6  1 */ (n213 ? (n410 ? n8 : !n8) : (n410 ? !n8 : n8));
assign n4779 = /* LUT   14 13  4 */ (n1770 ? (n1772 ? 1'b0 : n1434) : !n1772);
assign n4780 = /* LUT    4  2  0 */ n233;
assign n4781 = /* LUT    8 14  3 */ (n1020 ? (n1026 ? (n621 ? n777 : 1'b0) : (n621 ? !n777 : 1'b0)) : (n1026 ? (n621 ? 1'b0 : n777) : (n621 ? 1'b0 : !n777)));
assign n4782 = /* LUT    2  2  7 */ n189;
assign n4783 = /* LUT   14  5  0 */ n354;
assign n4784 = /* LUT   16 16  2 */ (n2400 ? (n2270 ? 1'b0 : (n2272 ? 1'b0 : n2277)) : 1'b0);
assign n4785 = /* LUT   13 21  1 */ (n2021 ? (n5 ? 1'b0 : (n1491 ? n1655 : 1'b0)) : (n5 ? 1'b0 : n1655));
assign n4786 = /* LUT    8 13  7 */ (n1172 ? (n746 ? (n1167 ? 1'b0 : n1173) : 1'b1) : 1'b0);
assign n4789 = /* LUT    5  7  2 */ (n176 ? 1'b0 : !n200);
assign n4790 = /* LUT    4  3  1 */ (n516 ? (n506 ? (n41 ? !n6 : n6) : (n41 ? !n6 : 1'b1)) : (n506 ? (n41 ? 1'b1 : n6) : 1'b1));
assign n4793 = /* LUT   16 17  3 */ (n2279 ? (n1994 ? !n2280 : 1'b0) : 1'b0);
assign n4794 = /* LUT    7  2  2 */ (n679 ? n839 : (n837 ? (n806 ? !n839 : 1'b1) : (n806 ? !n839 : 1'b0)));
assign n4795 = /* LUT    8  6  4 */ (n861 ? (n852 ? 1'b0 : n973) : 1'b0);
assign n4796 = /* LUT    1 16  2 */ (n298 ? (n129 ? !n120 : 1'b0) : (n129 ? n120 : 1'b0));
assign n4797 = /* LUT   20 20  6 */ (n2293 ? (n2296 ? (n2297 ? n2156 : 1'b0) : 1'b0) : 1'b0);
assign n4798 = /* LUT   10 15  1 */ (n1495 ? !n984 : 1'b0);
assign n4799 = /* LUT   13 22  1 */ (n1491 ? 1'b0 : n1527);
assign n4802 = /* LUT    9 14  5 */ n354;
assign n4803 = /* LUT    8  2  6 */ (n936 ? (n1094 ? (n1093 ? 1'b1 : !n941) : 1'b0) : (n1093 ? 1'b1 : !n941));
assign n4804 = /* LUT   16  4  5 */ (n2333 ? (n2303 ? 1'b0 : n2172) : n2172);
assign n4805 = /* LUT   12 19  0 */ (n1652 ? !n1639 : 1'b0);
assign n4806 = /* LUT    7  3  2 */ n179;
assign n4807 = /* LUT   10 11  3 */ (n1316 ? (n1309 ? 1'b0 : n1456) : (n1309 ? (n1315 ? 1'b0 : n1456) : n1456));
assign n4808 = /* LUT   16  5  6 */ (n1453 ? (n1884 ? 1'b0 : !n1542) : (n1884 ? 1'b0 : n1542));
assign n4809 = /* LUT    2 16  4 */ (n294 ? 1'b0 : (n293 ? (n452 ? !n252 : 1'b0) : 1'b0));
assign n4810 = /* LUT    3 20  6 */ (n628 ? !n481 : (n627 ? 1'b1 : !n471));
assign n4811 = /* LUT   13  9  3 */ (n1751 ? (n1595 ? 1'b0 : !n1702) : (n1595 ? 1'b0 : n1702));
assign n4812 = /* LUT    3 12  2 */ (n128 ? 1'b1 : !n274);
assign n4813 = /* LUT   18 14  3 */ (n1 ? 1'b1 : n2274);
assign n4814 = /* LUT    1  4  5 */ (n27 ? (n41 ? 1'b1 : (n6 ? n29 : 1'b1)) : (n41 ? n6 : (n6 ? n29 : 1'b1)));
assign n4818 = /* LUT   12 14  6 */ (n1622 ? 1'b0 : n1623);
assign n4819 = /* LUT   22 17  6 */ (n2297 ? 1'b0 : (n2156 ? 1'b0 : (n2855 ? !n2293 : 1'b0)));
assign n4820 = /* LUT    2 17  5 */ (n124 ? (n295 ? n268 : 1'b0) : n268);
assign n4821 = /* LUT   13 10  4 */ n1753;
assign n4822 = /* LUT    2  9  1 */ (n209 ? !n208 : n208);
assign n4825 = /* LUT   13  2  0 */ n1862;
assign n4826 = /* LUT   11 15  2 */ (n1356 ? (n1498 ? (n1499 ? !n1333 : 1'b0) : n1499) : (n1498 ? 1'b0 : n1499));
assign n4827 = /* LUT    1  5  6 */ (n38 ? (n41 ? n6 : (n6 ? 1'b1 : !n40)) : (n41 ? 1'b1 : (n6 ? 1'b1 : !n40)));
assign n4828 = /* LUT   14 23  3 */ (n2163 ? (n2026 ? n1845 : !n1845) : (n2026 ? !n1845 : n1845));
assign n4831 = /* LUT   10  3  3 */ (n1404 ? (n1091 ? 1'b1 : !n1107) : (n1091 ? !n1246 : (n1107 ? 1'b0 : !n1246)));
assign n4832 = /* LUT   12 15  7 */ (n1181 ? 1'b0 : (n1633 ? (n1354 ? 1'b1 : !n1492) : 1'b0));
assign n4833 = /* LUT   18  6  4 */ (n2613 ? !n2468 : n2468);
assign n4834 = /* LUT   12  7  3 */ n354;
assign n4835 = /* LUT   13  3  1 */ (n1553 ? (n1417 ? 1'b0 : !n1874) : !n1417);
assign n4836 = /* LUT   21 13  4 */ (n2825 ? n2833 : n2962);
assign n4839 = /* LUT   21  5  0 */ (n2924 ? (n8 ? n2776 : !n2776) : (n8 ? !n2776 : n2776));
assign n4840 = /* LUT    8 16  3 */ !n931;
assign n4841 = /* LUT   21  6  1 */ n2606;
assign n4842 = /* LUT   18  2  6 */ n2311;
assign n4843 = /* LUT   15 14  7 */ (n2126 ? (n1473 ? 1'b1 : (n1494 ? 1'b0 : !n2117)) : (n1473 ? n1494 : 1'b0));
assign n4844 = /* LUT    5  9  2 */ (n811 ? (n711 ? (n565 ? 1'b0 : n5) : 1'b1) : 1'b0);
assign n4845 = /* LUT    4 13  5 */ (n751 ? (n575 ? (n266 ? !n744 : 1'b0) : n266) : 1'b0);
assign n4846 = /* LUT   11  4  1 */ (n1406 ? 1'b0 : (n212 ? !n1550 : 1'b1));
assign n4847 = /* LUT    4  5  1 */ n354;
assign n4848 = /* LUT    3  1  6 */ n175;
assign n4851 = /* LUT   17 15  1 */ !n2275;
assign n4852 = /* LUT   11  3  5 */ (n1407 ? (n1410 ? 1'b0 : n1399) : (n5 ? (n1410 ? 1'b0 : n1399) : n1399));
assign n4853 = /* LUT   14 11  6 */ (n423 ? 1'b1 : n577);
assign n4857 = /* LUT   15  7  4 */ (n2087 ? (n1876 ? 1'b0 : !n1691) : (n1876 ? !n1691 : 1'b0));
assign n4858 = /* LUT   23 17  7 */ (n3053 ? (n2404 ? !n3054 : 1'b0) : (n2404 ? !n3054 : 1'b1));
assign n4859 = /* LUT    5 10  3 */ (n63 ? (n711 ? 1'b0 : n811) : n811);
assign n4860 = /* LUT    7 21  5 */ (n5 ? (n159 ? 1'b0 : n249) : (n485 ? 1'b0 : (n159 ? 1'b0 : n249)));
assign n4863 = /* LUT   14  8  0 */ (n1920 ? (n1723 ? 1'b0 : (n1921 ? n1899 : 1'b0)) : 1'b0);
assign n4864 = /* LUT    4  9  7 */ (n565 ? !n406 : n406);
assign n4865 = /* LUT   15  8  5 */ (n1909 ? (n1932 ? 1'b0 : !n1929) : (n1932 ? 1'b0 : n1929));
assign n4868 = /* LUT   17 11  3 */ (n2355 ? 1'b0 : (n2499 ? (n2364 ? 1'b0 : !n2244) : (n2364 ? 1'b1 : !n2244)));
assign n4872 = /* LUT    4  6  1 */ n233;
assign n4873 = /* LUT    7 14  2 */ (n1033 ? (n904 ? 1'b1 : (n818 ? n1046 : 1'b0)) : (n818 ? n1046 : 1'b0));
assign n4874 = /* LUT   16 20  3 */ (n2154 ? 1'b0 : !n2155);
assign n4875 = /* LUT    7 13  6 */ (n698 ? (n610 ? !n564 : 1'b0) : !n564);
assign n4876 = /* LUT   14 12  6 */ (n1772 ? n1752 : (n1934 ? 1'b0 : n1770));
assign n4877 = /* LUT   14  4  2 */ (n1698 ? (n1679 ? (n1410 ? 1'b0 : !n956) : !n956) : (n1679 ? !n1410 : 1'b1));
assign n4878 = /* LUT    8  1  0 */ n15;
assign n4879 = /* LUT    1 19  2 */ (n326 ? (n136 ? 1'b0 : n150) : (n136 ? n150 : 1'b0));
assign n4882 = /* LUT    8  4  5 */ (n972 ? (n1107 ? n966 : 1'b1) : (n1107 ? (n966 ? !n1087 : 1'b0) : !n1087));
assign n4883 = /* LUT   20 18  7 */ (n2731 ? n2565 : (n2588 ? n2565 : (n2406 ? 1'b0 : n2565)));
assign n4884 = /* LUT   17  3  4 */ (io_19_0_1 ? (n2333 ? n2304 : 1'b0) : 1'b0);
assign n4885 = /* LUT   10 13  2 */ (n212 ? (n1146 ? 1'b1 : n1479) : 1'b0);
assign n4886 = /* LUT    9 17  5 */ (n277 ? (n1202 ? (n1201 ? n1200 : !n1200) : 1'b0) : (n1202 ? 1'b0 : (n1201 ? n1200 : !n1200)));
assign n4887 = /* LUT    9  9  1 */ (n811 ? n1146 : (n1146 ? !n876 : 1'b0));
assign n4888 = /* LUT   13 21  4 */ (n2025 ? (n1652 ? n1665 : 1'b0) : n1652);
assign n4889 = /* LUT    8  5  6 */ (n971 ? (n1109 ? 1'b0 : n969) : !n1109);
assign n4893 = /* LUT   20 11  4 */ n2635;
assign n4894 = /* LUT   10 14  3 */ n1342;
assign n4897 = /* LUT    9 10  2 */ (n1143 ? n1007 : (n1007 ? !n1152 : 1'b0));
assign n4898 = /* LUT   22 20  1 */ n2012;
assign n4899 = /* LUT    7  2  5 */ (n949 ? n200 : (n52 ? n200 : (n200 ? n943 : 1'b0)));
assign n4900 = /* LUT   21 16  0 */ (n2845 ? (n2844 ? !n2403 : (n2978 ? !n2403 : 1'b1)) : (n2844 ? 1'b0 : (n2978 ? 1'b0 : n2403)));
assign n4901 = /* LUT   16  8  6 */ (n1679 ? (n1701 ? !n2203 : (n1927 ? !n2203 : 1'b0)) : (n1701 ? !n2203 : (n1927 ? 1'b0 : !n2203)));
assign n4902 = /* LUT   13 13  5 */ n1954;
assign n4903 = /* LUT    3 15  2 */ (n280 ? 1'b0 : (n438 ? 1'b0 : (n303 ? !n442 : 1'b0)));
assign n4904 = /* LUT   20  4  1 */ !n2772;
assign n4905 = /* LUT   18 17  3 */ (n2156 ? (n2293 ? 1'b0 : (n2297 ? 1'b0 : n2432)) : 1'b0);
assign n4906 = /* LUT    1  7  5 */ !n53;
assign n4907 = /* LUT   12 17  6 */ n1637;
assign n4908 = /* LUT    2 20  5 */ (n306 ? n93 : 1'b0);
assign n4909 = /* LUT   22 12  2 */ (n2814 ? 1'b1 : n2395);
assign n4910 = /* LUT    2 12  1 */ (n255 ? (n256 ? (n261 ? 1'b1 : !n112) : 1'b1) : (n256 ? !n112 : 1'b1));
assign n4911 = /* LUT   13  5  0 */ (n956 ? (n1696 ? 1'b0 : !n841) : !n841);
assign n4914 = /* LUT    1  8  6 */ (n214 ? (n8 ? n60 : !n60) : (n8 ? !n60 : n60));
assign n4915 = /* LUT   11 14  5 */ (n984 ? 1'b0 : (n4 ? n1563 : 1'b0));
assign n4916 = /* LUT   12 18  7 */ (n1647 ? 1'b0 : n1813);
assign n4917 = /* LUT    2 13  2 */ (n112 ? (n431 ? (n243 ? !n81 : 1'b0) : 1'b0) : 1'b0);
assign n4918 = /* LUT   13  6  1 */ (n1632 ? (n1891 ? !n1877 : (n1037 ? n1877 : !n1877)) : (n1891 ? (n1037 ? !n1877 : n1877) : n1877));
assign n4919 = /* LUT   10  2  6 */ (n41 ? (n6 ? 1'b1 : !n1247) : (n6 ? 1'b1 : !n1248));
assign n4920 = /* LUT    4 16  0 */ (n455 ? (n606 ? 1'b0 : n249) : (n606 ? 1'b0 : (n117 ? n249 : 1'b0)));
assign n4921 = /* LUT    2 16  7 */ (n252 ? n452 : (n293 ? 1'b0 : n452));
assign n4922 = /* LUT   13  9  6 */ (n1699 ? 1'b0 : (n1732 ? !n1885 : n1885));
assign n4926 = /* LUT    3 12  5 */ (n584 ? !n125 : 1'b0);
assign n4927 = /* LUT   21 12  7 */ (n2809 ? (n2522 ? !n2509 : 1'b0) : (n2522 ? (n2535 ? n2509 : 1'b0) : 1'b0));
assign n4928 = /* LUT   22  8  4 */ (n3014 ? (n2947 ? !n2693 : 1'b0) : 1'b0);
assign n4929 = /* LUT    3  4  1 */ (n52 ? n51 : (n526 ? (n369 ? 1'b0 : n51) : 1'b0));
assign n4930 = /* LUT   21  4  3 */ (n2919 ? (n2912 ? !n8 : n8) : (n2912 ? n8 : !n8));
assign n4938 = /* LUT   18  5  6 */ n2450;
assign n4939 = /* LUT    5 20  6 */ (n785 ? (n640 ? (n792 ? n795 : 1'b1) : n795) : n795);
assign n4940 = /* LUT   17 21  7 */ (n2426 ? (n2022 ? 1'b0 : (n2292 ? 1'b0 : n2427)) : 1'b0);
assign n4941 = /* LUT   11 15  5 */ (n1599 ? (n1357 ? 1'b1 : (n1436 ? 1'b1 : n1363)) : 1'b0);
assign n4942 = /* LUT   11  7  1 */ (n1432 ? n1564 : (n816 ? (n841 ? n1564 : 1'b0) : 1'b0));
assign n4943 = /* LUT    8 20  4 */ (n925 ? (n1043 ? n930 : (n1064 ? 1'b1 : n930)) : n930);
assign n4946 = /* LUT   17 18  1 */ (n2415 ? !n2409 : n2409);
assign n4947 = /* LUT   14 14  6 */ (n1463 ? n2102 : 1'b0);
assign n4948 = /* LUT   15 10  4 */ (n2098 ? 1'b0 : (n2091 ? !n2210 : 1'b1));
assign n4949 = /* LUT   15  2  0 */ n175;
assign n4950 = /* LUT    7 16  1 */ n1051;
assign n4951 = /* LUT   16 15  0 */ n1321;
assign n4952 = /* LUT   14 15  7 */ (n1651 ? (n1798 ? (n1812 ? n1796 : !n1796) : 1'b0) : (n1798 ? 1'b0 : (n1812 ? n1796 : !n1796)));
assign n4953 = /* LUT    8 16  6 */ !n1061;
assign n4954 = /* LUT   15  3  1 */ n175;
assign n4955 = /* LUT   17 14  3 */ (n2546 ? !n2392 : n2392);
assign n4956 = /* LUT    7 17  2 */ (n5 ? 1'b0 : (n302 ? (n131 ? n448 : 1'b0) : 1'b0));
assign n4957 = /* LUT   15  6  6 */ (n1728 ? (n1689 ? 1'b0 : !n1887) : (n1689 ? 1'b0 : n1887));
assign n4958 = /* LUT    2  1  4 */ (n161 ? (n176 ? n41 : (n164 ? 1'b1 : !n41)) : (n176 ? n41 : (n164 ? n41 : 1'b0)));
assign n4959 = /* LUT    5  9  5 */ (n711 ? (n568 ? 1'b0 : (n5 ? n811 : 1'b0)) : n811);
assign n4960 = /* LUT    4  5  4 */ (n212 ? !n101 : (n52 ? !n101 : (n101 ? 1'b0 : !n378)));
assign n4961 = /* LUT   14  7  2 */ (n1889 ? (n1452 ? 1'b0 : !n1903) : (n1452 ? !n1903 : 1'b0));
assign n4962 = /* LUT   16 19  6 */ (n2286 ? (n2145 ? (n1823 ? n2280 : !n2280) : !n2280) : (n2145 ? n2280 : (n1823 ? !n2280 : n2280)));
assign n4963 = /* LUT   13 23  3 */ (n2040 ? (n2033 ? n1842 : !n1842) : n2033);
assign n4966 = /* LUT    1 18  5 */ (n307 ? (n130 ? n93 : 1'b0) : 1'b1);
assign n4969 = /* LUT   10 16  2 */ (n1459 ? (n1367 ? n1268 : 1'b1) : 1'b0);
assign n4970 = /* LUT    9 20  5 */ (n1385 ? (n8 ? n1189 : !n1189) : (n8 ? !n1189 : n1189));
assign n4971 = /* LUT    9 12  1 */ (n817 ? (n1322 ? n8 : !n8) : (n1322 ? !n8 : n8));
assign n4972 = /* LUT   13 16  0 */ (n1126 ? n1983 : !n1983);
assign n4973 = /* LUT    7  4  4 */ n175;
assign n4974 = /* LUT    8  8  6 */ !n866;
assign n4975 = /* LUT   16 11  7 */ n1938;
assign n4976 = /* LUT   23  2  3 */ n3044;
assign n4977 = /* LUT   16  3  3 */ !n2178;
assign n4978 = /* LUT   20 14  4 */ n2660;
assign n4982 = /* LUT    9 13  2 */ (n1146 ? n984 : (n1046 ? 1'b0 : n984));
assign n4983 = /* LUT   17  2  6 */ (n2312 ? 1'b1 : n2306);
assign n4984 = /* LUT   22 23  1 */ (n2297 ? 1'b0 : (n2986 ? (n2293 ? n2156 : 1'b0) : 1'b0));
assign n4987 = /* LUT    7  5  5 */ (n679 ? (n373 ? n362 : !n362) : (n373 ? (n362 ? 1'b1 : n963) : (n362 ? 1'b0 : n963)));
assign n4988 = /* LUT    8  1  3 */ (n200 ? (n828 ? (n1081 ? 1'b1 : n1083) : 1'b0) : n828);
assign n4991 = /* LUT   20 15  5 */ (n2156 ? 1'b0 : (n2293 ? 1'b0 : (n2432 ? !n2297 : 1'b0)));
assign n4994 = /* LUT   10 10  0 */ (n1464 ? 1'b0 : !n984);
assign n4995 = /* LUT   18 20  3 */ n2012;
assign n4996 = /* LUT   12 21  2 */ (n1839 ? !n1834 : n1834);
assign n4997 = /* LUT   17  3  7 */ (n2305 ? (n2333 ? io_19_0_1 : 1'b0) : 1'b0);
assign n4998 = /* LUT    3 14  5 */ (n76 ? (n106 ? n249 : (n249 ? n80 : 1'b0)) : (n106 ? n249 : 1'b0));
assign n4999 = /* LUT   10 13  5 */ (n904 ? n1320 : (n984 ? n1320 : 1'b0));
assign n5000 = /* LUT    9  9  4 */ (n573 ? n711 : 1'b0);
assign n5001 = /* LUT    2 15  1 */ (n257 ? 1'b0 : (n159 ? 1'b0 : !n5));
assign n5002 = /* LUT   18 13  0 */ n2656;
assign n5003 = /* LUT    1  3  2 */ (n10 ? (n34 ? (n186 ? n191 : !n191) : 1'b0) : (n34 ? 1'b0 : (n186 ? n191 : !n191)));
assign n5004 = /* LUT   13 12  7 */ n45;
assign n5005 = /* LUT    2 18  6 */ (n314 ? 1'b0 : (n139 ? (n318 ? 1'b1 : !n142) : 1'b1));
assign n5006 = /* LUT   13  4  3 */ (n1685 ? (n1877 ? 1'b1 : !n1249) : (n1877 ? n1249 : 1'b0));
assign n5007 = /* LUT   11 17  5 */ n188;
assign n5008 = /* LUT   18 16  5 */ n2415;
assign n5009 = /* LUT   12 13  3 */ (n1783 ? (n1771 ? 1'b1 : n1349) : (n1349 ? 1'b1 : n1782));
assign n5010 = /* LUT    4 19  0 */ (n781 ? (n8 ? n477 : !n477) : (n8 ? !n477 : n477));
assign n5011 = /* LUT    9  1  5 */ n188;
assign n5012 = /* LUT    2 19  7 */ (n320 ? (n319 ? n323 : 1'b0) : 1'b0);
assign n5013 = /* LUT   14 22  0 */ !n2008;
assign n5014 = /* LUT   22 11  4 */ (n2954 ? (n2950 ? !n2952 : n2952) : 1'b0);
assign n5015 = /* LUT    2 11  3 */ (n242 ? (n90 ? 1'b0 : (n73 ? 1'b1 : !n70)) : (n90 ? n73 : (n73 ? 1'b1 : !n70)));
assign n5016 = /* LUT    3 15  5 */ (n442 ? n287 : (n287 ? n598 : 1'b0));
assign n5017 = /* LUT    3  7  1 */ (n93 ? !n363 : 1'b0);
assign n5018 = /* LUT   11 18  6 */ n151;
assign n5021 = /* LUT   11 10  2 */ (n1412 ? !n852 : 1'b0);
assign n5022 = /* LUT   12  6  0 */ (n1559 ? (n1697 ? (n841 ? !n1291 : 1'b0) : (n841 ? !n1291 : 1'b1)) : (n841 ? !n1291 : 1'b0));
assign n5023 = /* LUT   24 20  2 */ n2012;
assign n5024 = /* LUT    4 20  1 */ (n639 ? 1'b1 : (n638 ? (n636 ? n785 : 1'b0) : n785));
assign n5025 = /* LUT   18  8  6 */ n1757;
assign n5026 = /* LUT   12  9  5 */ (n1728 ? (n1135 ? 1'b0 : !n1429) : (n1135 ? !n1429 : 1'b0));
assign n5027 = /* LUT    2 12  4 */ (n272 ? (n142 ? 1'b0 : !n117) : 1'b0);
assign n5028 = /* LUT   13  5  3 */ (n1684 ? (n1886 ? (n1249 ? !n1714 : 1'b1) : 1'b0) : 1'b0);
assign n5029 = /* LUT   22  4  1 */ (n2771 ? (n2772 ? (n2770 ? n2769 : 1'b0) : 1'b0) : 1'b0);
assign n5030 = /* LUT    2  4  0 */ n195;
assign n5031 = /* LUT   21  8  4 */ (n2949 ? (n2940 ? (n2801 ? n2689 : !n2689) : !n2801) : (n2940 ? (n2801 ? n2689 : !n2689) : n2801));
assign n5032 = /* LUT   14 18  2 */ (n2142 ? 1'b0 : (n1997 ? 1'b0 : n1996));
assign n5036 = /* LUT   18  1  3 */ (n2597 ? (n8 ? n2448 : !n2448) : (n8 ? !n2448 : n2448));
assign n5037 = /* LUT    8 18  5 */ (n477 ? (n1052 ? (n1055 ? 1'b0 : !n1207) : 1'b0) : (n1052 ? !n1207 : 1'b0));
assign n5038 = /* LUT   17 17  4 */ (n2409 ? (n2553 ? 1'b1 : n2011) : (n2553 ? !n2011 : 1'b0));
assign n5039 = /* LUT    7 19  1 */ n1059;
assign n5042 = /* LUT    5 11  4 */ (n815 ? (n583 ? 1'b0 : n764) : (n583 ? n764 : 1'b0));
assign n5043 = /* LUT    4 15  7 */ !n271;
assign n5047 = /* LUT   23 17  0 */ n2012;
assign n5048 = /* LUT    4  7  3 */ (n41 ? 1'b1 : (n400 ? (n44 ? 1'b0 : n6) : (n44 ? !n6 : 1'b1)));
assign n5051 = /* LUT   14 10  3 */ n1740;
assign n5052 = /* LUT    8 11  2 */ (n362 ? 1'b0 : (n679 ? n777 : 1'b1));
assign n5055 = /* LUT   15  9  6 */ (n2079 ? (n2075 ? (n2211 ? !n2082 : 1'b0) : 1'b0) : 1'b0);
assign n5056 = /* LUT    5 12  5 */ (n113 ? (n735 ? (n271 ? n579 : 1'b0) : 1'b0) : 1'b0);
assign n5057 = /* LUT    5  4  1 */ (n6 ? 1'b1 : (n541 ? (n213 ? 1'b0 : !n41) : (n213 ? n41 : 1'b1)));
assign n5058 = /* LUT    4  8  4 */ (n559 ? (n711 ? 1'b0 : n396) : !n711);
assign n5059 = /* LUT   16 22  6 */ n2012;
assign n5060 = /* LUT   16 14  2 */ n2250;
assign n5061 = /* LUT   17 18  4 */ (n2571 ? !n2412 : n2412);
assign n5065 = /* LUT   14  6  5 */ (n1895 ? 1'b0 : (n1894 ? 1'b0 : (n1897 ? 1'b0 : !n1898)));
assign n5066 = /* LUT    8  3  3 */ n189;
assign n5067 = /* LUT    1 21  5 */ (n156 ? 1'b0 : (n154 ? (n152 ? !n153 : 1'b0) : 1'b0));
assign n5068 = /* LUT   15  2  3 */ (n2053 ? (n1543 ? (n1890 ? 1'b0 : !n1863) : !n1863) : (n1543 ? !n1890 : 1'b1));
assign n5069 = /* LUT    1 13  1 */ (n96 ? (n94 ? 1'b0 : n99) : (n94 ? n99 : 1'b0));
assign n5070 = /* LUT   20 17  5 */ (n2727 ? (n2406 ? (n2856 ? n2403 : 1'b0) : 1'b0) : (n2406 ? (n2856 ? 1'b1 : !n2403) : 1'b0));
assign n5074 = /* LUT   23 13  7 */ (n3052 ? 1'b0 : n2841);
assign n5075 = /* LUT   16  6  3 */ n188;
assign n5076 = /* LUT   17  5  6 */ n2172;
assign n5077 = /* LUT   20 13  7 */ (n2702 ? (n2500 ? 1'b0 : (n2817 ? n2531 : 1'b0)) : 1'b1);
assign n5080 = /* LUT    7  8  5 */ (n994 ? (n869 ? 1'b0 : n981) : (n869 ? n981 : 1'b0));
assign n5081 = /* LUT   13 23  6 */ (n2043 ? (n2036 ? n1842 : !n1842) : n2036);
assign n5082 = /* LUT   20 10  1 */ (n2341 ? (n2345 ? n2375 : 1'b0) : 1'b0);
assign n5083 = /* LUT    3 18  1 */ (n309 ? !n312 : n312);
assign n5084 = /* LUT   17  6  7 */ n2476;
assign n5085 = /* LUT   16  2  5 */ n354;
assign n5086 = /* LUT    7  1  2 */ (n6 ? (n41 ? !n935 : 1'b1) : (n937 ? !n41 : 1'b1));
assign n5087 = /* LUT    9 12  4 */ n733;
assign n5088 = /* LUT    7  4  7 */ (n962 ? (n827 ? (n679 ? 1'b1 : !n806) : !n679) : (n827 ? n679 : (n679 ? 1'b0 : n806)));
assign n5089 = /* LUT    4 22  1 */ (n804 ? !n490 : n490);
assign n5090 = /* LUT   16  3  6 */ n189;
assign n5091 = /* LUT   11 21  1 */ (n1391 ? (n1511 ? n1522 : (n1521 ? 1'b1 : n1522)) : (n1511 ? 1'b0 : n1521));
assign n5092 = /* LUT   13 15  7 */ n1964;
assign n5093 = /* LUT   13  7  3 */ (n1896 ? 1'b0 : (n1916 ? 1'b0 : (n1908 ? 1'b0 : !n1568)));
assign n5094 = /* LUT   20  6  3 */ (n2786 ? !n2679 : n2679);
assign n5095 = /* LUT   18 11  1 */ (n2500 ? (n2509 ? 1'b0 : n2519) : (n2512 ? 1'b1 : n2509));
assign n5099 = /* LUT   10  8  6 */ n984;
assign n5100 = /* LUT    9  4  5 */ (n6 ? (n41 ? 1'b1 : !n1104) : (n41 ? !n1105 : 1'b1));
assign n5101 = /* LUT   22 14  4 */ n3028;
assign n5102 = /* LUT    2 14  3 */ (n277 ? (n267 ? !n281 : 1'b1) : (n267 ? (n281 ? 1'b0 : !n437) : !n437));
assign n5103 = /* LUT   13  8  4 */ (n1301 ? 1'b0 : (n1579 ? !n1740 : n1740));
assign n5104 = /* LUT   10  1  3 */ n179;
assign n5105 = /* LUT   11 16  7 */ (n1478 ? !n1459 : 1'b0);
assign n5106 = /* LUT   12 12  5 */ n1349;
assign n5107 = /* LUT   18  3  2 */ (n852 ? (n2455 ? (n2340 ? n2066 : 1'b1) : (n2340 ? 1'b0 : !n2066)) : (n2455 ? (n2340 ? 1'b1 : n2066) : (n2340 ? !n2066 : 1'b0)));
assign n5108 = /* LUT   22 15  5 */ (n2976 ? 1'b0 : (n3022 ? 1'b0 : (n2966 ? 1'b0 : !n3024)));
assign n5109 = /* LUT    2 15  4 */ (n282 ? (n258 ? (n288 ? !n257 : 1'b0) : !n257) : 1'b0);
assign n5110 = /* LUT   12  4  1 */ (n1126 ? 1'b0 : (n973 ? (n852 ? n1125 : 1'b0) : 1'b0));
assign n5111 = /* LUT   22  7  1 */ (n2938 ? n2940 : 1'b1);
assign n5112 = /* LUT    2  7  0 */ (n391 ? (n225 ? 1'b1 : !n222) : (n397 ? 1'b1 : (n225 ? 1'b1 : !n222)));
assign n5113 = /* LUT   21 11  4 */ n1965;
assign n5114 = /* LUT   24 18  3 */ n2012;
assign n5118 = /* LUT   15 17  0 */ (n1822 ? 1'b0 : !n5);
assign n5119 = /* LUT   13  4  6 */ (n1880 ? (n1422 ? n1435 : !n1881) : (n1422 ? n1435 : 1'b1));
assign n5120 = /* LUT   17 21  0 */ (n2022 ? 1'b0 : (n2292 ? 1'b0 : (n2427 ? 1'b0 : !n2426)));
assign n5121 = /* LUT   11  9  4 */ (n984 ? (n1135 ? n1146 : (n1146 ? 1'b1 : n5)) : 1'b0);
assign n5122 = /* LUT    8 21  5 */ (n1067 ? n929 : (n929 ? 1'b1 : (n1074 ? 1'b0 : n1064)));
assign n5123 = /* LUT   12  5  2 */ (n1545 ? (n1548 ? n841 : 1'b0) : (n1548 ? (n841 ? 1'b1 : !n1551) : (n841 ? 1'b0 : !n1551)));
assign n5124 = /* LUT   17 20  4 */ (n5 ? 1'b1 : !n2022);
assign n5125 = /* LUT   15 12  7 */ (n2238 ? (n2122 ? 1'b0 : !n2094) : (n2122 ? 1'b0 : !n1740));
assign n5128 = /* LUT   21  7  6 */ n2943;
assign n5129 = /* LUT    4 10  3 */ n189;
assign n5130 = /* LUT   14 13  3 */ (n1936 ? (n1770 ? 1'b0 : !n2102) : !n1770);
assign n5131 = /* LUT    8 14  2 */ n45;
assign n5132 = /* LUT    2  2  6 */ n354;
assign n5135 = /* LUT    5 15  5 */ (n597 ? 1'b0 : n603);
assign n5136 = /* LUT    5  7  1 */ n354;
assign n5137 = /* LUT   17 16  6 */ n1480;
assign n5138 = /* LUT    4 11  4 */ (n88 ? (n736 ? (n729 ? !n737 : 1'b0) : n729) : (n736 ? !n737 : 1'b1));
assign n5139 = /* LUT    4  3  0 */ (n176 ? 1'b0 : (n667 ? n660 : 1'b0));
assign n5142 = /* LUT    2  3  7 */ n184;
assign n5146 = /* LUT   14  9  5 */ n1755;
assign n5147 = /* LUT   15  5  3 */ n354;
assign n5148 = /* LUT    5  8  2 */ (n811 ? (n711 ? (n5 ? !n60 : 1'b0) : 1'b1) : 1'b0);
assign n5149 = /* LUT   17 17  7 */ (n2011 ? n2413 : n2551);
assign n5150 = /* LUT    7 19  4 */ !n490;
assign n5151 = /* LUT    4  4  1 */ (n678 ? (n6 ? 1'b1 : (n41 ? 1'b0 : !n680)) : (n6 ? 1'b1 : (n41 ? 1'b1 : !n680)));
assign n5152 = /* LUT    7 11  0 */ (n698 ? 1'b0 : (n1020 ? !n362 : 1'b1));
assign n5153 = /* LUT    5 11  7 */ (n764 ? !n733 : 1'b0);
assign n5156 = /* LUT    4  7  6 */ (n402 ? (n545 ? n372 : (n694 ? 1'b0 : n372)) : (n694 ? 1'b0 : n372));
assign n5157 = /* LUT   13 22  0 */ (n1842 ? (n1846 ? (n2030 ? n1835 : 1'b1) : (n2030 ? 1'b0 : !n1835)) : (n1846 ? (n2030 ? 1'b1 : n1835) : (n2030 ? !n1835 : 1'b0)));
assign n5158 = /* LUT   14 10  6 */ n1933;
assign n5159 = /* LUT   14  2  2 */ (n852 ? n1001 : 1'b0);
assign n5160 = /* LUT    1 17  2 */ (n308 ? (n122 ? 1'b0 : n307) : (n122 ? n307 : 1'b0));
assign n5161 = /* LUT   17  9  2 */ (n2366 ? (n2498 ? 1'b0 : !n2494) : n2349);
assign n5162 = /* LUT    8  2  5 */ (n41 ? (n953 ? !n6 : 1'b1) : (n6 ? 1'b1 : !n944));
assign n5163 = /* LUT    1 20  7 */ (n329 ? 1'b1 : (n150 ? (n137 ? !n149 : 1'b1) : 1'b1));
assign n5164 = /* LUT    7  3  1 */ (n959 ? (n841 ? (n5 ? 1'b1 : n954) : 1'b1) : (n841 ? (n5 ? 1'b1 : n954) : 1'b0));
assign n5165 = /* LUT   10 11  2 */ n1471;
assign n5166 = /* LUT    9 15  5 */ (n1146 ? n984 : (n1359 ? n984 : 1'b0));
assign n5167 = /* LUT   13 18  2 */ (n1812 ? (n1982 ? (n1808 ? n5 : 1'b1) : (n1808 ? 1'b0 : !n5)) : (n1982 ? (n1808 ? 1'b1 : n5) : (n1808 ? !n5 : 1'b0)));
assign n5168 = /* LUT    3 21  1 */ (n45 ? n482 : 1'b0);
assign n5169 = /* LUT    8  3  6 */ n179;
assign n5170 = /* LUT    1 13  4 */ (n87 ? 1'b0 : (n278 ? !n62 : (n62 ? 1'b0 : !n266)));
assign n5171 = /* LUT   17  1  3 */ (n2442 ? (n2314 ? !n2439 : 1'b0) : 1'b0);
assign n5172 = /* LUT   20  9  4 */ n1754;
assign n5173 = /* LUT   18 14  2 */ n2659;
assign n5174 = /* LUT    9  7  0 */ (n208 ? 1'b0 : !n811);
assign n5175 = /* LUT    7  7  7 */ !n869;
assign n5176 = /* LUT   21 21  2 */ (n2875 ? n2408 : (n2408 ? (n2431 ? 1'b1 : !n2404) : 1'b0));
assign n5177 = /* LUT   16  6  6 */ (n1890 ? 1'b0 : (n1463 ? !n1731 : n1731));
assign n5180 = /* LUT   10 12  2 */ (n1330 ? 1'b0 : n1473);
assign n5181 = /* LUT    1  5  5 */ n37;
assign n5182 = /* LUT   15 19  0 */ n2284;
assign n5183 = /* LUT    3 16  7 */ (n80 ? (n612 ? (n605 ? n111 : 1'b0) : 1'b0) : 1'b0);
assign n5184 = /* LUT   21 22  3 */ n2012;
assign n5185 = /* LUT   22 18  0 */ (n2855 ? (n2293 ? 1'b0 : (n2156 ? 1'b0 : n2297)) : 1'b0);
assign n5186 = /* LUT   12 15  6 */ (n1493 ? (n1181 ? 1'b0 : (n1489 ? n1613 : 1'b0)) : (n1181 ? 1'b0 : n1613));
assign n5187 = /* LUT   12  7  2 */ (n1427 ? 1'b0 : (n1576 ? !n1454 : n1454));
assign n5188 = /* LUT   13  3  0 */ (n1543 ? (n1863 ? (n1691 ? 1'b0 : !n1689) : !n1689) : (n1863 ? !n1691 : 1'b1));
assign n5189 = /* LUT    4 21  3 */ n799;
assign n5190 = /* LUT   18 15  2 */ n2012;
assign n5191 = /* LUT   22 13  7 */ (n3017 ? (n3016 ? 1'b0 : (n2825 ? 1'b0 : !n2818)) : (n3016 ? (n2825 ? !n2818 : 1'b0) : !n2818));
assign n5192 = /* LUT    3  9  4 */ n572;
assign n5193 = /* LUT   11 19  7 */ (n1511 ? (n1380 ? !n1520 : 1'b0) : (n1514 ? 1'b1 : (n1380 ? !n1520 : 1'b0)));
assign n5194 = /* LUT    2 10  0 */ (n106 ? n65 : (n65 ? 1'b1 : n244));
assign n5195 = /* LUT    5 18  1 */ (n648 ? (n785 ? !n642 : 1'b0) : (n627 ? n785 : (n785 ? !n642 : 1'b0)));
assign n5196 = /* LUT    9  3  7 */ (n1107 ? (n1095 ? (n1244 ? !n841 : 1'b0) : !n841) : (n1244 ? !n841 : 1'b0));
assign n5197 = /* LUT   21  6  0 */ n2608;
assign n5198 = /* LUT   18  2  5 */ n2310;
assign n5199 = /* LUT   13  7  6 */ (n1037 ? (n1912 ? !n1722 : 1'b1) : (n1722 ? n1915 : 1'b0));
assign n5200 = /* LUT    3  2  1 */ n233;
assign n5201 = /* LUT   11 12  4 */ (n212 ? 1'b0 : n1457);
assign n5202 = /* LUT   12  8  2 */ n189;
assign n5203 = /* LUT   11  4  0 */ (n1415 ? 1'b0 : n1106);
assign n5204 = /* LUT   15 16  3 */ !n1790;
assign n5205 = /* LUT    3  1  5 */ n15;
assign n5206 = /* LUT   22 14  7 */ n3030;
assign n5207 = /* LUT   15 15  7 */ (n1645 ? (n1517 ? !n1608 : 1'b1) : 1'b1);
assign n5208 = /* LUT    5 10  2 */ (n811 ? (n711 ? (n566 ? 1'b0 : n5) : 1'b1) : 1'b0);
assign n5209 = /* LUT    7 21  4 */ (n927 ? (n1060 ? 1'b0 : n151) : (n1060 ? 1'b0 : (n277 ? n151 : 1'b1)));
assign n5210 = /* LUT   11  5  1 */ (n1125 ? 1'b0 : (n1416 ? (n1126 ? 1'b0 : !n1541) : 1'b0));
assign n5213 = /* LUT    5 13  7 */ (n271 ? (n128 ? (n747 ? !n113 : 1'b0) : 1'b0) : 1'b0);
assign n5214 = /* LUT   23 19  3 */ n2012;
assign n5215 = /* LUT    4  9  6 */ (n221 ? !n711 : (n559 ? 1'b0 : !n711));
assign n5216 = /* LUT   15  8  4 */ n2204;
assign n5217 = /* LUT   17 19  6 */ n2579;
assign n5218 = /* LUT   17 11  2 */ (n2520 ? (n2341 ? 1'b0 : n577) : (n2341 ? n577 : 1'b0));
assign n5219 = /* LUT    4  6  0 */ (n693 ? (n41 ? !n6 : (n6 ? 1'b1 : !n692)) : (n41 ? 1'b1 : (n6 ? 1'b1 : !n692)));
assign n5220 = /* LUT    7 14  1 */ (n4 ? (n564 ? (n816 ? 1'b0 : !n906) : !n906) : !n906);
assign n5221 = /* LUT    2  6  7 */ (n200 ? 1'b1 : (n207 ? (n176 ? !n388 : 1'b1) : (n176 ? !n388 : 1'b0)));
assign n5222 = /* LUT   16 20  2 */ (n2297 ? 1'b0 : (n2156 ? 1'b0 : (n2293 ? 1'b0 : n2428)));
assign n5223 = /* LUT   14 12  5 */ (n1740 ? (n2104 ? !n2102 : (n2102 ? 1'b0 : n2100)) : (n2102 ? 1'b0 : n2100));
assign n5224 = /* LUT   14  4  1 */ n233;
assign n5225 = /* LUT   17 20  7 */ (n2293 ? (n2422 ? (n2412 ? n2022 : 1'b0) : (n2412 ? 1'b1 : !n2022)) : (n2422 ? (n2412 ? 1'b1 : !n2022) : (n2412 ? n2022 : 1'b0)));
assign n5226 = /* LUT   17 12  3 */ n2389;
assign n5227 = /* LUT   23  3  0 */ n3047;
assign n5228 = /* LUT   15  4  6 */ (n1249 ? (n2052 ? !n2179 : 1'b0) : n2052);
assign n5229 = /* LUT    5  6  3 */ (n699 ? (n5 ? 1'b1 : (n698 ? n365 : 1'b1)) : (n5 ? n698 : (n698 ? n365 : 1'b0)));
assign n5230 = /* LUT   14 13  6 */ (n1772 ? n1761 : (n1494 ? n1761 : n1948));
assign n5231 = /* LUT    4  2  2 */ (n510 ? 1'b0 : !n513);
assign n5232 = /* LUT   14  5  2 */ (n1541 ? (n1126 ? 1'b0 : (n1416 ? !n1125 : 1'b0)) : 1'b0);
assign n5233 = /* LUT   16 16  4 */ (n2274 ? 1'b0 : (n2277 ? n2272 : 1'b0));
assign n5234 = /* LUT   13 21  3 */ (n1491 ? (n5 ? 1'b0 : !n1833) : (n5 ? 1'b0 : (n2021 ? 1'b0 : !n1833)));
assign n5235 = /* LUT    8  5  5 */ (n976 ? (n958 ? (n807 ? 1'b1 : n980) : n807) : (n958 ? n980 : 1'b0));
assign n5236 = /* LUT   24  3  4 */ !n2901;
assign n5237 = /* LUT   10 14  2 */ (n1356 ? (n1341 ? (n1344 ? !n1183 : 1'b1) : 1'b0) : (n1341 ? !n1344 : 1'b0));
assign n5240 = /* LUT    9 10  1 */ (n362 ? (n698 ? 1'b0 : !n1021) : !n698);
assign n5241 = /* LUT   16  9  1 */ (n2355 ? (n2364 ? !n2199 : !n2207) : n2364);
assign n5242 = /* LUT    7  2  4 */ (n200 ? (n948 ? 1'b0 : !n942) : 1'b0);
assign n5243 = /* LUT    8  6  6 */ (n891 ? !n852 : 1'b0);
assign n5244 = /* LUT   16  8  5 */ (n2206 ? 1'b0 : (n2198 ? (n2205 ? !n2208 : 1'b0) : 1'b0));
assign n5245 = /* LUT   10 15  3 */ (n1356 ? (n1352 ? (n1361 ? !n1191 : 1'b1) : 1'b0) : (n1352 ? !n1361 : 1'b0));
assign n5246 = /* LUT   20  4  0 */ !n2481;
assign n5247 = /* LUT   18 17  2 */ (n2589 ? (n2557 ? 1'b0 : n2404) : (n2557 ? !n2404 : 1'b1));
assign n5248 = /* LUT   13 22  3 */ (n1491 ? (n2025 ? (n1835 ? 1'b0 : !n5) : 1'b0) : (n1835 ? 1'b0 : !n5));
assign n5252 = /* LUT    9 14  7 */ n189;
assign n5255 = /* LUT   16  4  7 */ (n2303 ? (io_19_0_1 ? n2182 : 1'b0) : 1'b0);
assign n5256 = /* LUT    1  8  5 */ (n56 ? (n58 ? 1'b1 : !n65) : n58);
assign n5257 = /* LUT    9 11  1 */ (n711 ? (n60 ? n811 : 1'b0) : n811);
assign n5258 = /* LUT    7  3  4 */ (n371 ? (n51 ? 1'b1 : (n833 ? 1'b0 : !n830)) : (n51 ? (n833 ? 1'b0 : !n830) : 1'b0));
assign n5259 = /* LUT   12 18  6 */ (n1642 ? 1'b0 : n1640);
assign n5260 = /* LUT    2 13  1 */ (n96 ? (n94 ? (n95 ? n80 : 1'b0) : 1'b0) : 1'b0);
assign n5261 = /* LUT   13  6  0 */ (n1554 ? 1'b0 : (n1418 ? !n1705 : n1705));
assign n5262 = /* LUT    2 16  6 */ (n258 ? n112 : 1'b0);
assign n5263 = /* LUT   13  9  5 */ (n1751 ? (n1729 ? (n1291 ? 1'b1 : n1281) : 1'b0) : (n1729 ? (n1291 ? n1281 : 1'b1) : 1'b0));
assign n5264 = /* LUT    3 12  4 */ (n5 ? 1'b0 : (n584 ? !n277 : (n138 ? !n277 : 1'b0)));
assign n5265 = /* LUT    1  4  7 */ n36;
assign n5266 = /* LUT   15 18  2 */ n2281;
assign n5267 = /* LUT    4 17  0 */ (n111 ? (n448 ? (n612 ? 1'b0 : n454) : 1'b0) : 1'b0);
assign n5268 = /* LUT    2 17  7 */ (n363 ? 1'b0 : (io_4_31_0 ? n114 : !n114));
assign n5269 = /* LUT   13 10  6 */ n1593;
assign n5270 = /* LUT   13  2  2 */ n188;
assign n5271 = /* LUT    2  9  3 */ !n421;
assign n5274 = /* LUT    3  5  1 */ (n6 ? !n41 : 1'b0);
assign n5275 = /* LUT   11 15  4 */ (n258 ? (n1491 ? n1623 : 1'b0) : (n1491 ? n1623 : (n1500 ? n1623 : 1'b0)));
assign n5276 = /* LUT   14 23  5 */ (n2165 ? (n1847 ? n8 : !n8) : (n1847 ? !n8 : n8));
assign n5277 = /* LUT   11  7  0 */ (n841 ? n1577 : !n1574);
assign n5280 = /* LUT   10  3  5 */ n175;
assign n5281 = /* LUT   18  6  6 */ (n2615 ? !n2470 : n2470);
assign n5282 = /* LUT   12  7  5 */ (n1427 ? 1'b0 : (n1732 ? !n1576 : n1576));
assign n5283 = /* LUT   22  9  3 */ n2616;
assign n5284 = /* LUT   21 13  6 */ (n2824 ? !n2818 : n2818);
assign n5285 = /* LUT    4 21  6 */ (n801 ? !n477 : n477);
assign n5286 = /* LUT   21  5  2 */ (n2931 ? (n8 ? !n2926 : n2926) : (n8 ? n2926 : !n2926));
assign n5287 = /* LUT    8 16  5 */ !n1019;
assign n5288 = /* LUT   15  3  0 */ n179;
assign n5289 = /* LUT   17 22  6 */ (n2297 ? (n2156 ? 1'b0 : (n2432 ? n2293 : 1'b0)) : 1'b0);
assign n5290 = /* LUT   22  2  0 */ (n2324 ? 1'b0 : (io_19_0_1 ? 1'b1 : !n2757));
assign n5291 = /* LUT    7 17  1 */ (n448 ? (n465 ? (n302 ? n5 : 1'b1) : 1'b1) : 1'b1);
assign n5292 = /* LUT   15  6  5 */ (n2196 ? (n1541 ? (n2066 ? n2192 : 1'b0) : (n2066 ? n2192 : 1'b1)) : (n1541 ? (n2066 ? n2192 : 1'b1) : (n2066 ? n2192 : 1'b0)));
assign n5293 = /* LUT    5  9  4 */ (n717 ? (n810 ? (n560 ? 1'b0 : n725) : n725) : (n560 ? 1'b0 : n725));
assign n5294 = /* LUT    4 13  7 */ (n440 ? (n121 ? (n592 ? !n445 : 1'b0) : 1'b0) : 1'b0);
assign n5295 = /* LUT    4  5  3 */ (n522 ? (n6 ? 1'b0 : !n365) : (n6 ? 1'b1 : !n390));
assign n5296 = /* LUT   16 19  5 */ (n2156 ? 1'b0 : (n2293 ? 1'b0 : (n2297 ? 1'b0 : n2298)));
assign n5297 = /* LUT   17 15  3 */ (n2397 ? n2395 : (n2270 ? (n2395 ? !n2272 : 1'b0) : 1'b0));
assign n5298 = /* LUT   11  3  7 */ n354;
assign n5301 = /* LUT   15  7  6 */ (n1692 ? (n1593 ? 1'b0 : !n1904) : (n1593 ? !n1904 : 1'b0));
assign n5302 = /* LUT    9 21  0 */ (n1388 ? (n932 ? n8 : !n8) : (n932 ? !n8 : n8));
assign n5303 = /* LUT    7 21  7 */ (n1031 ? n15 : 1'b0);
assign n5304 = /* LUT   14  8  2 */ (n1752 ? (n1888 ? 1'b0 : !n2049) : (n1888 ? !n2049 : 1'b0));
assign n5305 = /* LUT    8  9  1 */ (n812 ? !n880 : n880);
assign n5306 = /* LUT   20 23  3 */ (n2297 ? 1'b0 : (n2293 ? (n2156 ? n2432 : 1'b0) : 1'b0));
assign n5307 = /* LUT   17  8  0 */ n2204;
assign n5308 = /* LUT    5  2  0 */ (n355 ? (n41 ? !n6 : (n6 ? 1'b1 : !n666)) : (n41 ? 1'b1 : (n6 ? 1'b1 : !n666)));
assign n5309 = /* LUT   23  2  2 */ (n3043 ? (n8 ? n3005 : !n3005) : (n8 ? !n3005 : n3005));
assign n5310 = /* LUT    4  6  3 */ (n372 ? (n402 ? (n213 ? 1'b1 : n385) : n385) : 1'b0);
assign n5311 = /* LUT   17 11  5 */ n2345;
assign n5312 = /* LUT    9 13  1 */ (n1044 ? (n806 ? 1'b0 : !n679) : !n679);
assign n5313 = /* LUT   16 12  1 */ n1754;
assign n5317 = /* LUT    7  5  4 */ (n684 ? (n698 ? 1'b1 : n844) : (n5 ? (n698 ? 1'b1 : n844) : (n698 ? 1'b0 : n844)));
assign n5318 = /* LUT   14  4  4 */ (n1871 ? (n1875 ? 1'b0 : (n1874 ? !n1647 : 1'b1)) : (n1874 ? !n1647 : 1'b1));
assign n5319 = /* LUT    8  1  2 */ n188;
assign n5320 = /* LUT    1 19  4 */ (n135 ? (n151 ? 1'b0 : !n136) : !n151);
assign n5323 = /* LUT    1 11  0 */ (n70 ? !n75 : 1'b0);
assign n5324 = /* LUT    8  4  7 */ (n51 ? 1'b0 : n52);
assign n5328 = /* LUT   12 21  1 */ (n1833 ? !n1831 : n1831);
assign n5329 = /* LUT   17  3  6 */ (io_19_0_1 ? (n2304 ? n2182 : 1'b0) : 1'b0);
assign n5330 = /* LUT    7  6  5 */ (n861 ? (n967 ? !n852 : 1'b0) : 1'b0);
assign n5331 = /* LUT   10 13  4 */ (n1459 ? 1'b0 : !n5);
assign n5332 = /* LUT    9 17  7 */ !n907;
assign n5333 = /* LUT    9  9  3 */ n811;
assign n5334 = /* LUT   13 21  6 */ (n1656 ? (n2021 ? (n5 ? 1'b0 : n1491) : !n5) : 1'b0);
assign n5335 = /* LUT    1 12  1 */ (n69 ? (n244 ? !n84 : 1'b0) : 1'b0);
assign n5338 = /* LUT   12 22  2 */ (n1850 ? !n1843 : n1843);
assign n5339 = /* LUT   20 11  6 */ n2644;
assign n5340 = /* LUT   10 14  5 */ (n1351 ? (n1356 ? 1'b0 : n1345) : (n1356 ? (n1345 ? !n1283 : 1'b0) : n1345));
assign n5341 = /* LUT   10  6  1 */ (n1126 ? (n1125 ? n1424 : 1'b0) : 1'b0);
assign n5342 = /* LUT   18 16  4 */ n2412;
assign n5343 = /* LUT    9 10  4 */ (n1008 ? (n1306 ? 1'b0 : (n1154 ? n727 : 1'b0)) : n727);
assign n5344 = /* LUT    9  2  0 */ (n1080 ? (n1245 ? n1251 : 1'b1) : (n1245 ? (n1107 ? 1'b0 : n1251) : !n1107));
assign n5345 = /* LUT   22 20  3 */ (n2293 ? (n2156 ? 1'b0 : (n2848 ? !n2297 : 1'b0)) : 1'b0);
assign n5346 = /* LUT    7  2  7 */ n188;
assign n5347 = /* LUT   21 24  6 */ n2012;
assign n5348 = /* LUT    2 19  6 */ (n323 ? 1'b0 : n307);
assign n5349 = /* LUT   13 13  7 */ n1949;
assign n5350 = /* LUT    3 15  4 */ (n446 ? n80 : 1'b0);
assign n5351 = /* LUT   20  4  3 */ !n2775;
assign n5352 = /* LUT    3  7  0 */ n179;
assign n5353 = /* LUT   11 18  5 */ (n1490 ? !n264 : 1'b0);
assign n5354 = /* LUT   18  9  1 */ (n2355 ? (n2364 ? 1'b0 : n2371) : (n2489 ? !n2364 : 1'b0));
assign n5355 = /* LUT    4 20  0 */ (n626 ? n785 : (n785 ? !n480 : 1'b0));
assign n5356 = /* LUT    2 20  7 */ (n148 ? (n151 ? (n146 ? n149 : 1'b1) : 1'b0) : n151);
assign n5357 = /* LUT   12  9  4 */ (n1281 ? !n1588 : (n1291 ? (n1749 ? !n1588 : 1'b0) : (n1749 ? 1'b0 : !n1588)));
assign n5358 = /* LUT   22 12  4 */ (n2809 ? 1'b0 : (n2509 ? 1'b0 : n2500));
assign n5359 = /* LUT    2 12  3 */ (n151 ? (n257 ? 1'b0 : n256) : (n249 ? (n257 ? 1'b0 : n256) : 1'b0));
assign n5360 = /* LUT   13  5  2 */ (n1682 ? (n1887 ? 1'b1 : (n1410 ? !n1693 : 1'b1)) : (n1887 ? (n1410 ? 1'b1 : !n1693) : !n1693));
assign n5361 = /* LUT    3  8  1 */ (n66 ? !n53 : n53);
assign n5364 = /* LUT   14 18  1 */ (n1993 ? (n2140 ? (n1823 ? 1'b1 : !n2000) : (n1823 ? 1'b0 : !n2000)) : (n2140 ? (n1823 ? 1'b0 : n2000) : (n1823 ? 1'b1 : n2000)));
assign n5365 = /* LUT    3 11  6 */ (n271 ? 1'b0 : (n575 ? (n17 ? n113 : 1'b0) : 1'b0));
assign n5366 = /* LUT   11 14  7 */ (n1464 ? 1'b0 : (n1487 ? 1'b0 : (n1171 ? 1'b0 : !n904)));
assign n5367 = /* LUT   18  1  2 */ (n2596 ? (n2447 ? n8 : !n8) : (n2447 ? !n8 : n8));
assign n5368 = /* LUT    2 13  4 */ (n282 ? !n5 : 1'b0);
assign n5369 = /* LUT   13  6  3 */ (n1871 ? 1'b0 : (n1694 ? !n1753 : n1753));
assign n5370 = /* LUT    2  5  0 */ (n199 ? (n196 ? n383 : 1'b0) : 1'b0);
assign n5371 = /* LUT    4 16  2 */ (n91 ? !n612 : 1'b0);
assign n5374 = /* LUT   14 19  2 */ (n2148 ? (n2006 ? n1982 : !n1982) : (n2006 ? !n1982 : n1982));
assign n5375 = /* LUT   22  8  6 */ (n2946 ? (n1 ? 1'b0 : !n1645) : 1'b0);
assign n5379 = /* LUT    3  4  3 */ (n525 ? (n376 ? (n199 ? n205 : 1'b0) : n205) : (n199 ? n205 : 1'b0));
assign n5380 = /* LUT   21  4  5 */ (n2921 ? (n2773 ? n8 : !n8) : (n2773 ? !n8 : n8));
assign n5385 = /* LUT   22  5  0 */ (n2675 ? n2928 : (n2928 ? (n2673 ? 1'b1 : n2674) : 1'b0));
assign n5388 = /* LUT    4  8  3 */ (n559 ? (n711 ? 1'b0 : n44) : !n711);
assign n5389 = /* LUT    8 20  6 */ (n1044 ? (n8 ? (n1064 ? n1043 : 1'b0) : (n1064 ? !n1043 : 1'b0)) : (n8 ? (n1064 ? !n1043 : 1'b0) : (n1064 ? n1043 : 1'b0)));
assign n5390 = /* LUT   11  7  3 */ (n1575 ? (n1444 ? (n841 ? 1'b1 : !n1443) : 1'b1) : (n1444 ? (n841 ? 1'b0 : !n1443) : !n841));
assign n5391 = /* LUT   17 18  3 */ (n2570 ? !n2411 : n2411);
assign n5392 = /* LUT   15 10  6 */ n1755;
assign n5393 = /* LUT   15  2  2 */ n179;
assign n5394 = /* LUT    5  5  1 */ (n684 ? (n683 ? !n6 : (n41 ? !n6 : 1'b1)) : (n683 ? (n41 ? 1'b1 : !n6) : 1'b1));
assign n5395 = /* LUT    4  1  0 */ n354;
assign n5396 = /* LUT   16 15  2 */ n2131;
assign n5397 = /* LUT   15  3  3 */ (n1541 ? n1416 : 1'b0);
assign n5398 = /* LUT   23 13  6 */ (n2810 ? 1'b1 : n2711);
assign n5399 = /* LUT   17 14  5 */ (n2548 ? !n2267 : n2267);
assign n5400 = /* LUT    1 14  1 */ (n244 ? (n116 ? n76 : 1'b0) : 1'b0);
assign n5401 = /* LUT    7 17  4 */ (n133 ? (n448 ? (n5 ? 1'b0 : n302) : 1'b0) : 1'b0);
assign n5405 = /* LUT    2  1  6 */ (n166 ? (n162 ? n41 : (n6 ? 1'b1 : n41)) : (n162 ? (n6 ? n41 : 1'b1) : 1'b1));
assign n5409 = /* LUT   14  7  4 */ n189;
assign n5410 = /* LUT   13 23  5 */ (n2042 ? (n2035 ? n1842 : !n1842) : n2035);
assign n5416 = /* LUT   10 16  4 */ (n1201 ? !n1268 : 1'b0);
assign n5417 = /* LUT    7  1  1 */ (n41 ? (n836 ? !n6 : 1'b1) : (n6 ? !n835 : 1'b1));
assign n5418 = /* LUT    9 20  7 */ (n1387 ? (n8 ? n907 : !n907) : (n8 ? !n907 : n907));
assign n5419 = /* LUT    9 12  3 */ (n1141 ? n1331 : (n1331 ? !n1174 : 1'b0));
assign n5420 = /* LUT    7  4  6 */ (n5 ? (n831 ? 1'b1 : n362) : (n357 ? (n831 ? 1'b1 : n362) : (n831 ? !n362 : 1'b0)));
assign n5421 = /* LUT    3 19  1 */ (n621 ? !n620 : n620);
assign n5422 = /* LUT   20 14  6 */ n2653;
assign n5423 = /* LUT   10 17  5 */ n179;
assign n5424 = /* LUT   20  6  2 */ (n2785 ? !n2678 : n2678);
assign n5425 = /* LUT   10  9  1 */ (n1288 ? !n1289 : 1'b0);
assign n5426 = /* LUT    9 13  4 */ (n806 ? (n679 ? 1'b0 : !n1043) : !n679);
assign n5427 = /* LUT    9  5  0 */ (n1114 ? (n5 ? (n1266 ? 1'b0 : !n841) : (n1266 ? 1'b1 : n841)) : (n5 ? 1'b0 : !n841));
assign n5428 = /* LUT    7  5  7 */ (n958 ? (n976 ? (n960 ? 1'b1 : n975) : n975) : (n976 ? n960 : 1'b0));
assign n5431 = /* LUT   13  8  3 */ (n1741 ? (n1701 ? 1'b0 : !n1679) : (n1701 ? 1'b0 : n1679));
assign n5432 = /* LUT   18 12  1 */ (n2527 ? (n2509 ? !n2500 : (n2526 ? 1'b1 : !n2500)) : (n2509 ? !n2500 : (n2526 ? n2500 : 1'b0)));
assign n5433 = /* LUT    3 14  7 */ (n284 ? (n113 ? 1'b1 : n271) : 1'b0);
assign n5434 = /* LUT   10  1  2 */ n15;
assign n5435 = /* LUT   22 15  4 */ (n3037 ? (n8 ? n2974 : !n2974) : (n8 ? !n2974 : n2974));
assign n5436 = /* LUT    2 15  3 */ (n249 ? (n289 ? !n117 : 1'b0) : 1'b0);
assign n5437 = /* LUT   10  4  7 */ n177;
assign n5438 = /* LUT   21 11  3 */ n1789;
assign n5439 = /* LUT   14 21  1 */ (n2021 ? (n2020 ? 1'b0 : (n5 ? 1'b0 : n1491)) : (n2020 ? 1'b0 : !n5));
assign n5440 = /* LUT    1  3  4 */ n18;
assign n5441 = /* LUT   13  4  5 */ (n1676 ? (n1427 ? (n1422 ? 1'b1 : !n1681) : (n1422 ? 1'b0 : !n1681)) : (n1427 ? 1'b1 : !n1422));
assign n5442 = /* LUT   11 17  7 */ (n212 ? (n1359 ? n1510 : 1'b0) : (n1510 ? n1328 : 1'b0));
assign n5443 = /* LUT   11  9  3 */ (n1297 ? (n1438 ? (n718 ? 1'b0 : n1437) : n1437) : (n1438 ? 1'b0 : n1437));
assign n5444 = /* LUT   12 13  5 */ (n1783 ? (n1774 ? 1'b1 : n1349) : (n1627 ? 1'b1 : n1349));
assign n5445 = /* LUT   12  5  1 */ n175;
assign n5449 = /* LUT    4 19  2 */ n789;
assign n5450 = /* LUT    9  1  7 */ n177;
assign n5451 = /* LUT    2 11  5 */ (n264 ? (n272 ? !n304 : 1'b0) : (n272 ? !n117 : 1'b0));
assign n5454 = /* LUT   11 10  4 */ (n1425 ? n852 : 1'b1);
assign n5455 = /* LUT   15 21  5 */ n2134;
assign n5456 = /* LUT   12  6  2 */ (n1435 ? 1'b0 : (n1718 ? !n1548 : n1548));
assign n5457 = /* LUT   15 13  1 */ (n2117 ? (n2116 ? n1474 : 1'b0) : (n2237 ? (n2116 ? n1474 : 1'b0) : n2116));
assign n5458 = /* LUT    5 16  0 */ (n267 ? n760 : 1'b0);
assign n5459 = /* LUT   12  9  7 */ (n1270 ? 1'b0 : (n1463 ? !n1577 : n1577));
assign n5460 = /* LUT   22 12  7 */ (n2809 ? 1'b0 : (n2500 ? 1'b0 : !n2509));
assign n5461 = /* LUT   22  4  3 */ (n2675 ? 1'b1 : (n7 ? 1'b1 : (n2673 ? 1'b1 : n2674)));
assign n5462 = /* LUT    2  4  2 */ (n22 ? (n181 ? (n36 ? n194 : 1'b0) : (n36 ? !n194 : 1'b0)) : (n181 ? (n36 ? 1'b0 : n194) : (n36 ? 1'b0 : !n194)));
assign n5463 = /* LUT   21  8  6 */ (n2803 ? (n2940 ? n2688 : !n2800) : (n2940 ? !n2688 : n2800));
assign n5464 = /* LUT    4 11  3 */ (n128 ? n297 : 1'b0);
assign n5467 = /* LUT    2  3  6 */ n181;
assign n5468 = /* LUT    8 18  7 */ (n777 ? 1'b0 : (n642 ? 1'b0 : (n630 ? 1'b0 : !n621)));
assign n5469 = /* LUT   18  1  5 */ (n2599 ? (n2314 ? n2439 : 1'b0) : 1'b0);
assign n5470 = /* LUT   15  5  2 */ (n1691 ? 1'b0 : (n1876 ? !n1892 : n1892));
assign n5471 = /* LUT    5  8  1 */ (n564 ? (n5 ? 1'b0 : (n542 ? 1'b0 : !n712)) : !n712);
assign n5472 = /* LUT    4  4  0 */ (n520 ? (n232 ? !n379 : 1'b0) : n232);
assign n5473 = /* LUT   16 18  2 */ n2416;
assign n5474 = /* LUT    4  7  5 */ (n213 ? (n693 ? (n200 ? !n687 : 1'b0) : (n200 ? 1'b0 : !n687)) : (n200 ? !n687 : 1'b0));
assign n5475 = /* LUT   14 10  5 */ (n1454 ? (n2049 ? 1'b0 : !n1888) : (n2049 ? 1'b0 : n1888));
assign n5476 = /* LUT    8 11  4 */ (n1018 ? (n1145 ? (n1014 ? 1'b0 : n1015) : n1015) : (n1014 ? 1'b0 : n1015));
assign n5477 = /* LUT   14  2  1 */ (n1861 ? n1550 : 1'b0);
assign n5478 = /* LUT   16 21  7 */ (n2293 ? (n2298 ? (n2156 ? 1'b0 : !n2297) : 1'b0) : 1'b0);
assign n5479 = /* LUT   23  8  2 */ (n3015 ? 1'b0 : (n2947 ? n2945 : 1'b0));
assign n5482 = /* LUT   17  9  1 */ n1789;
assign n5483 = /* LUT    5 12  7 */ (n580 ? n579 : 1'b0);
assign n5484 = /* LUT    5  4  3 */ (n6 ? (n41 ? 1'b0 : n222) : (n41 ? n222 : 1'b0));
assign n5485 = /* LUT    4  8  6 */ (n44 ? (n212 ? n51 : 1'b0) : (n212 ? (n51 ? n548 : !n548) : 1'b0));
assign n5486 = /* LUT   16 14  4 */ (n212 ? 1'b0 : (n2129 ? !n2128 : 1'b0));
assign n5487 = /* LUT   17 10  2 */ (n2511 ? (n1765 ? n1618 : !n1618) : (n1765 ? !n1618 : n1618));
assign n5488 = /* LUT   14  6  7 */ n179;
assign n5489 = /* LUT    3 21  0 */ (n277 ? (n482 ? 1'b1 : !n487) : (n482 ? (n487 ? !n333 : 1'b1) : !n487));
assign n5490 = /* LUT    8  3  5 */ n188;
assign n5491 = /* LUT    1 21  7 */ (n152 ? (n154 ? 1'b0 : n335) : (n154 ? (n153 ? 1'b0 : n335) : n335));
assign n5492 = /* LUT   15  2  5 */ (n1555 ? (n1875 ? 1'b0 : (n2044 ? n2047 : 1'b0)) : (n2044 ? n2047 : 1'b0));
assign n5493 = /* LUT   18 23  1 */ n2012;
assign n5494 = /* LUT    1 13  3 */ (n96 ? 1'b0 : n99);
assign n5495 = /* LUT   20 17  7 */ (n2297 ? (n2855 ? (n2156 ? n2293 : 1'b0) : 1'b0) : 1'b0);
assign n5496 = /* LUT   14  3  1 */ n233;
assign n5497 = /* LUT   12 23  4 */ (n1855 ? (n5 ? 1'b0 : (n1835 ? n1659 : 1'b1)) : (n5 ? 1'b0 : (n1835 ? n1659 : 1'b0)));
assign n5498 = /* LUT   13 19  2 */ (n2001 ? !n1553 : n1553);
assign n5499 = /* LUT    7  7  6 */ (n986 ? (n853 ? 1'b0 : (n871 ? n857 : 1'b0)) : 1'b0);
assign n5500 = /* LUT    1 14  4 */ (n225 ? !n115 : (n108 ? !n115 : 1'b0));
assign n5501 = /* LUT   16  6  5 */ n177;
assign n5505 = /* LUT   10 20  5 */ (n1380 ? (n5 ? 1'b0 : (n80 ? 1'b0 : n354)) : (n5 ? 1'b0 : n354));
assign n5506 = /* LUT   10 12  1 */ (n1181 ? 1'b0 : !n1326);
assign n5507 = /* LUT    9  8  0 */ (n811 ? 1'b0 : !n209);
assign n5508 = /* LUT   13 20  3 */ (n2014 ? (n1649 ? n8 : !n8) : (n1649 ? !n8 : n8));
assign n5509 = /* LUT    7  8  7 */ (n981 ? !n871 : 1'b0);
assign n5510 = /* LUT   18 18  7 */ (n2574 ? n2408 : (n2562 ? n2408 : (n2406 ? n2408 : 1'b0)));
assign n5511 = /* LUT   20 10  3 */ n1965;
assign n5512 = /* LUT   16  2  7 */ n189;
assign n5513 = /* LUT   12 16  0 */ (n1800 ? (n1349 ? 1'b1 : (n1791 ? 1'b1 : n1783)) : (n1349 ? 1'b1 : (n1791 ? !n1783 : 1'b0)));
assign n5514 = /* LUT    3 17  7 */ (n466 ? 1'b0 : (n257 ? 1'b0 : (n584 ? 1'b0 : !n159)));
assign n5515 = /* LUT   10 16  7 */ (n1457 ? 1'b0 : n1362);
assign n5516 = /* LUT   22 19  0 */ (n2986 ? (n2293 ? (n2297 ? 1'b0 : !n2156) : 1'b0) : 1'b0);
assign n5517 = /* LUT    9 12  6 */ (n806 ? n1179 : 1'b0);
assign n5518 = /* LUT    5 18  0 */ (n786 ? (n188 ? n631 : 1'b0) : (n188 ? (n631 ? 1'b1 : n774) : n774));
assign n5519 = /* LUT   11 21  3 */ (n426 ? (n1069 ? 1'b0 : n1524) : (n1069 ? 1'b0 : (n1522 ? n1524 : 1'b0)));
assign n5520 = /* LUT   12 11  7 */ (n1329 ? (n1466 ? 1'b1 : (n1330 ? 1'b1 : !n1475)) : (n1466 ? (n1330 ? 1'b1 : !n1475) : 1'b1));
assign n5521 = /* LUT   13  7  5 */ (n1876 ? (n1691 ? 1'b0 : !n1706) : (n1691 ? 1'b0 : n1706));
assign n5522 = /* LUT    3 10  4 */ (n45 ? (n92 ? (n79 ? 1'b0 : !n419) : 1'b0) : 1'b0);
assign n5523 = /* LUT    3  2  0 */ (n371 ? n51 : 1'b0);
assign n5524 = /* LUT   18 11  3 */ (n2508 ? (n2355 ? n2369 : (n2639 ? 1'b0 : n2369)) : (n2355 ? n2369 : (n2639 ? !n2369 : 1'b1)));
assign n5525 = /* LUT    1  2  7 */ n11;
assign n5526 = /* LUT   12  8  1 */ (n1271 ? (n1569 ? 1'b0 : (n1290 ? 1'b1 : n1452)) : (n1569 ? 1'b0 : (n1290 ? 1'b1 : !n1452)));
assign n5527 = /* LUT   15 16  2 */ (n2276 ? (n2128 ? 1'b0 : n1623) : (n2128 ? n1623 : 1'b0));
assign n5528 = /* LUT    9  4  7 */ (n1110 ? (n6 ? !n41 : (n1113 ? n41 : 1'b1)) : (n6 ? 1'b1 : (n1113 ? n41 : 1'b1)));
assign n5529 = /* LUT   22 14  6 */ (n3029 ? (n8 ? n2969 : !n2969) : (n8 ? !n2969 : n2969));
assign n5530 = /* LUT    2 14  5 */ (n91 ? (n117 ? 1'b0 : !n128) : (n117 ? 1'b0 : (n297 ? !n128 : 1'b1)));
assign n5531 = /* LUT   13  8  6 */ (n1689 ? !n1465 : (n1592 ? (n1465 ? 1'b0 : n1887) : (n1465 ? 1'b0 : !n1887)));
assign n5532 = /* LUT   21 10  5 */ n2628;
assign n5533 = /* LUT   21  2  1 */ io_19_0_1;
assign n5534 = /* LUT   11 13  4 */ n189;
assign n5535 = /* LUT   11  5  0 */ (n1106 ? (n1264 ? 1'b0 : n1539) : 1'b0);
assign n5536 = /* LUT    5 19  0 */ (n630 ? !n642 : n642);
assign n5537 = /* LUT   10  1  5 */ n189;
assign n5538 = /* LUT   12 12  7 */ (n1330 ? 1'b0 : n1474);
assign n5539 = /* LUT   22 15  7 */ (n2973 ? 1'b0 : (n3019 ? 1'b0 : (n2969 ? 1'b0 : !n2974)));
assign n5540 = /* LUT    2 15  6 */ (n287 ? (n290 ? 1'b1 : n443) : 1'b0);
assign n5541 = /* LUT   12  4  3 */ (n1540 ? 1'b0 : (n1423 ? (n1419 ? n1539 : 1'b0) : 1'b1));
assign n5542 = /* LUT   22  7  3 */ (n2940 ? (n2691 ? n2622 : !n2622) : (n2691 ? !n2793 : n2793));
assign n5543 = /* LUT    2  7  2 */ (n218 ? (n220 ? n397 : (n6 ? n397 : 1'b0)) : 1'b0);
assign n5544 = /* LUT   21 11  6 */ n1755;
assign n5545 = /* LUT   21  3  2 */ (n2903 ? (n8 ? n2762 : !n2762) : (n8 ? !n2762 : n2762));
assign n5546 = /* LUT   11  6  1 */ (n1566 ? !n5 : 1'b0);
assign n5547 = /* LUT    5 14  7 */ (n4 ? (n698 ? n816 : 1'b0) : 1'b0);
assign n5548 = /* LUT    8 21  7 */ (n928 ? 1'b1 : (n1064 ? (n1066 ? 1'b0 : !n1072) : 1'b0));
assign n5549 = /* LUT   17 20  6 */ (n2022 ? 1'b0 : (n2426 ? (n2292 ? 1'b0 : !n2427) : 1'b0));
assign n5550 = /* LUT   15  4  5 */ (n1903 ? (n1836 ? (n1874 ? 1'b0 : !n1543) : !n1543) : (n1836 ? !n1874 : 1'b1));
assign n5551 = /* LUT    5  6  2 */ (n809 ? (n52 ? (n693 ? 1'b0 : !n542) : (n693 ? 1'b1 : n542)) : (n52 ? (n693 ? 1'b0 : n542) : (n693 ? 1'b1 : !n542)));
assign n5552 = /* LUT    4 10  5 */ n177;
assign n5553 = /* LUT   14 13  5 */ (n1944 ? (n2119 ? (n1494 ? 1'b1 : n1772) : (n1494 ? 1'b0 : n1772)) : (n2119 ? n1494 : (n1494 ? 1'b0 : !n1772)));
assign n5554 = /* LUT    4  2  1 */ (n495 ? (n511 ? !n176 : 1'b0) : 1'b0);
assign n5555 = /* LUT    8 14  4 */ (n1044 ? (n910 ? n1040 : 1'b0) : (n910 ? 1'b0 : n1040));
assign n5556 = /* LUT   14  5  1 */ (n1410 ? (n1888 ? 1'b0 : (n1901 ? !n956 : 1'b1)) : (n1901 ? !n956 : 1'b1));
assign n5557 = /* LUT   16 24  7 */ n2012;
assign n5558 = /* LUT   16 16  3 */ (n1 ? 1'b1 : !n1807);
assign n5564 = /* LUT    5 15  7 */ (n449 ? (n597 ? n603 : 1'b0) : n603);
assign n5565 = /* LUT    5  7  3 */ n189;
assign n5568 = /* LUT    4 11  6 */ (n270 ? (n62 ? 1'b1 : n88) : 1'b0);
assign n5569 = /* LUT    4  3  2 */ (n176 ? (n517 ? (n504 ? 1'b0 : n200) : n200) : 1'b0);
assign n5572 = /* LUT   16  9  0 */ (n2364 ? (n2085 ? 1'b0 : !n2355) : (n1927 ? 1'b0 : !n2355));
assign n5573 = /* LUT   20 21  3 */ (n2291 ? (n2748 ? 1'b1 : n2404) : (n2748 ? !n2404 : 1'b0));
assign n5574 = /* LUT   14  9  7 */ n1965;
assign n5575 = /* LUT   17 13  2 */ (n2537 ? !n2385 : n2385);
assign n5576 = /* LUT    8  6  5 */ (n891 ? (n1122 ? n1106 : (n1106 ? n983 : 1'b0)) : (n1106 ? n983 : 1'b0));
assign n5577 = /* LUT   15  5  5 */ (n1541 ? (n1125 ? (n1416 ? 1'b0 : !n1126) : 1'b0) : 1'b0);
assign n5578 = /* LUT   20 20  7 */ (n2406 ? n2408 : (n2744 ? n2408 : (n2408 ? n2434 : 1'b0)));
assign n5579 = /* LUT    7 11  2 */ (n567 ? n811 : (n811 ? !n711 : 1'b0));
assign n5580 = /* LUT   10 15  2 */ (n984 ? 1'b0 : n1488);
assign n5581 = /* LUT   16 10  1 */ (n2228 ? (n2355 ? (n2366 ? 1'b0 : n2216) : !n2366) : (n2355 ? (n2366 ? 1'b0 : n2216) : 1'b0));
assign n5582 = /* LUT   13 22  2 */ (n1856 ? (n1660 ? !n5 : (n5 ? 1'b0 : !n1835)) : (n1660 ? (n5 ? 1'b0 : n1835) : 1'b0));
assign n5585 = /* LUT   14  2  4 */ (n2045 ? (n1678 ? (n1867 ? !n1875 : 1'b0) : n1867) : 1'b0);
assign n5586 = /* LUT    1 17  4 */ (n123 ? (n307 ? !n126 : 1'b0) : (n307 ? n126 : 1'b0));
assign n5587 = /* LUT    1  9  0 */ (n53 ? (n66 ? 1'b0 : n240) : (n66 ? n240 : 1'b0));
assign n5588 = /* LUT    8  2  7 */ (n951 ? (n947 ? 1'b1 : n841) : (n947 ? (n5 ? 1'b1 : !n841) : (n5 ? n841 : 1'b0)));
assign n5592 = /* LUT   12 19  1 */ (n5 ? 1'b0 : (n1646 ? n1824 : n1817));
assign n5593 = /* LUT    7  3  3 */ (n958 ? n960 : 1'b0);
assign n5594 = /* LUT   10 11  4 */ (n1163 ? 1'b0 : (n1287 ? 1'b0 : n1310));
assign n5595 = /* LUT   18 21  7 */ n2012;
assign n5596 = /* LUT    9 15  7 */ (n642 ? (n1028 ? (n1022 ? n334 : !n334) : 1'b0) : (n1028 ? 1'b0 : (n1022 ? n334 : !n334)));
assign n5597 = /* LUT    1 10  1 */ (n69 ? 1'b0 : !n75);
assign n5598 = /* LUT   13 18  4 */ (n1814 ? (n1822 ? 1'b0 : !n1836) : 1'b0);
assign n5599 = /* LUT    3 21  3 */ (n277 ? !n484 : (n484 ? 1'b0 : !n437));
assign n5600 = /* LUT    1 13  6 */ (n273 ? 1'b0 : !n5);
assign n5601 = /* LUT   16  5  7 */ (n1931 ? 1'b0 : (n1892 ? !n1700 : n1700));
assign n5602 = /* LUT   17  1  5 */ n2194;
assign n5603 = /* LUT   20  9  6 */ n1965;
assign n5604 = /* LUT   18 14  4 */ n2651;
assign n5605 = /* LUT    9  7  2 */ (n973 ? (n852 ? 1'b1 : (n1126 ? 1'b1 : !n1125)) : 1'b1);
assign n5606 = /* LUT   13 11  1 */ n1598;
assign n5607 = /* LUT   21 21  4 */ (n2404 ? (n3002 ? (n2870 ? 1'b0 : !n2403) : (n2870 ? n2403 : 1'b1)) : n2403);
assign n5608 = /* LUT    2 17  6 */ (n126 ? (n122 ? n123 : 1'b0) : 1'b0);
assign n5609 = /* LUT   13 10  5 */ n1741;
assign n5612 = /* LUT    3  5  0 */ (n5 ? n362 : (n380 ? (n389 ? n362 : 1'b1) : (n389 ? 1'b0 : !n362)));
assign n5613 = /* LUT   10  4  0 */ (n1260 ? (n1249 ? (n5 ? 1'b0 : !n1235) : 1'b1) : 1'b0);
assign n5614 = /* LUT    1  5  7 */ n26;
assign n5615 = /* LUT   15 19  2 */ n2288;
assign n5616 = /* LUT   22 18  2 */ (n2403 ? (n3039 ? !n2404 : 1'b0) : (n2994 ? !n2404 : 1'b0));
assign n5617 = /* LUT   10  3  4 */ (n1403 ? (n1409 ? !n6 : (n6 ? !n41 : 1'b1)) : (n1409 ? (n6 ? n41 : 1'b1) : 1'b1));
assign n5618 = /* LUT   21 14  1 */ (n2829 ? (n2832 ? 1'b0 : (n2825 ? n2818 : 1'b0)) : (n2832 ? (n2825 ? 1'b0 : n2818) : n2818));
assign n5619 = /* LUT   12  7  4 */ (n1730 ? (n1703 ? !n1572 : (n1570 ? !n1572 : 1'b0)) : (n1703 ? !n1572 : (n1570 ? 1'b0 : !n1572)));
assign n5620 = /* LUT   13  3  2 */ (n1671 ? (n1874 ? !n1648 : 1'b1) : 1'b0);
assign n5621 = /* LUT   21 13  5 */ (n2827 ? 1'b1 : n2841);
assign n5622 = /* LUT    3  6  1 */ (n6 ? (n41 ? 1'b0 : n410) : (n41 ? 1'b0 : n542));
assign n5623 = /* LUT    4 21  5 */ (n800 ? !n620 : n620);
assign n5624 = /* LUT   11  8  0 */ n212;
assign n5625 = /* LUT   15 20  3 */ (n8 ? (n1822 ? n1836 : !n1836) : (n1822 ? !n1836 : n1836));
assign n5626 = /* LUT    3  9  6 */ (n414 ? (n408 ? (n53 ? n418 : 1'b0) : 1'b0) : (n408 ? (n53 ? 1'b0 : n418) : 1'b0));
assign n5627 = /* LUT   17 23  1 */ n2012;
assign n5628 = /* LUT   22 10  3 */ (n2952 ? (n2951 ? 1'b0 : (n2066 ? n2950 : 1'b0)) : 1'b0);
assign n5629 = /* LUT    2 10  2 */ (n106 ? 1'b1 : !n249);
assign n5630 = /* LUT    5 18  3 */ (n630 ? (n627 ? (n648 ? !n642 : 1'b0) : 1'b0) : (n627 ? (n648 ? n642 : 1'b0) : 1'b0));
assign n5631 = /* LUT   21  6  2 */ n2609;
assign n5632 = /* LUT   18  2  7 */ (n2440 ? 1'b0 : !n2441);
assign n5633 = /* LUT   21  9  7 */ n2192;
assign n5634 = /* LUT   17 24  2 */ n2012;
assign n5635 = /* LUT   11 12  6 */ n45;
assign n5636 = /* LUT   12  8  4 */ n188;
assign n5637 = /* LUT   11  4  2 */ (n852 ? n975 : 1'b0);
assign n5638 = /* LUT    3  1  7 */ n179;
assign n5639 = /* LUT   22  3  0 */ (n2899 ? 1'b0 : (n2896 ? 1'b0 : (n3005 ? 1'b0 : !n2897)));
assign n5640 = /* LUT    4 14  1 */ (n596 ? 1'b0 : (n297 ? 1'b0 : (n103 ? 1'b0 : !n594)));
assign n5643 = /* LUT   22  6  5 */ (n2936 ? !n2916 : 1'b0);
assign n5644 = /* LUT    5 10  4 */ n728;
assign n5645 = /* LUT   21  2  4 */ (n2757 ? !io_19_0_1 : n2889);
assign n5646 = /* LUT    7 21  6 */ (n354 ? n1031 : 1'b0);
assign n5652 = /* LUT   18  3  7 */ (n2066 ? n2454 : (n2343 ? !n2178 : n2178));
assign n5653 = /* LUT   15  8  6 */ (n2169 ? 1'b0 : (n2179 ? !n1597 : n1597));
assign n5657 = /* LUT    4  6  2 */ (n371 ? (n374 ? n372 : (n685 ? 1'b0 : n372)) : (n685 ? 1'b0 : n372));
assign n5658 = /* LUT    8 10  1 */ (n750 ? (n564 ? 1'b0 : !n711) : (n564 ? 1'b0 : (n698 ? 1'b0 : !n711)));
assign n5659 = /* LUT   16 20  4 */ n2012;
assign n5660 = /* LUT   16 12  0 */ (n2245 ? n1790 : (n2247 ? !n1790 : 1'b1));
assign n5661 = /* LUT   14 12  7 */ (n2105 ? (n1753 ? 1'b1 : !n1770) : (n1942 ? (n1753 ? n1770 : 1'b0) : (n1753 ? 1'b1 : !n1770)));
assign n5662 = /* LUT   14  4  3 */ (n1422 ? (n1428 ? 1'b0 : n1865) : n1865);
assign n5663 = /* LUT    5  3  0 */ n188;
assign n5664 = /* LUT   23  3  2 */ n3048;
assign n5665 = /* LUT   17 12  5 */ (n2378 ? (n2237 ? !n1329 : 1'b1) : (n2237 ? !n1329 : 1'b0));
assign n5666 = /* LUT   17  4  1 */ n2170;
assign n5667 = /* LUT    5  6  5 */ (n5 ? (n564 ? 1'b0 : !n712) : (n564 ? (n712 ? 1'b0 : !n695) : !n712));
assign n5668 = /* LUT   16 13  1 */ (n2251 ? n2254 : 1'b0);
assign n5669 = /* LUT    4  2  4 */ (n356 ? (n41 ? (n6 ? 1'b1 : !n381) : n6) : (n41 ? (n6 ? 1'b1 : !n381) : 1'b1));
assign n5670 = /* LUT    7  6  4 */ (n698 ? (n5 ? 1'b1 : n541) : n850);
assign n5671 = /* LUT   14  5  4 */ (n1914 ? (n1249 ? 1'b0 : n1879) : n1879);
assign n5672 = /* LUT   16 16  6 */ n2268;
assign n5673 = /* LUT    1 12  0 */ (n272 ? (n110 ? (n252 ? !n117 : 1'b0) : n252) : 1'b0);
assign n5674 = /* LUT    8  5  7 */ (n806 ? !n5 : 1'b0);
assign n5675 = /* LUT   20  8  0 */ n2798;
assign n5676 = /* LUT   12 22  1 */ (n1846 ? !n1528 : n1528);
assign n5677 = /* LUT   20 11  5 */ (n2704 ? (n2705 ? (n2699 ? 1'b0 : !n2701) : !n2701) : (n2705 ? !n2699 : 1'b1));
assign n5678 = /* LUT   10 14  4 */ (n1342 ? !n1457 : 1'b0);
assign n5681 = /* LUT    9 10  3 */ (n362 ? (n698 ? 1'b0 : !n1022) : !n698);
assign n5682 = /* LUT   22 20  2 */ (n2156 ? (n2293 ? 1'b0 : (n2297 ? n2296 : 1'b0)) : 1'b0);
assign n5683 = /* LUT    7  2  6 */ (n52 ? (n829 ? 1'b0 : n832) : n832);
assign n5684 = /* LUT   21 16  1 */ (n2983 ? (n2404 ? (n2550 ? 1'b1 : n2406) : 1'b0) : (n2404 ? (n2550 ? !n2406 : 1'b0) : 1'b0));
assign n5685 = /* LUT   16  8  7 */ n1938;
assign n5686 = /* LUT   20 12  6 */ (n2500 ? 1'b0 : (n2509 ? 1'b0 : n2809));
assign n5687 = /* LUT   10 15  5 */ (n1268 ? (n1358 ? 1'b1 : n984) : 1'b0);
assign n5688 = /* LUT   10  7  1 */ (n1290 ? (n1146 ? !n1267 : 1'b0) : (n1146 ? (n5 ? 1'b1 : !n1267) : 1'b0));
assign n5689 = /* LUT   18  9  0 */ (n2366 ? (n2492 ? 1'b0 : !n2493) : n2497);
assign n5690 = /* LUT   22 21  3 */ n2012;
assign n5691 = /* LUT    2 21  2 */ (n491 ? (n150 ? !n325 : 1'b0) : (n150 ? n325 : 1'b0));
assign n5692 = /* LUT   20  5  3 */ (n2675 ? !n2674 : n2674);
assign n5696 = /* LUT    1  8  7 */ (n54 ? (n69 ? n235 : 1'b0) : 1'b0);
assign n5697 = /* LUT   18 10  1 */ (n2630 ? (n2364 ? (n2355 ? !n2479 : 1'b1) : 1'b0) : (n2364 ? (n2355 ? !n2479 : 1'b1) : n2355));
assign n5698 = /* LUT   12 11  0 */ (n1609 ? 1'b0 : (n1637 ? (n1477 ? n1608 : 1'b0) : 1'b0));
assign n5699 = /* LUT   21 17  1 */ (n2848 ? (n2156 ? 1'b0 : (n2297 ? 1'b0 : !n2293)) : 1'b0);
assign n5700 = /* LUT   12 10  4 */ n175;
assign n5701 = /* LUT   13  6  2 */ (n1704 ? !n1037 : (n1696 ? (n1892 ? !n1037 : 1'b0) : (n1892 ? 1'b0 : !n1037)));
assign n5702 = /* LUT   10  2  7 */ n175;
assign n5706 = /* LUT   13  9  7 */ n1752;
assign n5707 = /* LUT   14 19  1 */ (n2147 ? (n2009 ? n1956 : !n1956) : (n2009 ? !n1956 : n1956));
assign n5708 = /* LUT    3 12  6 */ (n259 ? (n132 ? 1'b0 : !n257) : (n132 ? 1'b0 : (n391 ? 1'b0 : !n257)));
assign n5709 = /* LUT    3  4  2 */ n188;
assign n5710 = /* LUT   15 18  4 */ n2282;
assign n5713 = /* LUT   24 17  3 */ n2012;
assign n5714 = /* LUT    4 17  2 */ (n142 ? (n462 ? !n772 : 1'b0) : n462);
assign n5715 = /* LUT   18  5  7 */ n2173;
assign n5716 = /* LUT    2  9  5 */ (n60 ? (n53 ? (n63 ? n66 : 1'b0) : (n63 ? 1'b0 : n66)) : (n53 ? (n63 ? !n66 : 1'b0) : (n63 ? 1'b0 : !n66)));
assign n5717 = /* LUT   13  2  4 */ (n1478 ? n1550 : 1'b0);
assign n5718 = /* LUT    3  5  3 */ (n364 ? 1'b0 : (n203 ? (n52 ? 1'b1 : !n384) : 1'b0));
assign n5719 = /* LUT   11 15  6 */ (n1195 ? 1'b1 : (n1464 ? n1033 : 1'b0));
assign n5720 = /* LUT   16 23  0 */ (n2293 ? (n2297 ? 1'b0 : (n2296 ? n2156 : 1'b0)) : 1'b0);
assign n5721 = /* LUT   11  7  2 */ (n1271 ? (n1565 ? n841 : 1'b1) : (n1565 ? 1'b0 : !n841));
assign n5722 = /* LUT    8 20  5 */ (n1031 ? (n1063 ? (n189 ? 1'b1 : n925) : n189) : (n1063 ? n925 : 1'b0));
assign n5723 = /* LUT   15 19  5 */ n2012;
assign n5724 = /* LUT   15 11  1 */ (n1892 ? (n2238 ? (n2233 ? !n2239 : 1'b1) : 1'b0) : (n2238 ? (n2233 ? 1'b0 : n2239) : 1'b0));
assign n5725 = /* LUT   10  3  7 */ (n1257 ? (n1410 ? 1'b1 : n1408) : (n1410 ? n5 : n1408));
assign n5726 = /* LUT   23 21  4 */ n2012;
assign n5727 = /* LUT    5 14  0 */ (n752 ? (n439 ? !n578 : 1'b0) : (n439 ? (n604 ? !n578 : 1'b0) : 1'b0));
assign n5728 = /* LUT   12  7  7 */ (n1573 ? (n1731 ? (n956 ? 1'b0 : !n1410) : !n956) : (n1731 ? !n1410 : 1'b1));
assign n5729 = /* LUT   21  5  4 */ (n2933 ? (n2780 ? n8 : !n8) : (n2780 ? !n8 : n8));
assign n5730 = /* LUT   11  8  3 */ (n1146 ? (n1267 ? (n5 ? !n1301 : 1'b0) : 1'b1) : 1'b0);
assign n5731 = /* LUT   23 14  1 */ (n2819 ? !n2827 : 1'b0);
assign n5732 = /* LUT    8 16  7 */ !n1050;
assign n5733 = /* LUT   15  3  2 */ n188;
assign n5734 = /* LUT   22  2  2 */ (n2757 ? 1'b1 : n2889);
assign n5735 = /* LUT   17 14  4 */ (n2547 ? !n2265 : n2265);
assign n5736 = /* LUT    7 17  3 */ !n620;
assign n5737 = /* LUT   15  6  7 */ (n1901 ? (n1923 ? 1'b0 : !n1727) : (n1923 ? !n1727 : 1'b0));
assign n5738 = /* LUT    8 13  1 */ n189;
assign n5739 = /* LUT    2  1  5 */ n233;
assign n5740 = /* LUT    5  9  6 */ (n562 ? (n700 ? 1'b0 : (n723 ? n715 : 1'b0)) : n723);
assign n5741 = /* LUT    4  5  5 */ (n401 ? (n6 ? 1'b0 : !n396) : (n6 ? 1'b1 : !n396));
assign n5742 = /* LUT   14  7  3 */ (n1678 ? 1'b0 : (n1926 ? !n1573 : n1573));
assign n5743 = /* LUT   16 19  7 */ (n1987 ? (n2285 ? (n2144 ? n1823 : 1'b0) : (n2144 ? 1'b1 : !n1823)) : (n2285 ? (n2144 ? !n1823 : 1'b1) : (n2144 ? 1'b0 : n1823)));
assign n5744 = /* LUT   23  6  2 */ n2936;
assign n5745 = /* LUT   17  7  1 */ n2485;
assign n5748 = /* LUT    5 10  7 */ (n711 ? (n64 ? 1'b0 : n811) : n811);
assign n5749 = /* LUT    9 21  2 */ (n1218 ? 1'b0 : (n924 ? 1'b0 : (n1069 ? 1'b1 : n437)));
assign n5750 = /* LUT   20 20  0 */ (n2297 ? 1'b0 : (n2855 ? (n2293 ? 1'b0 : n2156) : 1'b0));
assign n5751 = /* LUT   14  8  4 */ (n1918 ? 1'b0 : (n1906 ? 1'b0 : (n1919 ? 1'b0 : !n1922)));
assign n5752 = /* LUT    8  9  3 */ (n1148 ? !n876 : n876);
assign n5753 = /* LUT   13 16  1 */ (n1983 ? 1'b1 : n1126);
assign n5754 = /* LUT    8  8  7 */ (n985 ? (n866 ? (n873 ? n870 : 1'b0) : (n873 ? 1'b0 : n870)) : (n866 ? (n873 ? !n870 : 1'b0) : (n873 ? 1'b0 : !n870)));
assign n5758 = /* LUT    5  2  2 */ n179;
assign n5761 = /* LUT   10 17  4 */ n15;
assign n5762 = /* LUT    9 13  3 */ (n806 ? n1050 : 1'b0);
assign n5763 = /* LUT   16 12  3 */ (n1891 ? (n2239 ? (n2358 ? 1'b0 : n2238) : n2238) : (n2239 ? (n2358 ? 1'b0 : n2238) : 1'b0));
assign n5764 = /* LUT   13 17  2 */ n1988;
assign n5765 = /* LUT    7  5  6 */ (n390 ? (n846 ? 1'b1 : n698) : (n846 ? (n5 ? 1'b1 : !n698) : (n5 ? n698 : 1'b0)));
assign n5766 = /* LUT    8  1  4 */ n189;
assign n5767 = /* LUT    1 19  6 */ (n93 ? (n142 ? (n139 ? !n150 : 1'b1) : !n150) : !n150);
assign n5768 = /* LUT    1 11  2 */ (n89 ? (n70 ? (n258 ? 1'b0 : !n75) : !n258) : (n70 ? !n75 : 1'b1));
assign n5769 = /* LUT   20  7  2 */ n2795;
assign n5770 = /* LUT   10 10  1 */ (n812 ? (n811 ? n1146 : 1'b0) : n1146);
assign n5771 = /* LUT   12 21  3 */ (n1840 ? !n1832 : n1832);
assign n5772 = /* LUT    7  6  7 */ (n5 ? (n698 ? 1'b1 : n848) : (n698 ? n527 : n848));
assign n5773 = /* LUT   10 13  6 */ (n1328 ? (n1459 ? n1349 : (n1349 ? !n212 : 1'b0)) : (n1459 ? n1349 : 1'b0));
assign n5774 = /* LUT    3 20  0 */ (n631 ? (n478 ? n233 : (n489 ? 1'b1 : n233)) : (n478 ? 1'b0 : n489));
assign n5775 = /* LUT   21 20  2 */ (n2404 ? n2874 : (n2999 ? (n2860 ? 1'b0 : !n2874) : (n2860 ? n2874 : 1'b1)));
assign n5776 = /* LUT    9  9  5 */ (n1285 ? (n1129 ? 1'b0 : !n1155) : 1'b0);
assign n5779 = /* LUT   21 23  7 */ (n2296 ? (n2156 ? 1'b0 : (n2297 ? n2293 : 1'b0)) : 1'b0);
assign n5780 = /* LUT   12 22  4 */ (n1852 ? !n1848 : n1848);
assign n5781 = /* LUT   18 13  1 */ n2649;
assign n5785 = /* LUT   10  6  3 */ (n852 ? 1'b1 : !n975);
assign n5786 = /* LUT   18 16  6 */ n2410;
assign n5787 = /* LUT    9  2  2 */ (n176 ? 1'b0 : (n1098 ? n1252 : 1'b0));
assign n5788 = /* LUT   21 16  4 */ (n2406 ? (n2847 ? !n2404 : 1'b1) : (n2723 ? 1'b0 : n2404));
assign n5789 = /* LUT    3 15  6 */ (n303 ? 1'b0 : (n446 ? 1'b0 : (n91 ? 1'b0 : !n452)));
assign n5790 = /* LUT    3  7  2 */ n188;
assign n5791 = /* LUT   11 10  3 */ (n1457 ? !n212 : (n1459 ? 1'b0 : !n212));
assign n5792 = /* LUT   18  9  3 */ (n2355 ? 1'b0 : (n2491 ? (n2370 ? 1'b1 : !n2364) : (n2370 ? n2364 : 1'b0)));
assign n5793 = /* LUT   12  6  1 */ (n1695 ? (n1570 ? 1'b1 : !n956) : (n1570 ? n956 : 1'b0));
assign n5794 = /* LUT   15 13  0 */ (n2104 ? (n1728 ? n1892 : (n1892 ? !n2102 : 1'b0)) : (n1728 ? 1'b1 : !n2102));
assign n5795 = /* LUT    4 20  2 */ (n648 ? (n625 ? (n488 ? n627 : 1'b0) : (n488 ? 1'b0 : n627)) : 1'b0);
assign n5796 = /* LUT   12  9  6 */ (n423 ? (n212 ? (n1742 ? 1'b1 : !n1733) : n1742) : 1'b0);
assign n5797 = /* LUT    2 12  5 */ (n423 ? n262 : (n101 ? n262 : 1'b0));
assign n5798 = /* LUT   13  5  4 */ (n1683 ? (n1885 ? 1'b1 : !n1410) : (n1885 ? n1410 : 1'b0));
assign n5799 = /* LUT   22  4  2 */ (n2913 ? (n2900 ? (n2898 ? n2783 : 1'b0) : 1'b0) : 1'b0);
assign n5800 = /* LUT    3  8  3 */ (n556 ? (n83 ? (n227 ? 1'b0 : n43) : 1'b0) : (n83 ? (n227 ? n43 : 1'b0) : 1'b0));
assign n5801 = /* LUT    2  4  1 */ n192;
assign n5802 = /* LUT   21  8  5 */ !n2623;
assign n5803 = /* LUT   14 18  3 */ (n2141 ? (n2143 ? (n1823 ? n1995 : !n1995) : n1995) : (n2143 ? !n1995 : (n1823 ? !n1995 : n1995)));
assign n5804 = /* LUT   15 14  1 */ (n1970 ? 1'b1 : n2113);
assign n5805 = /* LUT    5 17  0 */ (n159 ? 1'b0 : (n304 ? 1'b0 : (n252 ? n292 : 1'b0)));
assign n5806 = /* LUT   12 10  7 */ n233;
assign n5807 = /* LUT   18  1  4 */ n2598;
assign n5808 = /* LUT   12  2  3 */ (n1539 ? (n1537 ? (n1425 ? !n5 : 1'b0) : !n5) : (n1537 ? 1'b0 : !n5));
assign n5809 = /* LUT    2  5  2 */ (n212 ? (n211 ? !n52 : (n52 ? n371 : 1'b1)) : 1'b0);
assign n5810 = /* LUT   24 16  5 */ n2012;
assign n5811 = /* LUT    4 16  4 */ (n455 ? n264 : (n758 ? (n264 ? n266 : 1'b0) : n264));
assign n5814 = /* LUT   14 19  4 */ (n2150 ? !n1984 : n1984);
assign n5815 = /* LUT   14 11  0 */ n1463;
assign n5816 = /* LUT   21  4  7 */ (n2923 ? (n2671 ? !n8 : n8) : (n2671 ? n8 : !n8));
assign n5819 = /* LUT   20 22  0 */ n2012;
assign n5820 = /* LUT    8 11  3 */ (n1026 ? (n698 ? 1'b0 : !n362) : !n698);
assign n5821 = /* LUT   22  5  2 */ (n2673 ? (n7 ? (n2675 ? 1'b1 : n2674) : 1'b1) : 1'b1);
assign n5822 = /* LUT   21  1  1 */ !n2314;
assign n5825 = /* LUT   15  9  7 */ (n1927 ? (n1931 ? !n2073 : (n2073 ? 1'b0 : n1700)) : (n1931 ? !n2073 : (n2073 ? 1'b0 : !n1700)));
assign n5826 = /* LUT    5 12  6 */ (n128 ? (n455 ? 1'b1 : n266) : 1'b0);
assign n5827 = /* LUT    5  4  2 */ (n506 ? (n666 ? 1'b0 : n362) : (n666 ? (n362 ? 1'b0 : n679) : (n362 ? 1'b1 : n679)));
assign n5828 = /* LUT    4  8  5 */ (n398 ? (n200 ? (n554 ? n44 : 1'b0) : (n554 ? !n44 : 1'b0)) : (n200 ? n554 : 1'b0));
assign n5829 = /* LUT   16 14  3 */ !n1766;
assign n5830 = /* LUT   17 18  5 */ (n2572 ? !n2413 : n2413);
assign n5831 = /* LUT   17 10  1 */ (n2510 ? (n1617 ? n1766 : !n1766) : (n1617 ? !n1766 : n1766));
assign n5832 = /* LUT   14  6  6 */ (n1883 ? 1'b0 : (n1893 ? !n1740 : n1740));
assign n5833 = /* LUT    7 13  0 */ (n1019 ? (n679 ? 1'b0 : !n806) : !n679);
assign n5834 = /* LUT   15  2  4 */ n233;
assign n5835 = /* LUT    5  5  3 */ n233;
assign n5836 = /* LUT    4  1  2 */ (n515 ? (n41 ? n6 : (n6 ? 1'b1 : !n658)) : (n41 ? 1'b1 : (n6 ? 1'b1 : !n658)));
assign n5837 = /* LUT   14  3  0 */ (n2049 ? (n1863 ? (n1882 ? 1'b0 : !n1543) : !n1543) : (n1863 ? !n1882 : 1'b1));
assign n5838 = /* LUT   16 15  4 */ n1323;
assign n5839 = /* LUT   16  7  0 */ (n1716 ? !n2201 : (n1877 ? (n2201 ? 1'b0 : n2069) : (n2201 ? 1'b0 : !n2069)));
assign n5840 = /* LUT   20 18  1 */ (n2858 ? (n2724 ? n2407 : 1'b0) : (n2733 ? (n2724 ? n2407 : 1'b0) : (n2724 ? 1'b1 : !n2407)));
assign n5841 = /* LUT   15  3  5 */ (n1179 ? n1543 : 1'b0);
assign n5842 = /* LUT   17 14  7 */ !n2394;
assign n5843 = /* LUT    1 14  3 */ (n109 ? (n80 ? n99 : (n99 ? n107 : 1'b0)) : (n99 ? n107 : 1'b0));
assign n5844 = /* LUT    7  9  2 */ (n1002 ? (n997 ? n8 : !n8) : (n997 ? !n8 : n8));
assign n5845 = /* LUT   13 20  2 */ (n2013 ? (n8 ? n1553 : !n1553) : (n8 ? !n1553 : n1553));
assign n5846 = /* LUT    7  8  6 */ (n995 ? (n981 ? !n870 : 1'b0) : (n981 ? n870 : 1'b0));
assign n5847 = /* LUT   14  7  6 */ (n1900 ? 1'b0 : (n1913 ? 1'b0 : (n1907 ? 1'b0 : !n1905)));
assign n5848 = /* LUT   13 23  7 */ (n1662 ? (n5 ? 1'b0 : (n1835 ? 1'b1 : n1858)) : (n5 ? 1'b0 : (n1835 ? 1'b0 : n1858)));
assign n5849 = /* LUT    3 18  2 */ (n622 ? !n461 : n461);
assign n5850 = /* LUT   10 16  6 */ (n1184 ? (n1203 ? 1'b0 : (n1370 ? 1'b1 : n212)) : (n1203 ? 1'b0 : (n1370 ? !n212 : 1'b0)));
assign n5851 = /* LUT    7  1  3 */ n189;
assign n5852 = /* LUT   18 19  7 */ (n2293 ? 1'b0 : (n2156 ? (n2297 ? 1'b0 : n2298) : 1'b0));
assign n5853 = /* LUT    9 12  5 */ (n1032 ? (n1177 ? 1'b0 : n1178) : (n1177 ? (n1178 ? n1176 : 1'b0) : n1178));
assign n5854 = /* LUT    1 15  3 */ (n93 ? 1'b1 : n5);
assign n5855 = /* LUT   13 16  4 */ n1981;
assign n5856 = /* LUT    3 19  3 */ (n633 ? !n334 : n334);
assign n5857 = /* LUT   11 21  2 */ (n80 ? !n1519 : 1'b0);
assign n5858 = /* LUT   16  3  7 */ n179;
assign n5859 = /* LUT   12 17  0 */ (n1645 ? (n1807 ? !n1643 : 1'b0) : 1'b0);
assign n5860 = /* LUT   10 17  7 */ n354;
assign n5861 = /* LUT   20  6  4 */ (n2787 ? !n2680 : n2680);
assign n5862 = /* LUT   10  9  3 */ (n1446 ? (n1288 ? (n1300 ? 1'b1 : n1447) : 1'b1) : 1'b0);
assign n5863 = /* LUT    9 13  6 */ (n642 ? !n362 : (n362 ? 1'b0 : !n679));
assign n5864 = /* LUT   18 11  2 */ (n2364 ? (n2092 ? 1'b0 : n2355) : (n2355 ? !n2353 : 1'b0));
assign n5865 = /* LUT    9  5  2 */ (n1110 ? (n1261 ? !n806 : 1'b0) : (n1112 ? !n806 : (n1261 ? !n806 : 1'b0)));
assign n5866 = /* LUT   21 19  4 */ n2012;
assign n5867 = /* LUT   13  8  5 */ (n1745 ? (n1746 ? 1'b0 : (n1917 ? !n1737 : 1'b1)) : !n1746);
assign n5868 = /* LUT   18 20  7 */ (n2296 ? (n2297 ? 1'b0 : (n2156 ? 1'b0 : !n2293)) : 1'b0);
assign n5869 = /* LUT   18 12  3 */ n2627;
assign n5870 = /* LUT   10  1  4 */ (n6 ? (n1237 ? n41 : 1'b1) : (n1239 ? !n41 : 1'b1));
assign n5871 = /* LUT   12 12  6 */ (n817 ? !n1475 : 1'b1);
assign n5872 = /* LUT   22 15  6 */ !n2976;
assign n5873 = /* LUT    2  7  1 */ (n41 ? (n6 ? (n62 ? n176 : 1'b0) : !n62) : 1'b0);
assign n5874 = /* LUT   21 11  5 */ n1938;
assign n5877 = /* LUT    1  3  6 */ (n12 ? (n9 ? (n30 ? n29 : 1'b0) : (n30 ? 1'b0 : n29)) : (n9 ? (n30 ? !n29 : 1'b0) : (n30 ? 1'b0 : !n29)));
assign n5878 = /* LUT   14 21  3 */ (n2019 ? 1'b0 : (n2025 ? (n1665 ? !n1491 : 1'b1) : 1'b1));
assign n5879 = /* LUT   11  6  0 */ (n1564 ? (n1122 ? (n983 ? 1'b1 : n1115) : n983) : 1'b0);
assign n5880 = /* LUT   13  4  7 */ (n1281 ? (n1422 ? 1'b1 : n1677) : (n1422 ? 1'b0 : n1677));
assign n5881 = /* LUT    5 20  0 */ (n794 ? 1'b1 : (n791 ? 1'b0 : (n785 ? n796 : 1'b0)));
assign n5882 = /* LUT   17 21  1 */ (n2293 ? (n2427 ? (n2297 ? n2156 : 1'b0) : 1'b0) : 1'b0);
assign n5883 = /* LUT   11  9  5 */ (n1429 ? n1267 : (n1267 ? !n5 : 1'b0));
assign n5884 = /* LUT   12 13  7 */ (n1783 ? (n1349 ? 1'b1 : n1773) : (n1349 ? 1'b1 : n1626));
assign n5885 = /* LUT   12  5  3 */ n189;
assign n5886 = /* LUT    2  8  2 */ (n411 ? (n226 ? 1'b0 : n240) : (n226 ? n240 : 1'b0));
assign n5889 = /* LUT    4 19  4 */ (n790 ? (n627 ? (n490 ? n648 : 1'b0) : 1'b0) : (n627 ? (n490 ? 1'b0 : n648) : 1'b0));
assign n5890 = /* LUT   14 22  4 */ !n2009;
assign n5891 = /* LUT    2 11  7 */ (n249 ? (n128 ? (n91 ? 1'b0 : n423) : (n91 ? 1'b1 : n423)) : 1'b0);
assign n5892 = /* LUT   14 14  0 */ (n1950 ? (n1770 ? n1556 : 1'b1) : (n1770 ? n1556 : 1'b0));
assign n5893 = /* LUT    3  7  5 */ n354;
assign n5896 = /* LUT   11 10  6 */ (n1425 ? n892 : 1'b0);
assign n5897 = /* LUT    8 22  7 */ (n1069 ? (n924 ? !n1230 : 1'b0) : (n924 ? !n1230 : (n1230 ? 1'b0 : !n437)));
assign n5898 = /* LUT   15 13  3 */ (n1624 ? 1'b0 : n2122);
assign n5899 = /* LUT    5 15  6 */ (n756 ? 1'b1 : (n753 ? 1'b0 : !n249));
assign n5900 = /* LUT   22  4  5 */ (n2774 ? 1'b0 : (n2764 ? 1'b0 : (n2773 ? 1'b0 : n2768)));
assign n5901 = /* LUT    4 11  5 */ (n729 ? n88 : 1'b0);
assign n5902 = /* LUT   11  2  1 */ n354;
assign n5908 = /* LUT   17 13  1 */ (n2257 ? !n2386 : n2386);
assign n5909 = /* LUT   20 21  2 */ n2012;
assign n5910 = /* LUT   14  9  6 */ n1754;
assign n5911 = /* LUT   15  5  4 */ n177;
assign n5912 = /* LUT    5  8  3 */ (n557 ? (n706 ? (n716 ? !n688 : 1'b0) : 1'b0) : n716);
assign n5913 = /* LUT    4  4  2 */ (n200 ? (n675 ? (n676 ? 1'b0 : !n176) : !n176) : 1'b0);
assign n5914 = /* LUT    7 11  1 */ (n711 ? 1'b1 : (n564 ? n885 : 1'b0));
assign n5915 = /* LUT   16 18  4 */ n2417;
assign n5916 = /* LUT    4  7  7 */ (n41 ? 1'b1 : (n692 ? (n6 ? !n693 : 1'b0) : (n6 ? !n693 : 1'b1)));
assign n5917 = /* LUT   16 10  0 */ n2204;
assign n5918 = /* LUT   14 10  7 */ (n1882 ? !n1935 : (n1935 ? 1'b0 : (n1763 ? n1714 : !n1714)));
assign n5919 = /* LUT    8 11  6 */ (n1061 ? (n679 ? 1'b0 : !n806) : !n679);
assign n5920 = /* LUT   14  2  3 */ n189;
assign n5921 = /* LUT    5  1  0 */ (n41 ? 1'b1 : (n6 ? !n650 : !n653));
assign n5924 = /* LUT   17  9  3 */ (n2355 ? (n2364 ? !n2502 : !n2352) : n2364);
assign n5925 = /* LUT    7 12  2 */ (n883 ? (n884 ? 1'b1 : (n738 ? !n890 : 1'b0)) : 1'b0);
assign n5926 = /* LUT    5  4  5 */ (n222 ? !n6 : 1'b0);
assign n5927 = /* LUT   16 11  1 */ n1755;
assign n5928 = /* LUT   10 19  7 */ (n1189 ? 1'b0 : (n648 ? (n1375 ? !n1050 : 1'b0) : 1'b0));
assign n5929 = /* LUT   16 14  6 */ (n1037 ? 1'b0 : (n212 ? !n2128 : 1'b0));
assign n5930 = /* LUT    9 15  6 */ (n249 ? 1'b0 : (n753 ? 1'b0 : n1144));
assign n5931 = /* LUT    1 10  0 */ (n69 ? 1'b0 : (n76 ? (n242 ? n235 : 1'b0) : 1'b0));
assign n5932 = /* LUT   17  2  0 */ (n2307 ? 1'b1 : n2320);
assign n5933 = /* LUT    3 21  2 */ (n483 ? n333 : 1'b0);
assign n5934 = /* LUT    8  3  7 */ (n5 ? (n1084 ? 1'b1 : n841) : (n1084 ? (n953 ? 1'b1 : !n841) : (n953 ? n841 : 1'b0)));
assign n5935 = /* LUT    1 13  5 */ (n106 ? n249 : 1'b0);
assign n5936 = /* LUT   12 20  1 */ (n1653 ? 1'b1 : (n1652 ? 1'b1 : (n5 ? 1'b1 : n1501)));
assign n5937 = /* LUT   20  9  5 */ (n2377 ? 1'b0 : n577);
assign n5938 = /* LUT    9  7  1 */ (n1125 ? (n892 ? (n973 ? !n1126 : 1'b0) : 1'b0) : 1'b0);
assign n5939 = /* LUT   13 19  4 */ (n2003 ? !n1715 : n1715);
assign n5940 = /* LUT   21 21  3 */ (n2156 ? (n2848 ? (n2293 ? !n2297 : 1'b0) : 1'b0) : 1'b0);
assign n5941 = /* LUT    1 14  6 */ (n110 ? n99 : (n99 ? n285 : 1'b0));
assign n5942 = /* LUT   16  6  7 */ (n1893 ? (n1705 ? 1'b0 : !n1883) : (n1705 ? !n1883 : 1'b0));
assign n5945 = /* LUT   10 20  7 */ !n1189;
assign n5946 = /* LUT   10 12  3 */ (n1338 ? (n1314 ? (n1181 ? 1'b0 : n1182) : !n1181) : (n1181 ? 1'b0 : n1182));
assign n5947 = /* LUT    9  8  2 */ n1128;
assign n5948 = /* LUT   22 18  1 */ (n2293 ? 1'b0 : (n2156 ? 1'b0 : (n2297 ? n2992 : 1'b0)));
assign n5949 = /* LUT    2 18  0 */ (n112 ? (n300 ? 1'b0 : (n309 ? 1'b0 : !n318)) : 1'b0);
assign n5950 = /* LUT   13 12  1 */ (n1772 ? n1592 : n1706);
assign n5951 = /* LUT   21 14  0 */ (n2813 ? 1'b1 : n2710);
assign n5952 = /* LUT   20 10  5 */ n1757;
assign n5953 = /* LUT    3  6  0 */ (n539 ? (n387 ? (n544 ? 1'b0 : !n200) : !n544) : 1'b0);
assign n5954 = /* LUT   10  5  0 */ (n852 ? n1425 : 1'b0);
assign n5955 = /* LUT   12 16  2 */ (n1483 ? 1'b0 : !n5);
assign n5956 = /* LUT   15 20  2 */ (n1646 ? (n2153 ? !n5 : 1'b0) : (n1816 ? !n5 : 1'b0));
assign n5957 = /* LUT    3  9  5 */ (n226 ? (n415 ? (n563 ? n66 : !n66) : 1'b0) : (n415 ? 1'b0 : (n563 ? n66 : !n66)));
assign n5958 = /* LUT    2 10  1 */ (n42 ? 1'b1 : (n128 ? n251 : 1'b0));
assign n5959 = /* LUT   18  8  0 */ n1789;
assign n5960 = /* LUT   13  7  7 */ (n1705 ? (n1691 ? !n1719 : (n1876 ? !n1719 : 1'b0)) : (n1691 ? !n1719 : (n1876 ? 1'b0 : !n1719)));
assign n5961 = /* LUT    3  2  2 */ (n351 ? (n6 ? !n41 : (n344 ? n41 : 1'b1)) : (n6 ? 1'b1 : (n344 ? n41 : 1'b1)));
assign n5962 = /* LUT   11 12  5 */ (n1475 ? !n1472 : 1'b0);
assign n5963 = /* LUT   18 11  5 */ n2638;
assign n5964 = /* LUT   12  8  3 */ (n1453 ? (n1428 ? 1'b0 : !n1575) : (n1428 ? 1'b0 : n1575));
assign n5965 = /* LUT   15 16  4 */ (n1790 ? 1'b0 : n1623);
assign n5966 = /* LUT    4 14  0 */ (n128 ? (n595 ? (n297 ? 1'b0 : n249) : 1'b0) : (n595 ? n249 : (n297 ? n249 : 1'b0)));
assign n5967 = /* LUT    2 14  7 */ (n252 ? (n151 ? n288 : 1'b0) : 1'b0);
assign n5968 = /* LUT   21  2  3 */ (n2889 ? !n2758 : 1'b0);
assign n5969 = /* LUT   11  5  2 */ (n1424 ? (n1126 ? 1'b0 : n1125) : 1'b0);
assign n5973 = /* LUT    5 19  2 */ (n631 ? (n776 ? n179 : (n793 ? 1'b1 : n179)) : (n776 ? 1'b0 : n793));
assign n5974 = /* LUT   10  1  7 */ n233;
assign n5975 = /* LUT    4 15  1 */ (n92 ? (n265 ? (n455 ? 1'b0 : n286) : 1'b0) : 1'b0);
assign n5976 = /* LUT   12  4  5 */ (n956 ? 1'b0 : (n1410 ? !n1692 : 1'b1));
assign n5977 = /* LUT   22  7  5 */ (n2693 ? (n1 ? 1'b0 : (n2936 ? n3014 : 1'b1)) : !n1);
assign n5978 = /* LUT    2  7  4 */ !n230;
assign n5979 = /* LUT   21  3  4 */ (n2905 ? (n8 ? n2764 : !n2764) : (n8 ? !n2764 : n2764));
assign n5980 = /* LUT   14 21  6 */ (n2020 ? 1'b0 : !n2155);
assign n5981 = /* LUT   11  6  3 */ n354;
assign n5982 = /* LUT    8 10  0 */ (n564 ? 1'b0 : (n757 ? !n711 : (n711 ? 1'b0 : !n698)));
assign n5983 = /* LUT   15  9  0 */ (n1596 ? (n1699 ? n2083 : (n1885 ? n2083 : 1'b0)) : (n1699 ? n2083 : (n1885 ? 1'b0 : n2083)));
assign n5984 = /* LUT   17 12  4 */ (n1632 ? (n2379 ? !n2239 : 1'b1) : (n2379 ? 1'b0 : n2239));
assign n5985 = /* LUT   17  4  0 */ n2173;
assign n5986 = /* LUT   15  4  7 */ (n1301 ? (n2050 ? !n1422 : 1'b0) : n2050);
assign n5987 = /* LUT    5  6  4 */ (n6 ? 1'b0 : n41);
assign n5988 = /* LUT    4 10  7 */ n15;
assign n5989 = /* LUT   16 13  0 */ (n2238 ? (n2122 ? 1'b0 : n2383) : (n1463 ? 1'b0 : !n2122));
assign n5990 = /* LUT   14 13  7 */ (n1951 ? (n1952 ? (n1758 ? n1946 : 1'b1) : !n1758) : (n1952 ? 1'b1 : !n1758));
assign n5991 = /* LUT    4  2  3 */ (n41 ? (n6 ? 1'b1 : !n516) : (n501 ? !n6 : 1'b1));
assign n5992 = /* LUT    8 14  6 */ (n1035 ? (n1022 ? (n1029 ? n931 : 1'b0) : (n1029 ? !n931 : 1'b0)) : 1'b0);
assign n5993 = /* LUT   14  5  3 */ n233;
assign n5999 = /* LUT    5  7  5 */ (n537 ? (n41 ? !n6 : (n6 ? !n695 : 1'b1)) : (n41 ? 1'b1 : (n6 ? !n695 : 1'b1)));
assign n6000 = /* LUT    9 19  2 */ (n907 ? (n931 ? 1'b0 : !n932) : 1'b0);
assign n6001 = /* LUT    4  3  4 */ (n507 ? (n508 ? (n662 ? 1'b0 : !n671) : 1'b1) : 1'b0);
assign n6002 = /* LUT   16  9  2 */ (n2212 ? (n2364 ? n2229 : 1'b1) : (n2364 ? n2229 : 1'b0));
assign n6003 = /* LUT   17 13  4 */ (n2539 ? !n2255 : n2255);
assign n6004 = /* LUT   17  5  0 */ n2331;
assign n6005 = /* LUT   20 13  1 */ (n2500 ? (n2817 ? !n2534 : 1'b1) : (n2532 ? !n2817 : 1'b1));
assign n6006 = /* LUT    8  6  7 */ (n978 ? n1106 : (n841 ? (n1106 ? n816 : 1'b0) : 1'b0));
assign n6007 = /* LUT   15  5  7 */ (n1541 ? (n1126 ? 1'b0 : (n1416 ? n1125 : 1'b0)) : 1'b0);
assign n6008 = /* LUT   10 15  4 */ (n1360 ? (n212 ? (n1186 ? n1477 : 1'b0) : n1477) : (n212 ? (n1186 ? n1477 : 1'b0) : 1'b0));
assign n6009 = /* LUT   10  7  0 */ (n876 ? !n1267 : (n811 ? !n1267 : (n1267 ? 1'b0 : !n5)));
assign n6010 = /* LUT   13 22  4 */ (n1857 ? (n1835 ? (n5 ? 1'b0 : n1661) : !n5) : (n1835 ? (n5 ? 1'b0 : n1661) : 1'b0));
assign n6011 = /* LUT    2 21  1 */ (n331 ? (n324 ? 1'b0 : n150) : (n324 ? n150 : 1'b0));
assign n6012 = /* LUT   13 14  0 */ (n1330 ? (n1494 ? 1'b1 : n1741) : (n1494 ? 1'b0 : n1741));
assign n6013 = /* LUT    1 17  6 */ (n123 ? (n132 ? !n122 : (n257 ? !n122 : 1'b0)) : (n132 ? 1'b1 : n257));
assign n6014 = /* LUT    1  9  2 */ (n75 ? n70 : (n67 ? n70 : (n70 ? n55 : 1'b0)));
assign n6015 = /* LUT   20  5  2 */ (n2784 ? !n2673 : n2673);
assign n6016 = /* LUT    9 11  2 */ (n587 ? !n564 : (n564 ? 1'b0 : !n698));
assign n6017 = /* LUT   12 19  3 */ (n1825 ? (n1646 ? !n5 : (n5 ? 1'b0 : n1821)) : (n1646 ? 1'b0 : (n5 ? 1'b0 : n1821)));
assign n6018 = /* LUT   18 10  0 */ (n2518 ? (n2500 ? (n2516 ? !n2509 : 1'b0) : 1'b1) : (n2500 ? (n2516 ? !n2509 : 1'b0) : n2509));
assign n6019 = /* LUT   13 15  1 */ (n1971 ? (n1969 ? n1787 : !n1787) : (n1969 ? !n1787 : n1787));
assign n6020 = /* LUT    7  3  5 */ n188;
assign n6021 = /* LUT   10 11  6 */ (n1311 ? (n1305 ? 1'b0 : !n1317) : 1'b0);
assign n6022 = /* LUT   13 18  6 */ (n1983 ? (n1780 ? (n1809 ? n5 : 1'b1) : (n1809 ? 1'b1 : n5)) : (n1780 ? (n1809 ? 1'b0 : !n5) : (n1809 ? !n5 : 1'b0)));
assign n6023 = /* LUT   10  8  0 */ (n1286 ? 1'b0 : (n1288 ? (n1285 ? n1118 : 1'b1) : 1'b0));
assign n6024 = /* LUT   21 21  6 */ (n2426 ? (n2292 ? (n2022 ? 1'b0 : !n2427) : 1'b0) : 1'b0);
assign n6025 = /* LUT    4 17  1 */ (n315 ? (n456 ? 1'b0 : n316) : 1'b0);
assign n6026 = /* LUT   11 16  1 */ (n1508 ? (n1459 ? n1268 : 1'b0) : n1459);
assign n6027 = /* LUT   13 10  7 */ n1454;
assign n6028 = /* LUT    2  9  4 */ (n68 ? !n106 : 1'b0);
assign n6029 = /* LUT   13  2  3 */ n179;
assign n6030 = /* LUT    3 13  6 */ n590;
assign n6031 = /* LUT    3  5  2 */ (n210 ? 1'b0 : (n204 ? (n200 ? 1'b1 : n206) : n200));
assign n6032 = /* LUT   14 23  6 */ (n2166 ? (n8 ? n1665 : !n1665) : (n8 ? !n1665 : n1665));
assign n6033 = /* LUT   15 19  4 */ n2289;
assign n6034 = /* LUT   15 11  0 */ (n2224 ? (n1473 ? 1'b1 : !n2237) : (n1473 ? n2237 : 1'b0));
assign n6035 = /* LUT   10  3  6 */ (n5 ? (n1410 ? 1'b0 : !n956) : (n1247 ? (n1410 ? 1'b0 : !n956) : !n956));
assign n6036 = /* LUT   12  7  6 */ n188;
assign n6037 = /* LUT   14 20  0 */ n1834;
assign n6038 = /* LUT   22  9  4 */ n2618;
assign n6039 = /* LUT   13  3  4 */ (n1595 ? (n1543 ? 1'b1 : !n1866) : (n1543 ? 1'b0 : !n1866));
assign n6040 = /* LUT   21 13  7 */ (n2820 ? (n8 ? n2824 : !n2824) : (n8 ? !n2824 : n2824));
assign n6041 = /* LUT    3  6  3 */ n177;
assign n6042 = /* LUT   21  5  3 */ (n2932 ? (n8 ? n2779 : !n2779) : (n8 ? !n2779 : n2779));
assign n6043 = /* LUT    4 21  7 */ (n802 ? !n334 : n334);
assign n6044 = /* LUT   11  8  2 */ (n5 ? (n1146 ? n984 : (n1579 ? n984 : 1'b0)) : n984);
assign n6045 = /* LUT   15 20  5 */ (n1491 ? 1'b0 : (n2021 ? !n1998 : 1'b0));
assign n6046 = /* LUT   15 12  1 */ (n2238 ? (n2117 ? n1632 : 1'b1) : (n2117 ? n1632 : !n1593));
assign n6047 = /* LUT   23 14  0 */ (n3032 ? !n3020 : (n2965 ? !n3020 : (n3020 ? 1'b0 : n3018)));
assign n6050 = /* LUT   22 10  5 */ (n2950 ? (n2951 ? 1'b0 : (n2952 ? n2953 : 1'b0)) : 1'b0);
assign n6051 = /* LUT    2 10  4 */ (n253 ? (n93 ? (n77 ? !n86 : 1'b1) : !n77) : !n77);
assign n6052 = /* LUT   22  2  1 */ (n2757 ? !io_19_0_1 : (n2889 ? 1'b0 : n3009));
assign n6053 = /* LUT    2  2  0 */ (n170 ? (n176 ? (n6 ? 1'b1 : n174) : !n6) : (n176 ? (n6 ? 1'b0 : n174) : !n6));
assign n6054 = /* LUT   21  6  4 */ n2607;
assign n6055 = /* LUT    8 13  0 */ n354;
assign n6056 = /* LUT   11  4  4 */ n179;
assign n6057 = /* LUT   22  3  2 */ (n3012 ? (n2889 ? !n2756 : n2896) : (n2889 ? !n2756 : !n2896));
assign n6058 = /* LUT   17 15  4 */ n2277;
assign n6061 = /* LUT   22  6  7 */ n2195;
assign n6062 = /* LUT   15  7  7 */ (n2056 ? 1'b0 : (n2057 ? 1'b0 : (n2061 ? 1'b0 : !n2059)));
assign n6063 = /* LUT    9 21  1 */ (n1233 ? n1226 : (n1223 ? n1226 : (n1226 ? 1'b1 : n1064)));
assign n6066 = /* LUT   14  8  3 */ (n1889 ? (n2070 ? 1'b0 : (n1750 ? 1'b1 : n1903)) : (n2070 ? 1'b0 : (n1750 ? n1903 : 1'b1)));
assign n6067 = /* LUT    8  9  2 */ (n1147 ? !n878 : n878);
assign n6068 = /* LUT   23 11  3 */ !n2500;
assign n6069 = /* LUT   20 23  4 */ n2012;
assign n6070 = /* LUT   17  8  1 */ n1965;
assign n6071 = /* LUT    9 22  2 */ (n1392 ? !n1189 : n1189);
assign n6072 = /* LUT   17 11  6 */ (n2367 ? (n2355 ? 1'b0 : (n2240 ? 1'b1 : n2364)) : (n2355 ? 1'b0 : (n2240 ? !n2364 : 1'b0)));
assign n6073 = /* LUT    4  6  4 */ (n402 ? (n545 ? 1'b0 : (n691 ? n694 : 1'b0)) : (n691 ? n694 : 1'b0));
assign n6074 = /* LUT    8 10  3 */ (n698 ? (n711 ? 1'b0 : (n761 ? !n564 : 1'b0)) : (n711 ? 1'b0 : !n564));
assign n6075 = /* LUT   14  1  0 */ (n1670 ? n5 : 1'b0);
assign n6076 = /* LUT   16 20  6 */ (n2297 ? (n2156 ? 1'b0 : (n2293 ? 1'b0 : n2298)) : 1'b0);
assign n6077 = /* LUT    1 20  1 */ (n149 ? !n146 : n146);
assign n6078 = /* LUT   16 12  2 */ (n2237 ? 1'b0 : !n2122);
assign n6079 = /* LUT   14  4  5 */ (n1179 ? n1410 : 1'b0);
assign n6080 = /* LUT   10 19  0 */ n1516;
assign n6081 = /* LUT    1 19  5 */ (n135 ? (n136 ? n141 : 1'b0) : 1'b0);
assign n6082 = /* LUT    5  3  2 */ (n383 ? (n212 ? 1'b0 : (n669 ? n519 : 1'b1)) : !n212);
assign n6083 = /* LUT   23  3  4 */ (n3049 ? (n2887 ? n8 : !n8) : (n2887 ? !n8 : n8));
assign n6084 = /* LUT   17  4  3 */ n2172;
assign n6085 = /* LUT    5  6  7 */ (n176 ? 1'b0 : (n6 ? 1'b1 : (n398 ? n41 : 1'b1)));
assign n6086 = /* LUT   16 13  3 */ n1755;
assign n6087 = /* LUT    4  2  6 */ (n664 ? (n361 ? (n661 ? n62 : 1'b0) : n62) : n62);
assign n6088 = /* LUT   14  5  6 */ n179;
assign n6089 = /* LUT    1 12  2 */ (n261 ? (io_4_31_0 ? 1'b0 : !n246) : 1'b0);
assign n6090 = /* LUT   13 21  7 */ (n1981 ? !n1652 : 1'b0);
assign n6091 = /* LUT   20  8  2 */ n2805;
assign n6092 = /* LUT   12 22  3 */ (n1851 ? !n1845 : n1845);
assign n6093 = /* LUT   20 11  7 */ (n2517 ? (n2705 ? 1'b0 : (n2704 ? !n2695 : 1'b1)) : (n2704 ? !n2695 : 1'b1));
assign n6094 = /* LUT   10 14  6 */ (n1459 ? 1'b0 : !n1360);
assign n6095 = /* LUT   10  6  2 */ (n1115 ? !n852 : 1'b0);
assign n6096 = /* LUT    9 10  5 */ (n1146 ? (n989 ? n811 : 1'b1) : 1'b0);
assign n6097 = /* LUT    9  2  1 */ (n1238 ? (n176 ? n1234 : 1'b0) : 1'b0);
assign n6098 = /* LUT   22 20  4 */ (n2855 ? (n2156 ? 1'b0 : (n2297 ? n2293 : 1'b0)) : 1'b0);
assign n6099 = /* LUT    3 16  1 */ (n80 ? (n303 ? (n592 ? !n446 : 1'b0) : 1'b0) : (n592 ? n446 : 1'b0));
assign n6100 = /* LUT   21 16  3 */ (n2404 ? n2846 : (n2846 ? !n2854 : !n2839));
assign n6101 = /* LUT   12 15  0 */ n1181;
assign n6102 = /* LUT   20  4  4 */ (n2673 ? 1'b0 : (n2675 ? (n2674 ? n7 : 1'b0) : 1'b0));
assign n6103 = /* LUT   10 15  7 */ (n1275 ? (n1356 ? 1'b0 : n1365) : (n1356 ? (n1365 ? !n1353 : 1'b0) : n1365));
assign n6104 = /* LUT   10  7  3 */ (n1272 ? (n858 ? (n1273 ? 1'b0 : n1277) : n1277) : (n1273 ? 1'b0 : n1277));
assign n6105 = /* LUT   18 17  6 */ (n2558 ? (n2403 ? !n2406 : (n2406 ? 1'b0 : !n2564)) : (n2403 ? 1'b0 : (n2406 ? 1'b0 : !n2564)));
assign n6106 = /* LUT   18  9  2 */ (n2364 ? (n2355 ? n2496 : n2501) : 1'b0);
assign n6107 = /* LUT    3  8  2 */ (n555 ? !n226 : n226);
assign n6108 = /* LUT   18 10  3 */ (n2631 ? (n2480 ? n2355 : (n2355 ? !n2364 : 1'b0)) : (n2480 ? (n2355 ? n2364 : 1'b0) : 1'b0));
assign n6109 = /* LUT    9  3  1 */ (n176 ? (n1258 ? n1254 : 1'b0) : 1'b0);
assign n6110 = /* LUT   15 22  4 */ n2012;
assign n6111 = /* LUT    3 11  7 */ (n264 ? 1'b0 : !n260);
assign n6112 = /* LUT   15 14  0 */ (n2246 ? (n1494 ? n1329 : 1'b0) : (n1494 ? n1329 : (n2117 ? n1329 : 1'b1)));
assign n6113 = /* LUT   21 17  3 */ (n2408 ? 1'b0 : (n2850 ? !n2406 : (n2406 ? !n2851 : 1'b1)));
assign n6114 = /* LUT    2 13  5 */ (n274 ? (n113 ? !n271 : n271) : 1'b0);
assign n6115 = /* LUT   12  2  2 */ !n852;
assign n6116 = /* LUT   13  6  4 */ (n1561 ? 1'b0 : (n1709 ? (n1712 ? 1'b0 : !n1707) : 1'b0));
assign n6117 = /* LUT    4 16  3 */ (n249 ? (n128 ? (n606 ? !n608 : 1'b0) : (n606 ? 1'b1 : n608)) : 1'b0);
assign n6118 = /* LUT   11 11  2 */ n1602;
assign n6119 = /* LUT   14 19  3 */ (n2149 ? (n2008 ? n1983 : !n1983) : (n2008 ? !n1983 : n1983));
assign n6120 = /* LUT   22  8  7 */ (n2937 ? (n2803 ? 1'b1 : n2801) : 1'b1);
assign n6123 = /* LUT    3  4  4 */ (n368 ? (n200 ? (n197 ? 1'b0 : !n176) : 1'b0) : (n200 ? !n176 : 1'b0));
assign n6124 = /* LUT   21  4  6 */ (n2922 ? (n2774 ? n8 : !n8) : (n2774 ? !n8 : n8));
assign n6125 = /* LUT   15 18  6 */ n2283;
assign n6128 = /* LUT   22  5  1 */ !n2778;
assign n6129 = /* LUT    5 13  1 */ !n581;
assign n6130 = /* LUT    4 17  4 */ (n159 ? 1'b0 : (n158 ? 1'b0 : !n292));
assign n6131 = /* LUT   21  1  0 */ (n2314 ? (n2448 ? (n2447 ? 1'b0 : !n2595) : 1'b0) : 1'b0);
assign n6132 = /* LUT    2  9  7 */ (n68 ? (n235 ? 1'b1 : n106) : n106);
assign n6133 = /* LUT   13  2  6 */ (n1668 ? n1550 : 1'b0);
assign n6137 = /* LUT   11  7  4 */ (n1146 ? n984 : (n1576 ? n984 : (n984 ? !n5 : 1'b0)));
assign n6138 = /* LUT    8 20  7 */ (n1031 ? 1'b0 : !n466);
assign n6139 = /* LUT   15 11  3 */ (n1728 ? (n2238 ? (n2095 ? n2103 : 1'b0) : n2103) : (n2095 ? n2103 : 1'b0));
assign n6140 = /* LUT   14 20  3 */ n1832;
assign n6141 = /* LUT   15 10  7 */ (n2090 ? (n1882 ? !n2062 : (n1714 ? !n2062 : 1'b0)) : (n1882 ? !n2062 : (n1714 ? 1'b0 : !n2062)));
assign n6142 = /* LUT   22  9  7 */ n2619;
assign n6143 = /* LUT   21  5  6 */ (n2935 ? (n2782 ? n8 : !n8) : (n2782 ? !n8 : n8));
assign n6144 = /* LUT    5  5  2 */ n175;
assign n6145 = /* LUT    4  1  1 */ (n651 ? 1'b0 : (n200 ? 1'b0 : !n502));
assign n6146 = /* LUT    8 12  2 */ n175;
assign n6147 = /* LUT   16 15  3 */ n1366;
assign n6148 = /* LUT   20 18  0 */ (n2739 ? (n2729 ? 1'b0 : !n2405) : (n2729 ? n2405 : 1'b1));
assign n6149 = /* LUT   15  3  4 */ n15;
assign n6150 = /* LUT   17 14  6 */ (n2549 ? !n2393 : n2393);
assign n6151 = /* LUT    7 17  5 */ (n448 ? (n769 ? (n605 ? 1'b1 : n5) : n5) : 1'b1);
assign n6152 = /* LUT    7  9  1 */ (n875 ? (n996 ? n8 : !n8) : (n996 ? !n8 : n8));
assign n6153 = /* LUT    2  1  7 */ n15;
assign n6154 = /* LUT    8 13  3 */ n179;
assign n6155 = /* LUT    4  5  7 */ n179;
assign n6156 = /* LUT   20 19  1 */ (n2407 ? (n2743 ? !n2734 : 1'b0) : n2741);
assign n6157 = /* LUT   14  7  5 */ (n1909 ? (n1410 ? (n1889 ? 1'b0 : !n956) : !n956) : (n1410 ? !n1889 : 1'b1));
assign n6158 = /* LUT   17 15  7 */ (n1 ? 1'b0 : n2272);
assign n6159 = /* LUT   17  7  3 */ n2486;
assign n6160 = /* LUT    9 21  4 */ (n1064 ? (n1225 ? !n1224 : (n1224 ? 1'b0 : n1232)) : !n1224);
assign n6161 = /* LUT   14  8  6 */ (n1932 ? 1'b0 : (n1909 ? !n1925 : n1925));
assign n6162 = /* LUT    1 15  2 */ (n5 ? 1'b0 : (n108 ? 1'b0 : io_4_31_0));
assign n6163 = /* LUT   13 16  3 */ (n1984 ? !n852 : n852);
assign n6164 = /* LUT    3 19  2 */ (n632 ? !n477 : n477);
assign n6167 = /* LUT   20 14  7 */ (n2818 ? (n2834 ? !n2824 : 1'b0) : (n2822 ? 1'b0 : !n2824));
assign n6168 = /* LUT   10  9  2 */ (n1450 ? n1285 : (n1299 ? (n1285 ? !n720 : 1'b0) : 1'b0));
assign n6169 = /* LUT    9 13  5 */ (n1175 ? (n620 ? 1'b1 : !n679) : (n620 ? (n1187 ? 1'b1 : n679) : (n1187 ? !n679 : 1'b0)));
assign n6170 = /* LUT    9  5  1 */ (n807 ? !n852 : 1'b0);
assign n6171 = /* LUT   13 17  4 */ n1989;
assign n6172 = /* LUT   16  4  1 */ (n2177 ? 1'b1 : n2175);
assign n6173 = /* LUT    8  1  6 */ (n41 ? 1'b1 : (n938 ? (n933 ? 1'b0 : !n6) : (n933 ? n6 : 1'b1)));
assign n6174 = /* LUT   21 19  3 */ (n2427 ? 1'b0 : (n2292 ? (n2022 ? 1'b0 : !n2426) : 1'b0));
assign n6175 = /* LUT   12 18  0 */ n1641;
assign n6176 = /* LUT   20  7  4 */ n2796;
assign n6177 = /* LUT   10 10  3 */ (n1288 ? (n1010 ? !n1455 : (n1298 ? 1'b0 : !n1455)) : 1'b0);
assign n6178 = /* LUT   12 21  5 */ (n189 ? n1523 : 1'b0);
assign n6179 = /* LUT   18 12  2 */ n2626;
assign n6180 = /* LUT    9  6  2 */ (n1125 ? 1'b0 : n1126);
assign n6181 = /* LUT    2 16  0 */ (n80 ? (n294 ? 1'b0 : (n452 ? n293 : 1'b0)) : 1'b0);
assign n6182 = /* LUT   21 20  4 */ (n2404 ? n2996 : n2866);
assign n6183 = /* LUT    9  9  7 */ (n1292 ? (n488 ? !n1136 : (n679 ? 1'b0 : !n1136)) : (n488 ? 1'b1 : !n679));
assign n6184 = /* LUT   21 12  0 */ (n2509 ? (n2956 ? (n2513 ? !n2809 : 1'b0) : 1'b0) : (n2513 ? n2809 : 1'b0));
assign n6185 = /* LUT    1  4  1 */ (n38 ? (n33 ? (n16 ? n25 : 1'b0) : (n16 ? !n25 : 1'b0)) : (n33 ? (n16 ? 1'b0 : n25) : (n16 ? 1'b0 : !n25)));
assign n6186 = /* LUT   20  8  5 */ (n1 ? 1'b0 : n2693);
assign n6187 = /* LUT   18 13  3 */ n2654;
assign n6188 = /* LUT    1  3  5 */ (n35 ? (n14 ? (n18 ? n40 : 1'b0) : (n18 ? !n40 : 1'b0)) : (n14 ? (n18 ? 1'b0 : n40) : (n18 ? 1'b0 : !n40)));
assign n6189 = /* LUT   12 14  2 */ (n1793 ? (n1618 ? 1'b0 : n1623) : (n1618 ? n1623 : 1'b0));
assign n6190 = /* LUT   12 13  6 */ (n1615 ? (n1349 ? 1'b0 : (n1777 ? 1'b1 : !n1783)) : (n1349 ? 1'b0 : (n1777 ? n1783 : 1'b0)));
assign n6191 = /* LUT   22 20  7 */ (n2156 ? 1'b0 : (n2293 ? (n2992 ? n2297 : 1'b0) : 1'b0));
assign n6199 = /* LUT   14 22  3 */ !n2006;
assign n6203 = /* LUT    2 11  6 */ (n260 ? 1'b0 : !n259);
assign n6204 = /* LUT    3  7  4 */ (n410 ? (n542 ? n41 : (n41 ? n6 : 1'b0)) : (n542 ? (n41 ? !n6 : 1'b0) : 1'b0));
assign n6205 = /* LUT   11 10  5 */ (n1462 ? (n1468 ? (n1307 ? 1'b1 : n1448) : 1'b1) : 1'b0);
assign n6206 = /* LUT   18  9  5 */ n1965;
assign n6207 = /* LUT   12  6  3 */ (n1410 ? (n1702 ? 1'b0 : (n1418 ? !n956 : 1'b1)) : (n1418 ? !n956 : 1'b1));
assign n6208 = /* LUT   15 13  2 */ (n2104 ? 1'b0 : !n2102);
assign n6209 = /* LUT    4 20  4 */ (n628 ? !n641 : (n470 ? n627 : 1'b1));
assign n6213 = /* LUT    2 12  7 */ (n264 ? 1'b0 : (n212 ? (n422 ? 1'b0 : n426) : n426));
assign n6214 = /* LUT   13  5  6 */ (n1893 ? (n1687 ? 1'b1 : n1249) : (n1687 ? !n1249 : 1'b0));
assign n6215 = /* LUT   14 15  0 */ (n1966 ? !n1541 : n1541);
assign n6216 = /* LUT    2  4  3 */ (n37 ? !n193 : n193);
assign n6217 = /* LUT    3  8  5 */ (n43 ? (n83 ? n403 : 1'b0) : (n83 ? n238 : 1'b0));
assign n6218 = /* LUT   21  8  7 */ (n2940 ? (n2804 ? n2687 : !n2687) : (n2804 ? !n2799 : n2799));
assign n6219 = /* LUT   22  4  4 */ !n2771;
assign n6220 = /* LUT   14 18  5 */ (n1992 ? 1'b0 : (n1993 ? 1'b0 : (n1987 ? 1'b0 : !n1995)));
assign n6221 = /* LUT   11  2  0 */ (n1536 ? 1'b0 : (n960 ? !n1539 : 1'b1));
assign n6222 = /* LUT   15 14  3 */ (n2116 ? (n1624 ? !n2122 : 1'b1) : 1'b0);
assign n6225 = /* LUT    4 16  6 */ (n129 ? (n452 ? 1'b1 : n434) : 1'b0);
assign n6226 = /* LUT   11 11  5 */ (n1471 ? 1'b0 : (n277 ? n1268 : 1'b1));
assign n6227 = /* LUT   11  3  1 */ n188;
assign n6228 = /* LUT   14 11  2 */ (n2102 ? (n1940 ? (n2097 ? n1749 : 1'b0) : n1749) : (n1940 ? n2097 : 1'b1));
assign n6229 = /* LUT    8 11  5 */ (n1011 ? (n882 ? 1'b1 : (n1016 ? 1'b0 : n1012)) : 1'b0);
assign n6232 = /* LUT    7 12  1 */ n730;
assign n6233 = /* LUT    5  4  4 */ (n357 ? (n41 ? (n506 ? !n6 : 1'b1) : n6) : (n41 ? (n506 ? !n6 : 1'b1) : 1'b1));
assign n6234 = /* LUT    4  8  7 */ (n549 ? (n553 ? n52 : 1'b0) : (n553 ? (n44 ? n52 : !n52) : 1'b0));
assign n6235 = /* LUT   16 11  0 */ (n2239 ? (n2232 ? 1'b1 : n2220) : !n1705);
assign n6236 = /* LUT   16 14  5 */ (n1624 ? n2129 : (n2129 ? (n1790 ? !n2252 : 1'b1) : 1'b0));
assign n6237 = /* LUT   17 18  7 */ !n2415;
assign n6238 = /* LUT   17 10  3 */ n1754;
assign n6239 = /* LUT    7 13  2 */ (n887 ? (n564 ? 1'b1 : n711) : n711);
assign n6240 = /* LUT   15  2  6 */ (n1701 ? (n1549 ? 1'b0 : !n1543) : !n1549);
assign n6241 = /* LUT    5  5  5 */ (n41 ? (n382 ? (n6 ? !n221 : 1'b0) : (n6 ? !n221 : 1'b1)) : 1'b1);
assign n6245 = /* LUT    7 16  7 */ !n488;
assign n6246 = /* LUT    4  1  4 */ n233;
assign n6247 = /* LUT   14  3  2 */ n177;
assign n6248 = /* LUT    8  4  1 */ (n974 ? (n944 ? 1'b1 : (n841 ? n5 : 1'b1)) : (n944 ? n841 : (n841 ? n5 : 1'b0)));
assign n6249 = /* LUT   16 15  6 */ n1482;
assign n6250 = /* LUT   16  7  2 */ n1789;
assign n6251 = /* LUT   13 19  3 */ (n2002 ? !n1649 : n1649);
assign n6252 = /* LUT   20 18  3 */ (n2721 ? (n2581 ? 1'b0 : (n2404 ? 1'b0 : n2403)) : (n2581 ? (n2404 ? n2403 : 1'b0) : n2403));
assign n6253 = /* LUT   17  3  0 */ (n2304 ? (n2321 ? !n2182 : 1'b0) : n2321);
assign n6254 = /* LUT   23  5  6 */ n2457;
assign n6255 = /* LUT    1 14  5 */ (n110 ? n281 : 1'b0);
assign n6258 = /* LUT   10 20  6 */ (n177 ? (n1379 ? (n175 ? n189 : 1'b0) : 1'b0) : 1'b0);
assign n6259 = /* LUT    9  8  1 */ (n573 ? (n711 ? 1'b0 : n811) : (n5 ? n811 : (n711 ? 1'b0 : n811)));
assign n6260 = /* LUT   13 20  4 */ (n2015 ? (n1715 ? n8 : !n8) : (n1715 ? !n8 : n8));
assign n6261 = /* LUT   13 12  0 */ (n1772 ? (n1494 ? 1'b0 : !n1751) : !n1494);
assign n6262 = /* LUT    3 18  4 */ (n301 ? n132 : 1'b0);
assign n6263 = /* LUT   20  2  0 */ (n2333 ? (n2449 ? !n2313 : 1'b0) : n2449);
assign n6264 = /* LUT   12 16  1 */ (n1783 ? (n1349 ? 1'b0 : n1799) : (n1204 ? !n1349 : 1'b0));
assign n6265 = /* LUT   22 19  1 */ n2012;
assign n6269 = /* LUT    7  1  5 */ (n5 ? n679 : (n515 ? (n825 ? n679 : 1'b1) : (n825 ? 1'b0 : !n679)));
assign n6270 = /* LUT   13 13  1 */ n1760;
assign n6271 = /* LUT    9 12  7 */ (n1179 ? n362 : 1'b0);
assign n6272 = /* LUT   21 15  0 */ (n2818 ? 1'b0 : (n2824 ? (n2820 ? 1'b0 : n2821) : 1'b0));
assign n6273 = /* LUT    1  7  1 */ (n228 ? (n63 ? n49 : !n49) : (n63 ? !n49 : n49));
assign n6274 = /* LUT   13 16  6 */ (n212 ? (n1982 ? n1125 : !n1125) : (n1982 ? !n1125 : n1125));
assign n6275 = /* LUT   20  3  1 */ n2454;
assign n6276 = /* LUT   11 21  4 */ (n5 ? 1'b0 : (n80 ? (n1519 ? !n1525 : 1'b0) : 1'b1));
assign n6277 = /* LUT   12 17  2 */ (n1485 ? (n1638 ? 1'b1 : (n1652 ? 1'b1 : n1483)) : (n1652 ? 1'b1 : n1483));
assign n6278 = /* LUT   20  6  6 */ (n2789 ? !n2682 : n2682);
assign n6279 = /* LUT   10  9  5 */ (n1000 ? n1146 : (n811 ? n1146 : 1'b0));
assign n6280 = /* LUT   18 11  4 */ n2641;
assign n6281 = /* LUT    9  5  4 */ (n679 ? 1'b0 : (n5 ? !n806 : (n968 ? !n806 : 1'b1)));
assign n6282 = /* LUT   11 14  1 */ (n1181 ? 1'b0 : (n1460 ? 1'b1 : n1611));
assign n6283 = /* LUT    2 14  6 */ (n268 ? (n281 ? 1'b1 : n103) : 1'b0);
assign n6284 = /* LUT   13  8  7 */ (n1301 ? 1'b0 : (n1750 ? !n1579 : n1579));
assign n6285 = /* LUT   11 13  5 */ (n1334 ? 1'b0 : (n1599 ? !n1337 : 1'b0));
assign n6286 = /* LUT   18 12  5 */ n2645;
assign n6287 = /* LUT   18  4  1 */ n2321;
assign n6288 = /* LUT    5 19  1 */ (n822 ? 1'b0 : (n80 ? (n303 ? !n280 : 1'b0) : 1'b0));
assign n6289 = /* LUT   10  1  6 */ (n1235 ? (n6 ? n41 : (n1241 ? !n41 : 1'b1)) : (n6 ? 1'b1 : (n1241 ? !n41 : 1'b1)));
assign n6290 = /* LUT   24 15  1 */ n2012;
assign n6291 = /* LUT    4 15  0 */ (n446 ? 1'b0 : (n303 ? 1'b0 : (n87 ? 1'b0 : !n752)));
assign n6292 = /* LUT    2 15  7 */ (n290 ? 1'b0 : (n422 ? (n212 ? 1'b0 : !n264) : !n264));
assign n6293 = /* LUT   12  4  4 */ (n1249 ? (n1542 ? 1'b0 : n1546) : (n1686 ? 1'b0 : n1546));
assign n6294 = /* LUT   22  7  4 */ (n2794 ? 1'b0 : (n2939 ? !n2790 : 1'b0));
assign n6295 = /* LUT    2  7  3 */ (n51 ? (n52 ? 1'b0 : n372) : (n52 ? n232 : 1'b0));
assign n6296 = /* LUT    3  3  1 */ n15;
assign n6297 = /* LUT   21  3  3 */ (n2904 ? (n8 ? n2763 : !n2763) : (n8 ? !n2763 : n2763));
assign n6298 = /* LUT   14 21  5 */ (n5 ? 1'b0 : n1491);
assign n6299 = /* LUT   11  6  2 */ (n1416 ? 1'b0 : !n1541);
assign n6300 = /* LUT    5 20  2 */ (n648 ? (n627 ? (n619 ? !n620 : n620) : 1'b0) : 1'b0);
assign n6301 = /* LUT   17 21  3 */ n2012;
assign n6302 = /* LUT   11  9  7 */ (n1446 ? (n1295 ? 1'b1 : !n1449) : 1'b0);
assign n6303 = /* LUT   12  5  5 */ n179;
assign n6304 = /* LUT    2  8  4 */ (n413 ? (n240 ? !n230 : 1'b0) : (n240 ? n230 : 1'b0));
assign n6307 = /* LUT    4 19  6 */ (n464 ? 1'b0 : !n249);
assign n6308 = /* LUT   14 22  6 */ (n1846 ? (n8 ? n2018 : !n2018) : (n8 ? !n2018 : n2018));
assign n6309 = /* LUT   14 14  2 */ (n1494 ? n1961 : (n1947 ? n1772 : (n1961 ? 1'b0 : !n1772)));
assign n6310 = /* LUT   15 10  0 */ n1757;
assign n6311 = /* LUT    8 14  5 */ (n1050 ? (n1023 ? (n1025 ? n1189 : 1'b0) : (n1025 ? !n1189 : 1'b0)) : (n1023 ? (n1025 ? 1'b0 : n1189) : (n1025 ? 1'b0 : !n1189)));
assign n6312 = /* LUT   15 13  5 */ (n2117 ? !n2115 : (n2122 ? 1'b1 : (n2115 ? !n2242 : 1'b1)));
assign n6313 = /* LUT   23 16  6 */ n2012;
assign n6316 = /* LUT    5  7  4 */ n15;
assign n6317 = /* LUT    9 19  1 */ (n1378 ? !n1212 : 1'b0);
assign n6318 = /* LUT    4 11  7 */ (n446 ? 1'b0 : (n62 ? 1'b0 : (n87 ? 1'b0 : !n452)));
assign n6319 = /* LUT   23 13  0 */ (n2713 ? 1'b1 : n2959);
assign n6320 = /* LUT   11  2  3 */ (n41 ? (n966 ? n6 : 1'b1) : (n1253 ? 1'b0 : !n6));
assign n6321 = /* LUT    4  3  3 */ (n176 ? (n668 ? n505 : 1'b0) : 1'b0);
assign n6326 = /* LUT   16 17  5 */ (n1823 ? 1'b1 : !n2271);
assign n6327 = /* LUT   17 13  3 */ (n2538 ? !n2387 : n2387);
assign n6328 = /* LUT   20 13  0 */ (n2814 ? n2543 : 1'b0);
assign n6329 = /* LUT   15  5  6 */ n179;
assign n6330 = /* LUT    5  8  5 */ (n722 ? (n558 ? 1'b0 : n704) : (n558 ? (n704 ? n709 : 1'b0) : n704));
assign n6331 = /* LUT    7 19  7 */ (n490 ? 1'b0 : !n488);
assign n6332 = /* LUT   16 18  6 */ n2418;
assign n6333 = /* LUT   16 10  2 */ (n1756 ? (n2364 ? (n2355 ? 1'b0 : !n2090) : 1'b0) : (n2364 ? (n2355 ? 1'b0 : !n2090) : !n2355));
assign n6337 = /* LUT   14  2  5 */ (n1863 ? (n1883 ? 1'b0 : (n1550 ? !n212 : 1'b1)) : (n1550 ? !n212 : 1'b1));
assign n6340 = /* LUT    1 17  5 */ (n134 ? 1'b0 : (n306 ? 1'b0 : (n288 ? n113 : 1'b1)));
assign n6341 = /* LUT   17  9  5 */ (n2364 ? (n2355 ? !n2372 : 1'b0) : (n2354 ? 1'b0 : n2355));
assign n6342 = /* LUT    7 12  4 */ n583;
assign n6343 = /* LUT    7  4  0 */ (n967 ? (n861 ? n958 : 1'b0) : 1'b0);
assign n6347 = /* LUT   10 11  5 */ (n483 ? (n212 ? !n1268 : (n261 ? !n1268 : 1'b0)) : (n261 ? !n1268 : 1'b0));
assign n6348 = /* LUT   13 18  5 */ (n1648 ? 1'b0 : (n1553 ? 1'b0 : (n1649 ? 1'b0 : !n1715)));
assign n6349 = /* LUT    3 21  4 */ (n483 ? 1'b0 : (n486 ? n5 : 1'b1));
assign n6350 = /* LUT    1 13  7 */ (n110 ? (n273 ? n263 : 1'b0) : n263);
assign n6351 = /* LUT   20  9  7 */ n2067;
assign n6352 = /* LUT   21 18  0 */ n2012;
assign n6353 = /* LUT   13 19  6 */ (n2005 ? !n1647 : n1647);
assign n6354 = /* LUT   13 11  2 */ n1453;
assign n6355 = /* LUT   21 21  5 */ (n2404 ? n2872 : (n2872 ? (n2871 ? 1'b1 : n3001) : 1'b0));
assign n6358 = /* LUT   11 16  0 */ (n1369 ? 1'b0 : !n1459);
assign n6361 = /* LUT   10 12  5 */ (n1181 ? 1'b0 : (n1313 ? 1'b0 : n1470));
assign n6362 = /* LUT   10  4  1 */ (n5 ? 1'b0 : n956);
assign n6363 = /* LUT    9  8  4 */ (n1128 ? (n5 ? 1'b0 : !n1267) : !n1267);
assign n6364 = /* LUT   22 18  3 */ (n2156 ? 1'b0 : (n2297 ? (n2848 ? !n2293 : 1'b0) : 1'b0));
assign n6365 = /* LUT    2 18  2 */ (n301 ? n268 : (n139 ? n268 : 1'b0));
assign n6366 = /* LUT   21 14  2 */ (n2712 ? 1'b1 : n2816);
assign n6367 = /* LUT   13  3  3 */ (n1688 ? (n1422 ? n1429 : 1'b1) : (n1673 ? (n1422 ? n1429 : 1'b0) : (n1422 ? n1429 : 1'b1)));
assign n6368 = /* LUT    3  6  2 */ (n530 ? (n232 ? !n543 : 1'b0) : (n232 ? (n41 ? 1'b1 : !n543) : 1'b0));
assign n6369 = /* LUT   18 15  5 */ (n2432 ? (n2156 ? (n2297 ? !n2293 : 1'b0) : 1'b0) : 1'b0);
assign n6370 = /* LUT    3  9  7 */ (n69 ? 1'b1 : (n106 ? 1'b0 : n419));
assign n6371 = /* LUT   15 12  0 */ (n2241 ? (n2116 ? (n2117 ? n2106 : 1'b1) : 1'b0) : (n2116 ? (n2117 ? n2106 : !n2106) : 1'b0));
assign n6372 = /* LUT   17 23  2 */ (n2297 ? 1'b0 : (n2432 ? (n2156 ? 1'b0 : n2293) : 1'b0));
assign n6376 = /* LUT   22 10  4 */ (n2953 ? 1'b0 : (n2951 ? 1'b0 : n2066));
assign n6377 = /* LUT    2 10  3 */ (n250 ? (n253 ? (n80 ? 1'b0 : n246) : (n80 ? 1'b1 : n246)) : 1'b0);
assign n6378 = /* LUT    5 18  4 */ (n617 ? (n648 ? (n627 ? !n777 : 1'b0) : 1'b0) : (n648 ? (n627 ? n777 : 1'b0) : 1'b0));
assign n6379 = /* LUT   21  6  3 */ n2604;
assign n6380 = /* LUT   14 16  1 */ (n1956 ? (n1978 ? (n1980 ? n5 : 1'b1) : (n1980 ? 1'b1 : n5)) : (n1978 ? (n1980 ? 1'b0 : !n5) : (n1980 ? !n5 : 1'b0)));
assign n6381 = /* LUT    3  2  4 */ (n347 ? (n41 ? n6 : (n349 ? !n6 : 1'b1)) : (n41 ? 1'b1 : (n349 ? !n6 : 1'b1)));
assign n6382 = /* LUT   11 12  7 */ n1329;
assign n6383 = /* LUT   23 15  0 */ (n3032 ? 1'b1 : n2841);
assign n6384 = /* LUT   11  4  3 */ (n1126 ? 1'b0 : (n1541 ? (n1125 ? 1'b0 : !n1416) : 1'b0));
assign n6385 = /* LUT   12  8  5 */ (n1741 ? (n1271 ? !n1583 : (n1290 ? !n1583 : 1'b0)) : (n1271 ? (n1290 ? !n1583 : 1'b0) : !n1583));
assign n6386 = /* LUT   15 16  6 */ (n1491 ? (n1623 ? n2251 : 1'b1) : !n1623);
assign n6387 = /* LUT    2  3  0 */ n187;
assign n6388 = /* LUT    4 14  2 */ (n597 ? 1'b0 : (n598 ? 1'b0 : (n449 ? 1'b0 : !n443)));
assign n6389 = /* LUT    8 18  1 */ (n1208 ? (n212 ? 1'b0 : n1199) : 1'b0);
assign n6390 = /* LUT   21  2  5 */ (n2757 ? 1'b1 : n2756);
assign n6391 = /* LUT   11  5  4 */ (n1541 ? (n1539 ? (n1421 ? n1106 : 1'b0) : 1'b0) : 1'b0);
assign n6399 = /* LUT   12  4  7 */ (n1541 ? 1'b0 : n1416);
assign n6400 = /* LUT   15  8  7 */ (n1689 ? !n2068 : (n2068 ? 1'b0 : (n1887 ? n1929 : !n1929)));
assign n6401 = /* LUT   22  7  7 */ (n2804 ? 1'b0 : (n2691 ? 1'b0 : (n2690 ? 1'b0 : !n2692)));
assign n6402 = /* LUT    9 22  1 */ (n1019 ? !n1050 : n1050);
assign n6403 = /* LUT   21  3  6 */ (n2907 ? (n2766 ? n8 : !n8) : (n2766 ? !n8 : n8));
assign n6404 = /* LUT   16 21  1 */ (n1526 ? !n2022 : 1'b0);
assign n6405 = /* LUT    7 14  4 */ n304;
assign n6406 = /* LUT    8 10  2 */ (n852 ? 1'b0 : n1001);
assign n6410 = /* LUT    5  3  1 */ n175;
assign n6411 = /* LUT   17  4  2 */ n2311;
assign n6412 = /* LUT    5  6  6 */ (n564 ? 1'b0 : (n5 ? 1'b1 : (n698 ? n683 : 1'b1)));
assign n6413 = /* LUT    1 21  1 */ (n156 ? (n152 ? 1'b0 : n157) : (n152 ? n157 : 1'b0));
assign n6414 = /* LUT   16 13  2 */ n2067;
assign n6415 = /* LUT    4  2  5 */ n175;
assign n6416 = /* LUT   14  5  5 */ (n1126 ? (n1416 ? 1'b0 : (n1125 ? n1541 : 1'b0)) : 1'b0);
assign n6417 = /* LUT   16 16  7 */ (n2278 ? 1'b0 : n2125);
assign n6420 = /* LUT    7  7  0 */ (n869 ? !n864 : n864);
assign n6421 = /* LUT    5  7  7 */ (n690 ? (n710 ? (n702 ? !n689 : 1'b0) : n702) : (n702 ? !n689 : 1'b0));
assign n6422 = /* LUT    9 19  4 */ (n907 ? 1'b0 : (n1213 ? n1210 : 1'b0));
assign n6423 = /* LUT    4  3  6 */ n354;
assign n6424 = /* LUT   16  9  4 */ n1755;
assign n6425 = /* LUT   17  5  2 */ n2330;
assign n6426 = /* LUT    3 16  0 */ (n445 ? n287 : (n449 ? n287 : 1'b0));
assign n6427 = /* LUT   18 18  1 */ (n2404 ? (n2561 ? (n2403 ? 1'b1 : n2567) : (n2403 ? 1'b0 : n2567)) : 1'b0);
assign n6428 = /* LUT   20 12  7 */ n1755;
assign n6429 = /* LUT   10 15  6 */ n1268;
assign n6430 = /* LUT   10  7  2 */ (n841 ? (n1135 ? n1280 : 1'b0) : n1280);
assign n6431 = /* LUT   13 22  6 */ (n1859 ? (n1835 ? (n5 ? 1'b0 : n1663) : !n5) : (n1835 ? (n5 ? 1'b0 : n1663) : 1'b0));
assign n6432 = /* LUT   22 21  4 */ (n3041 ? (n2403 ? (n2406 ? !n3042 : 1'b0) : 1'b0) : (n2403 ? (n2406 ? !n3042 : 1'b0) : n2406));
assign n6433 = /* LUT    2 21  3 */ (n331 ? 1'b0 : n150);
assign n6434 = /* LUT   13 14  2 */ (n1790 ? 1'b0 : (n1957 ? !n1624 : 1'b0));
assign n6435 = /* LUT   22 13  0 */ (n2716 ? n2814 : 1'b0);
assign n6436 = /* LUT    3 17  1 */ (n465 ? !n614 : n614);
assign n6437 = /* LUT   16  1  5 */ io_16_0_0;
assign n6438 = /* LUT    9 11  4 */ (n1169 ? (n564 ? 1'b1 : n711) : n711);
assign n6439 = /* LUT   18 10  2 */ (n2505 ? (n2366 ? 1'b0 : n2362) : (n2506 ? (n2366 ? 1'b0 : n2362) : (n2366 ? 1'b1 : n2362)));
assign n6440 = /* LUT    9  3  0 */ n179;
assign n6441 = /* LUT   12 11  1 */ n1732;
assign n6442 = /* LUT    7  3  7 */ (n657 ? (n679 ? 1'b1 : (n5 ? 1'b0 : !n835)) : (n679 ? n5 : (n5 ? 1'b0 : !n835)));
assign n6443 = /* LUT   13 15  3 */ (n1975 ? (n1801 ? n1802 : !n1802) : (n1801 ? !n1802 : n1802));
assign n6444 = /* LUT   11 20  1 */ (n1520 ? 1'b0 : !n1380);
assign n6445 = /* LUT   10  8  2 */ (n1267 ? 1'b0 : (n812 ? 1'b1 : (n811 ? 1'b1 : !n5)));
assign n6446 = /* LUT    9  4  1 */ (n1104 ? (n1103 ? !n806 : 1'b0) : (n1103 ? !n806 : (n806 ? 1'b0 : n1112)));
assign n6447 = /* LUT   22 22  4 */ n2012;
assign n6451 = /* LUT   21 18  3 */ (n2746 ? (n2991 ? 1'b1 : (n2988 ? 1'b1 : !n2406)) : 1'b0);
assign n6452 = /* LUT    9  7  6 */ n177;
assign n6455 = /* LUT    5 13  0 */ (n128 ? (n455 ? n745 : 1'b0) : 1'b0);
assign n6456 = /* LUT    4 17  3 */ (n446 ? n268 : (n607 ? n268 : (n268 ? n291 : 1'b0)));
assign n6457 = /* LUT   11 16  3 */ (n1457 ? 1'b0 : n1497);
assign n6458 = /* LUT    2  9  6 */ (n241 ? (n226 ? n64 : !n64) : 1'b0);
assign n6459 = /* LUT   13  2  5 */ (n1550 ? n1669 : 1'b0);
assign n6460 = /* LUT    3  5  4 */ (n200 ? (n533 ? (n176 ? 1'b0 : !n534) : !n534) : 1'b0);
assign n6461 = /* LUT   11 15  7 */ (n1599 ? (n1481 ? 1'b1 : (n1436 ? 1'b1 : n1496)) : 1'b0);
assign n6462 = /* LUT   15 11  2 */ (n2237 ? !n1330 : n2227);
assign n6466 = /* LUT    5 14  1 */ (n249 ? (n753 ? !n756 : 1'b0) : !n756);
assign n6467 = /* LUT   14 20  2 */ n1833;
assign n6468 = /* LUT    8 21  1 */ (n1075 ? n926 : (n1064 ? (n926 ? 1'b1 : !n1222) : n926));
assign n6469 = /* LUT   13  3  6 */ (n1703 ? (n1716 ? (n1875 ? 1'b0 : !n1863) : !n1875) : (n1716 ? !n1863 : 1'b1));
assign n6470 = /* LUT   22  9  6 */ n2620;
assign n6471 = /* LUT   21  5  5 */ (n2934 ? (n8 ? !n2929 : n2929) : (n8 ? n2929 : !n2929));
assign n6472 = /* LUT   17 20  0 */ (n2580 ? (n2297 ? (n2022 ? n2413 : 1'b0) : (n2022 ? n2413 : 1'b1)) : (n2297 ? (n2022 ? n2413 : 1'b1) : (n2022 ? n2413 : 1'b0)));
assign n6473 = /* LUT   11  8  4 */ (n1575 ? !n212 : (n5 ? (n212 ? 1'b0 : n1146) : !n212));
assign n6474 = /* LUT   15 12  3 */ (n2117 ? 1'b0 : !n2104);
assign n6475 = /* LUT   23 14  2 */ (n3021 ? (n3025 ? n3020 : (n3020 ? 1'b1 : n2968)) : (n3025 ? n3020 : (n3020 ? 1'b1 : !n2968)));
assign n6478 = /* LUT    2 10  6 */ (n235 ? (n93 ? 1'b0 : !n254) : 1'b0);
assign n6479 = /* LUT   22  2  3 */ (n2890 ? 1'b0 : (n2891 ? 1'b0 : (n2893 ? n2895 : 1'b0)));
assign n6480 = /* LUT    2  2  2 */ (n165 ? (n172 ? 1'b1 : n176) : (n172 ? !n176 : 1'b0));
assign n6481 = /* LUT   21  6  6 */ n2605;
assign n6484 = /* LUT    8 13  2 */ n233;
assign n6485 = /* LUT    5  9  7 */ (n714 ? (n574 ? (n561 ? 1'b0 : n724) : n724) : (n561 ? 1'b0 : n724));
assign n6486 = /* LUT    4  5  6 */ (n6 ? 1'b1 : (n684 ? (n41 ? 1'b0 : !n683) : (n41 ? 1'b1 : !n683)));
assign n6487 = /* LUT   11  4  6 */ n15;
assign n6492 = /* LUT    7 10  1 */ (n5 ? (n711 ? (n811 ? !n567 : 1'b0) : n811) : (n711 ? 1'b0 : n811));
assign n6493 = /* LUT    9 21  3 */ (n924 ? 1'b0 : (n1069 ? !n1217 : (n1217 ? 1'b0 : n437)));
assign n6494 = /* LUT   20 20  1 */ (n2869 ? 1'b1 : (n2867 ? !n2408 : (n2750 ? !n2408 : 1'b0)));
assign n6495 = /* LUT   14  8  5 */ n2067;
assign n6496 = /* LUT    8  9  4 */ (n1149 ? !n989 : n989);
assign n6497 = /* LUT   11 30  0 */ (n1502 ? (n466 ? 1'b1 : n188) : (n466 ? 1'b1 : n5));
assign n6498 = /* LUT   17  8  3 */ n1754;
assign n6501 = /* LUT    9 22  4 */ (n1394 ? !n907 : n907);
assign n6502 = /* LUT   23  2  5 */ n3045;
assign n6503 = /* LUT    4  6  6 */ (n686 ? (n546 ? n51 : 1'b0) : (n546 ? (n693 ? n51 : !n51) : 1'b0));
assign n6504 = /* LUT   14  1  2 */ n15;
assign n6505 = /* LUT    8  2  1 */ (n943 ? n957 : (n957 ? (n200 ? 1'b1 : n949) : 1'b0));
assign n6506 = /* LUT   16 12  4 */ (n2384 ? (n1453 ? (n2238 ? n2237 : 1'b1) : (n2238 ? n2237 : 1'b0)) : (n1453 ? 1'b1 : n2238));
assign n6507 = /* LUT   16  4  0 */ (n2174 ? 1'b1 : n2176);
assign n6510 = /* LUT   14  4  7 */ (n1543 ? (n1863 ? (n1904 ? 1'b0 : !n1884) : !n1904) : (n1863 ? !n1884 : 1'b1));
assign n6511 = /* LUT   20 16  3 */ n2012;
assign n6512 = /* LUT    8  1  5 */ n179;
assign n6513 = /* LUT    1 19  7 */ (n150 ? !n141 : 1'b0);
assign n6514 = /* LUT   18 21  1 */ (n2404 ? !n2587 : (n2587 ? !n2159 : !n2585));
assign n6515 = /* LUT    1 11  3 */ (n75 ? 1'b1 : n260);
assign n6516 = /* LUT   20 15  7 */ (n2818 ? (n2840 ? 1'b0 : (n2715 ? 1'b1 : n2827)) : (n2840 ? 1'b1 : (n2715 ? 1'b1 : n2827)));
assign n6517 = /* LUT   17  4  5 */ n2318;
assign n6518 = /* LUT   10 10  2 */ (n811 ? n1146 : (n1146 ? !n880 : 1'b0));
assign n6519 = /* LUT    9  6  1 */ (n5 ? (n1123 ? 1'b0 : !n1267) : !n1267);
assign n6520 = /* LUT   16  5  1 */ (n2180 ? 1'b0 : (n2188 ? 1'b0 : (n2181 ? 1'b0 : !n1902)));
assign n6521 = /* LUT   10 13  7 */ (n1186 ? n984 : (n1146 ? n984 : 1'b0));
assign n6522 = /* LUT    3 20  1 */ (n318 ? 1'b0 : (n80 ? (n473 ? 1'b0 : !n330) : 1'b0));
assign n6523 = /* LUT    9  9  6 */ (n811 ? n1146 : (n878 ? 1'b0 : n1146));
assign n6524 = /* LUT    1 12  4 */ (n260 ? 1'b0 : (n252 ? !n261 : 1'b1));
assign n6525 = /* LUT    1  4  0 */ n34;
assign n6526 = /* LUT   20  8  4 */ n2806;
assign n6527 = /* LUT   12 22  5 */ (n1853 ? !n1847 : n1847);
assign n6528 = /* LUT   18 13  2 */ n2658;
assign n6529 = /* LUT   12 14  1 */ (n1622 ? (n1617 ? 1'b0 : n1623) : (n1617 ? n1623 : 1'b0));
assign n6530 = /* LUT   22 17  1 */ (n2156 ? (n2855 ? (n2293 ? 1'b0 : n2297) : 1'b0) : 1'b0);
assign n6534 = /* LUT   10  6  4 */ (n1281 ? n1267 : (n1267 ? !n5 : 1'b0));
assign n6535 = /* LUT    9 10  7 */ (n1138 ? (n1157 ? n1119 : 1'b0) : n1157);
assign n6536 = /* LUT    9  2  3 */ (n961 ? (n6 ? (n41 ? 1'b1 : !n964) : !n41) : (n6 ? (n41 ? 1'b1 : !n964) : 1'b1));
assign n6537 = /* LUT   22 20  6 */ (n2297 ? 1'b0 : (n2992 ? (n2156 ? n2293 : 1'b0) : 1'b0));
assign n6538 = /* LUT    3 16  3 */ (n612 ? 1'b0 : n80);
assign n6539 = /* LUT   21 16  5 */ (n2297 ? (n2156 ? (n2293 ? 1'b0 : n2428) : 1'b0) : 1'b0);
assign n6542 = /* LUT    3 15  7 */ (n447 ? (n453 ? (n602 ? n305 : 1'b0) : 1'b0) : 1'b0);
assign n6543 = /* LUT   10  7  5 */ (n5 ? (n1267 ? (n1427 ? 1'b0 : n1146) : n1146) : (n1267 ? 1'b0 : n1146));
assign n6544 = /* LUT   18  9  4 */ (n2624 ? (n2355 ? (n2348 ? 1'b0 : !n2364) : n2364) : (n2355 ? (n2348 ? n2364 : 1'b1) : n2364));
assign n6545 = /* LUT   22 21  7 */ (n2293 ? (n2297 ? (n2156 ? 1'b0 : n2848) : 1'b0) : 1'b0);
assign n6546 = /* LUT   22 13  3 */ (n2814 ? n2533 : 1'b0);
assign n6547 = /* LUT    4 20  3 */ (n627 ? (n624 ? n785 : (n648 ? 1'b0 : n785)) : n785);
assign n6548 = /* LUT    2 12  6 */ (n103 ? (n117 ? 1'b0 : n249) : (n117 ? 1'b0 : (n282 ? 1'b0 : n249)));
assign n6549 = /* LUT   13  5  5 */ n233;
assign n6550 = /* LUT    3  8  4 */ (n83 ? (n66 ? (n43 ? 1'b0 : !n209) : (n43 ? 1'b1 : !n209)) : 1'b0);
assign n6551 = /* LUT   18 10  5 */ (n2355 ? 1'b0 : (n2488 ? (n2629 ? 1'b1 : !n2364) : (n2629 ? n2364 : 1'b0)));
assign n6552 = /* LUT   18  2  1 */ n2449;
assign n6553 = /* LUT   15 14  2 */ n2113;
assign n6554 = /* LUT    5 17  1 */ (n93 ? !n5 : 1'b0);
assign n6558 = /* LUT    2 13  7 */ (n45 ? 1'b0 : n80);
assign n6559 = /* LUT   12  2  4 */ !n1541;
assign n6560 = /* LUT   13  6  6 */ (n1706 ? (n1704 ? 1'b0 : !n1696) : (n1704 ? 1'b0 : n1696));
assign n6561 = /* LUT    2  5  3 */ (n6 ? (n41 ? n194 : 1'b1) : (n41 ? 1'b1 : n36));
assign n6562 = /* LUT    3  1  1 */ n188;
assign n6563 = /* LUT    4 16  5 */ (n592 ? (n280 ? !n434 : 1'b1) : 1'b0);
assign n6564 = /* LUT   11 11  4 */ (n1603 ? (n1475 ? n1601 : !n1601) : (n1475 ? (n1330 ? n1601 : !n1601) : !n1601));
assign n6565 = /* LUT   14 19  5 */ (n2151 ? !n1503 : n1503);
assign n6566 = /* LUT   11  3  0 */ (n852 ? n980 : 1'b0);
assign n6567 = /* LUT   14 11  1 */ n1934;
assign n6568 = /* LUT   15 15  3 */ (n2269 ? (n1624 ? (n2130 ? 1'b1 : n2128) : 1'b1) : 1'b0);
assign n6569 = /* LUT    3  4  6 */ (n523 ? n371 : (n512 ? n371 : (n521 ? n371 : 1'b0)));
assign n6574 = /* LUT   22  5  3 */ (n2781 ? (n2775 ? (n2910 ? n2778 : 1'b0) : 1'b0) : 1'b0);
assign n6575 = /* LUT    5 13  3 */ (n271 ? (n582 ? 1'b0 : (n581 ? 1'b0 : !n113)) : 1'b0);
assign n6576 = /* LUT    4 17  6 */ (n80 ? (n605 ? 1'b1 : !n448) : !n448);
assign n6577 = /* LUT    4  9  2 */ (n559 ? (n711 ? 1'b0 : n400) : !n711);
assign n6578 = /* LUT   17 19  2 */ n2577;
assign n6579 = /* LUT   11  7  6 */ (n1419 ? n852 : 1'b1);
assign n6580 = /* LUT   17 18  6 */ (n2404 ? (n2403 ? 1'b0 : !n2010) : (n2403 ? 1'b0 : !n1829));
assign n6581 = /* LUT    7 13  1 */ (n1025 ? (n362 ? 1'b0 : !n698) : !n698);
assign n6582 = /* LUT   14 12  1 */ (n1453 ? (n2104 ? 1'b0 : (n2102 ? !n1933 : 1'b1)) : (n2102 ? !n1933 : 1'b1));
assign n6583 = /* LUT    5  5  4 */ n177;
assign n6584 = /* LUT    4  1  3 */ (n41 ? (n6 ? 1'b1 : !n501) : (n6 ? !n389 : 1'b1));
assign n6585 = /* LUT    8 12  4 */ n15;
assign n6586 = /* LUT    8  4  0 */ n233;
assign n6587 = /* LUT   16 15  5 */ n1631;
assign n6588 = /* LUT   23 14  5 */ (n3018 ? !n3020 : (n3032 ? !n3020 : (n2967 ? !n3020 : 1'b0)));
assign n6589 = /* LUT   20 18  2 */ n2012;
assign n6590 = /* LUT   15  3  6 */ (n1875 ? n1179 : 1'b0);
assign n6593 = /* LUT    7 17  7 */ !n621;
assign n6594 = /* LUT    7  9  3 */ (n1003 ? (n8 ? n998 : !n998) : (n8 ? !n998 : n998));
assign n6595 = /* LUT    8 13  5 */ n188;
assign n6596 = /* LUT    8  5  1 */ n354;
assign n6597 = /* LUT   14  7  7 */ (n1911 ? (n1937 ? (n1924 ? n1725 : 1'b0) : 1'b0) : 1'b0);
assign n6598 = /* LUT   17  7  5 */ (n2487 ? (n2066 ? n2484 : !n2315) : (n2066 ? n2484 : n2315));
assign n6599 = /* LUT    3 18  3 */ (n318 ? 1'b0 : (n112 ? (n300 ? 1'b0 : n460) : 1'b0));
assign n6600 = /* LUT    7  2  0 */ (n824 ? (n939 ? (n176 ? 1'b0 : !n499) : !n499) : !n499);
assign n6601 = /* LUT    9 21  6 */ (n1069 ? (n1219 ? !n924 : 1'b0) : (n437 ? (n1219 ? !n924 : 1'b0) : 1'b0));
assign n6602 = /* LUT   16  8  1 */ (n1931 ? 1'b0 : (n1700 ? !n2085 : n2085));
assign n6603 = /* LUT   13 13  0 */ (n1957 ? (n1790 ? 1'b0 : n1624) : 1'b0);
assign n6607 = /* LUT   13 16  5 */ (n1984 ? n852 : 1'b0);
assign n6608 = /* LUT    3 19  4 */ (n634 ? !n488 : n488);
assign n6609 = /* LUT   12 17  1 */ (n1358 ? (n5 ? 1'b0 : !n1652) : n1506);
assign n6610 = /* LUT   20  6  5 */ (n2788 ? !n2681 : n2681);
assign n6611 = /* LUT    2 20  0 */ (n327 ? n150 : (n475 ? n150 : 1'b0));
assign n6612 = /* LUT   10  9  4 */ (n811 ? !n1267 : (n5 ? (n1267 ? 1'b0 : n880) : !n1267));
assign n6613 = /* LUT    9 13  7 */ (n362 ? (n698 ? 1'b0 : !n1028) : !n698);
assign n6614 = /* LUT    9  5  3 */ n354;
assign n6615 = /* LUT   13 17  6 */ n1990;
assign n6618 = /* LUT   22 23  6 */ n2012;
assign n6619 = /* LUT    1 11  6 */ (n45 ? (n247 ? 1'b0 : (n79 ? 1'b0 : !n92)) : 1'b0);
assign n6620 = /* LUT   12 18  2 */ (n5 ? 1'b0 : (n1188 ? !n1652 : (n1652 ? 1'b0 : !n1639)));
assign n6621 = /* LUT   20  7  6 */ n2797;
assign n6622 = /* LUT   10 10  5 */ (n1302 ? 1'b0 : (n1158 ? 1'b0 : n1311));
assign n6623 = /* LUT   10  2  1 */ (n1400 ? (n6 ? (n1080 ? 1'b0 : n1077) : n1077) : (n6 ? n1077 : 1'b0));
assign n6624 = /* LUT   12 21  7 */ (n1523 ? n1501 : 1'b1);
assign n6625 = /* LUT    9  6  4 */ (n852 ? 1'b0 : n1116);
assign n6626 = /* LUT   18 12  4 */ n2647;
assign n6627 = /* LUT   18  4  0 */ n2173;
assign n6628 = /* LUT   22 16  3 */ n2012;
assign n6629 = /* LUT   13  9  1 */ (n1731 ? (n1890 ? 1'b0 : !n1598) : (n1890 ? 1'b0 : n1598));
assign n6630 = /* LUT   21 20  6 */ n2012;
assign n6631 = /* LUT   21 12  2 */ (n2509 ? (n2718 ? (n2503 ? !n2809 : 1'b0) : 1'b0) : (n2503 ? n2809 : 1'b0));
assign n6632 = /* LUT    3  3  0 */ n354;
assign n6633 = /* LUT   18 13  5 */ n2655;
assign n6634 = /* LUT    1  3  7 */ n14;
assign n6635 = /* LUT   18  5  1 */ n2332;
assign n6636 = /* LUT    5 20  1 */ (n627 ? (n618 ? (n621 ? 1'b0 : n648) : (n621 ? n648 : 1'b0)) : 1'b0);
assign n6637 = /* LUT   17 21  2 */ (n2429 ? (n2292 ? n2426 : 1'b0) : 1'b0);
assign n6638 = /* LUT   12  5  4 */ n15;
assign n3056 = /* CARRY 13  1  2 */ (n8 & n1533) | ((n8 | n1533) & n3226);
assign n413  = /* CARRY  2  8  3 */ (n227 & 1'b0) | ((n227 | 1'b0) & n412);
assign n741  = /* CARRY  4 12  2 */ (1'b0 & n579) | ((1'b0 | n579) & n740);
assign n3057 = /* CARRY  8 15  5 */ (n1023 & n917) | ((n1023 | n917) & n3227);
assign n2424 = /* CARRY 16 19  1 */ (1'b0 & n1987) | ((1'b0 | n1987) & n3081);
assign n2418 = /* CARRY 16 18  5 */ (n1993 & 1'b0) | ((n1993 | 1'b0) & n3229);
assign n3058 = /* CARRY  9 20  0 */ (n1043 & 1'b0) | ((n1043 | 1'b0) & n3322);
assign n1065 = /* CARRY  7 20  7 */ (n820 & 1'b0) | ((n820 | 1'b0) & n3230);
assign n3059 = /* CARRY  9 16  2 */ (n921 & 1'b0) | ((n921 | 1'b0) & n3083);
assign n2005 = /* CARRY 13 19  5 */ (n1648 & 1'b0) | ((n1648 | 1'b0) & n2004);
assign n3060 = /* CARRY  3 14  0 */ (1'b0 & n433) | ((1'b0 | n433) & n3347);
assign n3061 = /* CARRY  1  6  3 */ (1'b0 & n50) | ((1'b0 | n50) & n3231);
assign n1208 = /* CARRY  8 18  0 */ (1'b0 & n923) | ((1'b0 | n923) & n1205);
assign n3062 = /* CARRY 12  1  1 */ (1'b0 & n1402) | ((1'b0 | n1402) & n3232);
assign n3063 = /* CARRY  8 19  1 */ (n1045 & 1'b0) | ((n1045 | 1'b0) & n3085);
assign n2907 = /* CARRY 21  3  5 */ (n2765 & n8) | ((n2765 | n8) & n2906);
assign n3064 = /* CARRY  1 21  0 */ (1'b0 & n156) | ((1'b0 | n156) & n3401);
assign n3051 = /* CARRY 23 12  1 */ (1'b0 & n2809) | ((1'b0 | n2809) & n3233);
assign n3065 = /* CARRY  7 15  3 */ (n1020 & n1047) | ((n1020 | n1047) & n3234);
assign n3066 = /* CARRY  8  7  4 */ (n860 & n864) | ((n860 | n864) & n3088);
assign n2541 = /* CARRY 17 13  5 */ (n2256 & 1'b0) | ((n2256 | 1'b0) & n2540);
assign n3067 = /* CARRY  7  8  0 */ (n871 & 1'b0) | ((n871 | 1'b0) & n3419);
assign n2039 = /* CARRY 13 23  1 */ (1'b0 & n2031) | ((1'b0 | n2031) & n3089);
assign n2474 = /* CARRY 17  6  2 */ (n1416 & 1'b0) | ((n1416 | 1'b0) & n3090);
assign n3068 = /* CARRY  3 17  0 */ (1'b0 & n465) | ((1'b0 | n465) & n3432);
assign n1975 = /* CARRY 13 15  2 */ (n1806 & n1788) | ((n1806 | n1788) & n1974);
assign n3069 = /* CARRY  3 14  3 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n599);
assign n1767 = /* CARRY 12 12  0 */ (n1607 & n212) | ((n1607 | n212) & n3454);
assign n3035 = /* CARRY 22 15  0 */ (n3024 & n8) | ((n3024 | n8) & n3031);
assign n3070 = /* CARRY  4 18  2 */ (n8 & 1'b0) | ((n8 | 1'b0) & n778);
assign n3071 = /* CARRY 11  1  0 */ (1'b0 & n1531) | ((1'b0 | n1531) & n3477);
assign n1205 = /* CARRY  8 17  7 */ (1'b0 & n821) | ((1'b0 | n821) & n3238);
assign n3072 = /* CARRY 10 18  0 */ (1'b0 & n188) | ((1'b0 | n188) & n3493);
assign n1394 = /* CARRY  9 22  3 */ (1'b0 & n931) | ((1'b0 | n931) & n1393);
assign n3073 = /* CARRY  7 15  6 */ (n1022 & n920) | ((n1022 | n920) & n3096);
assign n3074 = /* CARRY 20  1  0 */ (n2314 & 1'b0) | ((n2314 | 1'b0) & n3525);
assign n3027 = /* CARRY 22 14  2 */ (n8 & n2966) | ((n8 | n2966) & n3026);
assign n2269 = /* CARRY 15 15  2 */ (n1979 & n1766) | ((n1979 | n1766) & n3242);
assign n2284 = /* CARRY 15 18  7 */ (n1995 & n8) | ((n1995 | n8) & n3243);
assign n3075 = /* CARRY 12  3  4 */ (1'b0 & n1532) | ((1'b0 | n1532) & n3244);
assign n2577 = /* CARRY 17 19  1 */ (1'b0 & n2292) | ((1'b0 | n2292) & n3245);
assign n393  = /* CARRY  2  6  2 */ (1'b0 & n176) | ((1'b0 | n176) & n392);
assign n3076 = /* CARRY 11  1  3 */ (n1535 & n8) | ((n1535 | n8) & n3098);
assign n3077 = /* CARRY  9 18  0 */ (1'b0 & n1034) | ((1'b0 | n1034) & n3588);
assign n1058 = /* CARRY  7 18  7 */ (n821 & 1'b0) | ((n821 | 1'b0) & n3099);
assign n2487 = /* CARRY 17  7  4 */ (1'b0 & n2178) | ((1'b0 | n2178) & n3246);
assign n3078 = /* CARRY 10 18  3 */ (n15 & 1'b0) | ((n15 | 1'b0) & n3100);
assign n3047 = /* CARRY 23  2  7 */ (n2892 & n8) | ((n2892 | n8) & n3046);
assign n3079 = /* CARRY  1  8  0 */ (n209 & n57) | ((n209 | n57) & n3611);
assign n1990 = /* CARRY 13 17  5 */ (1'b0 & n1780) | ((1'b0 | n1780) & n3247);
assign n2797 = /* CARRY 20  7  5 */ (n8 & n2692) | ((n8 | n2692) & n3248);
assign n2161 = /* CARRY 14 23  0 */ (n1846 & n2018) | ((n1846 | n2018) & n3640);
assign n2611 = /* CARRY 18  6  1 */ (1'b0 & n2465) | ((1'b0 | n2465) & n3250);
assign n2963 = /* CARRY 21 13  1 */ (1'b0 & n2824) | ((1'b0 | n2824) & n3101);
assign n740  = /* CARRY  4 12  1 */ (n113 & 1'b0) | ((n113 | 1'b0) & n3251);
assign n1198 = /* CARRY  8 16  0 */ (n923 & 1'b0) | ((n923 | 1'b0) & n1197);
assign n3080 = /* CARRY  4 13  2 */ (n8 & n433) | ((n8 | n433) & n3252);
assign n3081 = /* CARRY 16 19  0 */ (1'b0 & n8) | ((1'b0 | n8) & n2419);
assign n3082 = /* CARRY 17 11  0 */ (1'b0 & n2377) | ((1'b0 | n2377) & n3687);
assign n3083 = /* CARRY  9 16  1 */ (1'b0 & n1045) | ((1'b0 | n1045) & n3254);
assign n3084 = /* CARRY  7  9  5 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1005);
assign n2017 = /* CARRY 13 20  5 */ (n1648 & n8) | ((n1648 | n8) & n2016);
assign n476  = /* CARRY  2 19  1 */ (n319 & 1'b0) | ((n319 | 1'b0) & n3256);
assign n237  = /* CARRY  1  8  3 */ (1'b0 & n8) | ((1'b0 | n8) & n236);
assign n2917 = /* CARRY 21  4  0 */ (n2672 & n8) | ((n2672 | n8) & n2909);
assign n3085 = /* CARRY  8 19  0 */ (n922 & 1'b0) | ((n922 | 1'b0) & n3742);
assign n3086 = /* CARRY 13  1  4 */ (n8 & n1530) | ((n8 | n1530) & n3257);
assign n743  = /* CARRY  4 12  4 */ (1'b0 & n581) | ((1'b0 | n581) & n742);
assign n3087 = /* CARRY 17 14  0 */ (n2394 & 1'b0) | ((n2394 | 1'b0) & n3765);
assign n1197 = /* CARRY  8 15  7 */ (n1021 & n821) | ((n1021 | n821) & n3259);
assign n3088 = /* CARRY  8  7  3 */ (n863 & n855) | ((n863 | n855) & n3260);
assign n3089 = /* CARRY 13 23  0 */ (n2030 & 1'b0) | ((n2030 | 1'b0) & n3775);
assign n2419 = /* CARRY 16 18  7 */ (1'b0 & n1995) | ((1'b0 | n1995) & n3261);
assign n3090 = /* CARRY 17  6  1 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2473);
assign n1383 = /* CARRY  9 20  2 */ (n8 & n1061) | ((n8 | n1061) & n1382);
assign n2837 = /* CARRY 20 14  1 */ (n2820 & n8) | ((n2820 | n8) & n3109);
assign n3091 = /* CARRY  9 16  4 */ (n919 & 1'b0) | ((n919 | 1'b0) & n3110);
assign n599  = /* CARRY  3 14  2 */ (1'b0 & n588) | ((1'b0 | n588) & n3263);
assign n3092 = /* CARRY  1  6  5 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n216);
assign n3093 = /* CARRY 21  7  0 */ (n2794 & 1'b0) | ((n2794 | 1'b0) & n3823);
assign n3094 = /* CARRY 18  1  0 */ (n2314 & 1'b0) | ((n2314 | 1'b0) & n3836);
assign n3095 = /* CARRY 12  1  3 */ (1'b0 & n1535) | ((1'b0 | n1535) & n3266);
assign n813  = /* CARRY  5 11  1 */ (n731 & 1'b0) | ((n731 | 1'b0) & n3267);
assign n2909 = /* CARRY 21  3  7 */ (n8 & n2767) | ((n8 | n2767) & n2908);
assign n713  = /* CARRY  4  8  1 */ (n401 & n8) | ((n401 | n8) & n3113);
assign n337  = /* CARRY  1 21  2 */ (n153 & 1'b0) | ((n153 | 1'b0) & n336);
assign n3096 = /* CARRY  7 15  5 */ (n1023 & n909) | ((n1023 | n909) & n3269);
assign n992  = /* CARRY  7  8  2 */ (n866 & 1'b0) | ((n866 | 1'b0) & n991);
assign n1977 = /* CARRY 13 15  4 */ (n1803 & n1804) | ((n1803 | n1804) & n1976);
assign n3026 = /* CARRY 22 14  1 */ (n8 & n3019) | ((n8 | n3019) & n3270);
assign n1769 = /* CARRY 12 12  2 */ (n1766 & n1600) | ((n1766 | n1600) & n1768);
assign n3036 = /* CARRY 22 15  2 */ (n3022 & n8) | ((n3022 | n8) & n3119);
assign n392  = /* CARRY  2  6  1 */ (1'b0 & n41) | ((1'b0 | n41) & n3272);
assign n3097 = /* CARRY  4 18  4 */ (n8 & 1'b0) | ((n8 | 1'b0) & n779);
assign n3098 = /* CARRY 11  1  2 */ (n8 & n1533) | ((n8 | n1533) & n3273);
assign n3099 = /* CARRY  7 18  6 */ (n913 & 1'b0) | ((n913 | 1'b0) & n3274);
assign n3100 = /* CARRY 10 18  2 */ (1'b0 & n179) | ((1'b0 | n179) & n3275);
assign n458  = /* CARRY  2 17  1 */ (n456 & 1'b0) | ((n456 | 1'b0) & n3278);
assign n2760 = /* CARRY 20  1  2 */ (n2447 & 1'b0) | ((n2447 | 1'b0) & n2759);
assign n3101 = /* CARRY 21 13  0 */ (n2818 & 1'b0) | ((n2818 | 1'b0) & n3975);
assign n3102 = /* CARRY  4 21  0 */ (n642 & 1'b0) | ((n642 | 1'b0) & n3979);
assign n570  = /* CARRY  3  9  1 */ (n407 & n566) | ((n407 | n566) & n569);
assign n1071 = /* CARRY  7 21  1 */ (1'b0 & n8) | ((1'b0 | n8) & n1070);
assign n1680 = /* CARRY 12  3  6 */ (1'b0 & n1529) | ((1'b0 | n1529) & n3280);
assign n2578 = /* CARRY 17 19  3 */ (n2426 & 1'b0) | ((n2426 | 1'b0) & n3281);
assign n395  = /* CARRY  2  6  4 */ (n51 & 1'b0) | ((n51 | 1'b0) & n394);
assign n3103 = /* CARRY  5  6  0 */ (1'b0 & n213) | ((1'b0 | n213) & n4019);
assign n3104 = /* CARRY  9 17  1 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1371);
assign n1005 = /* CARRY  7  9  4 */ (n999 & n8) | ((n999 | n8) & n1004);
assign n3105 = /* CARRY  9 18  2 */ (n914 & 1'b0) | ((n914 | 1'b0) & n3125);
assign n298  = /* CARRY  1 16  1 */ (1'b0 & n119) | ((1'b0 | n119) & n3126);
assign n3106 = /* CARRY 10 18  5 */ (1'b0 & n233) | ((1'b0 | n233) & n3127);
assign n236  = /* CARRY  1  8  2 */ (n234 & n47) | ((n234 | n47) & n3283);
assign n1991 = /* CARRY 13 17  7 */ (n1650 & 1'b0) | ((n1650 | 1'b0) & n3282);
assign n2798 = /* CARRY 20  7  7 */ (n8 & n2691) | ((n8 | n2691) & n3284);
assign n3107 = /* CARRY  2  9  0 */ (1'b0 & n209) | ((1'b0 | n209) & n4076);
assign n2163 = /* CARRY 14 23  2 */ (n1843 & n2028) | ((n1843 | n2028) & n2162);
assign n1220 = /* CARRY  8 20  0 */ (n911 & 1'b0) | ((n911 | 1'b0) & n1214);
assign n2613 = /* CARRY 18  6  3 */ (1'b0 & n2467) | ((1'b0 | n2467) & n2612);
assign n742  = /* CARRY  4 12  3 */ (1'b0 & n580) | ((1'b0 | n580) & n741);
assign n751  = /* CARRY  4 13  4 */ (1'b0 & n588) | ((1'b0 | n588) & n3129);
assign n3108 = /* CARRY 16 19  2 */ (1'b0 & n8) | ((1'b0 | n8) & n2424);
assign n3109 = /* CARRY 20 14  0 */ (n2824 & 1'b0) | ((n2824 | 1'b0) & n4116);
assign n3110 = /* CARRY  9 16  3 */ (n1047 & 1'b0) | ((n1047 | 1'b0) & n3059);
assign n326  = /* CARRY  1 19  1 */ (n135 & 1'b0) | ((n135 | 1'b0) & n3131);
assign n3111 = /* CARRY 21  8  0 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2944);
assign n2919 = /* CARRY 21  4  2 */ (n8 & n2914) | ((n8 | n2914) & n2918);
assign n3112 = /* CARRY  8 19  2 */ (1'b0 & n921) | ((1'b0 | n921) & n3063);
assign n3113 = /* CARRY  4  8  0 */ (1'b0 & n398) | ((1'b0 | n398) & n4183);
assign n3114 = /* CARRY 13  1  6 */ (n1534 & 1'b0) | ((n1534 | 1'b0) & n3133);
assign n3115 = /* CARRY 17 18  0 */ (1'b0 & n2415) | ((1'b0 | n2415) & n4191);
assign n1051 = /* CARRY  7 16  0 */ (1'b0 & n911) | ((1'b0 | n911) & n1048);
assign n2546 = /* CARRY 17 14  2 */ (n2391 & 1'b0) | ((n2391 | 1'b0) & n2545);
assign n1127 = /* CARRY  8  7  5 */ (n985 & n988) | ((n985 | n988) & n3066);
assign n991  = /* CARRY  7  8  1 */ (n865 & 1'b0) | ((n865 | 1'b0) & n3067);
assign n2040 = /* CARRY 13 23  2 */ (n2032 & 1'b0) | ((n2032 | 1'b0) & n2039);
assign n3116 = /* CARRY 17  6  3 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2474);
assign n1385 = /* CARRY  9 20  4 */ (n1050 & n8) | ((n1050 | n8) & n1384);
assign n3117 = /* CARRY  9 12  0 */ (1'b0 & n817) | ((1'b0 | n817) & n4219);
assign n3118 = /* CARRY  9 16  6 */ (n920 & n8) | ((n920 | n8) & n3134);
assign n1768 = /* CARRY 12 12  1 */ (n1765 & n1606) | ((n1765 | n1606) & n1767);
assign n3119 = /* CARRY 22 15  1 */ (1'b0 & n8) | ((1'b0 | n8) & n3035);
assign n3120 = /* CARRY 21  7  2 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2941);
assign n1059 = /* CARRY  7 19  0 */ (n923 & 1'b0) | ((n923 | 1'b0) & n1058);
assign n3121 = /* CARRY 12  1  5 */ (n1532 & 1'b0) | ((n1532 | 1'b0) & n3138);
assign n815  = /* CARRY  5 11  3 */ (n732 & 1'b0) | ((n732 | 1'b0) & n814);
assign n3122 = /* CARRY  1 13  0 */ (1'b0 & n96) | ((1'b0 | n96) & n4296);
assign n1048 = /* CARRY  7 15  7 */ (n1021 & n820) | ((n1021 | n820) & n3073);
assign n994  = /* CARRY  7  8  4 */ (n868 & 1'b0) | ((n868 | 1'b0) & n993);
assign n569  = /* CARRY  3  9  0 */ (n406 & n565) | ((n406 | n565) & n4314);
assign n804  = /* CARRY  4 22  0 */ (n488 & 1'b0) | ((n488 | 1'b0) & n803);
assign n3028 = /* CARRY 22 14  3 */ (n3023 & n8) | ((n3023 | n8) & n3027);
assign n394  = /* CARRY  2  6  3 */ (n200 & 1'b0) | ((n200 | 1'b0) & n393);
assign n3123 = /* CARRY  4 18  6 */ (n8 & 1'b0) | ((n8 | 1'b0) & n780);
assign n3124 = /* CARRY 11  1  4 */ (n8 & n1530) | ((n8 | n1530) & n3076);
assign n3125 = /* CARRY  9 18  1 */ (1'b0 & n1053) | ((1'b0 | n1053) & n3077);
assign n3126 = /* CARRY  1 16  0 */ (n294 & 1'b0) | ((n294 | 1'b0) & n4373);
assign n3127 = /* CARRY 10 18  4 */ (n354 & 1'b0) | ((n354 | 1'b0) & n3078);
assign n308  = /* CARRY  1 17  1 */ (1'b0 & n123) | ((1'b0 | n123) & n3145);
assign n3128 = /* CARRY  3 13  1 */ (n430 & 1'b0) | ((n430 | 1'b0) & n3146);
assign n2162 = /* CARRY 14 23  1 */ (n1528 & n2029) | ((n1528 | n2029) & n2161);
assign n2612 = /* CARRY 18  6  2 */ (n2466 & 1'b0) | ((n2466 | 1'b0) & n2611);
assign n2964 = /* CARRY 21 13  2 */ (n2820 & 1'b0) | ((n2820 | 1'b0) & n2963);
assign n799  = /* CARRY  4 21  2 */ (1'b0 & n777) | ((1'b0 | n777) & n798);
assign n572  = /* CARRY  3  9  3 */ (n405 & n567) | ((n405 | n567) & n571);
assign n3129 = /* CARRY  4 13  3 */ (n444 & 1'b0) | ((n444 | 1'b0) & n3080);
assign n3130 = /* CARRY  8 17  1 */ (n1053 & 1'b0) | ((n1053 | 1'b0) & n3147);
assign n2579 = /* CARRY 17 19  5 */ (n2156 & 1'b0) | ((n2156 | 1'b0) & n3148);
assign n2520 = /* CARRY 17 11  1 */ (n2375 & 1'b0) | ((n2375 | 1'b0) & n3082);
assign n3131 = /* CARRY  1 19  0 */ (n141 & 1'b0) | ((n141 | 1'b0) & n4455);
assign n3132 = /* CARRY  9 18  4 */ (1'b0 & n915) | ((1'b0 | n915) & n3150);
assign n2918 = /* CARRY 21  4  1 */ (n8 & n2915) | ((n8 | n2915) & n2917);
assign n2281 = /* CARRY 15 18  1 */ (n8 & n2142) | ((n8 | n2142) & n3152);
assign n421  = /* CARRY  2  9  2 */ (1'b0 & n8) | ((1'b0 | n8) & n420);
assign n2165 = /* CARRY 14 23  4 */ (n1848 & n8) | ((n1848 | n8) & n2164);
assign n3133 = /* CARRY 13  1  5 */ (1'b0 & n1532) | ((1'b0 | n1532) & n3086);
assign n2615 = /* CARRY 18  6  5 */ (n2469 & 1'b0) | ((n2469 | 1'b0) & n2614);
assign n2931 = /* CARRY 21  5  1 */ (n2777 & n8) | ((n2777 | n8) & n2930);
assign n2545 = /* CARRY 17 14  1 */ (n2266 & 1'b0) | ((n2266 | 1'b0) & n3087);
assign n1384 = /* CARRY  9 20  3 */ (n8 & n1019) | ((n8 | n1019) & n1383);
assign n3043 = /* CARRY 23  2  1 */ (n8 & n2890) | ((n8 | n2890) & n3157);
assign n2838 = /* CARRY 20 14  2 */ (n2821 & n8) | ((n2821 | n8) & n2837);
assign n3134 = /* CARRY  9 16  5 */ (n909 & n8) | ((n909 | n8) & n3091);
assign n3135 = /* CARRY 12 21  0 */ (1'b0 & n1833) | ((1'b0 | n1833) & n4557);
assign n2941 = /* CARRY 21  7  1 */ (n2790 & 1'b0) | ((n2790 | 1'b0) & n3093);
assign n3136 = /* CARRY 21  8  2 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2948);
assign n2596 = /* CARRY 18  1  1 */ (n2595 & n8) | ((n2595 | n8) & n3094);
assign n3137 = /* CARRY 12  2  0 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1667);
assign n3138 = /* CARRY 12  1  4 */ (n1530 & n8) | ((n1530 | n8) & n3095);
assign n814  = /* CARRY  5 11  2 */ (1'b0 & n730) | ((1'b0 | n730) & n813);
assign n2921 = /* CARRY 21  4  4 */ (n2670 & n8) | ((n2670 | n8) & n2920);
assign n3139 = /* CARRY  8 19  4 */ (n919 & 1'b0) | ((n919 | 1'b0) & n3160);
assign n3140 = /* CARRY  7 20  0 */ (n922 & 1'b0) | ((n922 | 1'b0) & n4609);
assign n2570 = /* CARRY 17 18  2 */ (1'b0 & n2410) | ((1'b0 | n2410) & n2569);
assign n993  = /* CARRY  7  8  3 */ (n867 & 1'b0) | ((n867 | 1'b0) & n992);
assign n2042 = /* CARRY 13 23  4 */ (n2034 & 1'b0) | ((n2034 | 1'b0) & n2041);
assign n3141 = /* CARRY 17  6  5 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2475);
assign n1387 = /* CARRY  9 20  6 */ (n8 & n931) | ((n8 | n931) & n1386);
assign n2785 = /* CARRY 20  6  1 */ (1'b0 & n2677) | ((1'b0 | n2677) & n3164);
assign n3142 = /* CARRY 12 12  3 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1769);
assign n3037 = /* CARRY 22 15  3 */ (n2973 & n8) | ((n2973 | n8) & n3036);
assign n789  = /* CARRY  4 19  1 */ (n334 & n8) | ((n334 | n8) & n788);
assign n780  = /* CARRY  4 18  5 */ (n621 & n8) | ((n621 | n8) & n3097);
assign n3143 = /* CARRY 21  7  4 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2942);
assign n3144 = /* CARRY  8 15  1 */ (n910 & n1053) | ((n910 | n1053) & n3165);
assign n1667 = /* CARRY 12  1  7 */ (n1529 & 1'b0) | ((n1529 | 1'b0) & n3167);
assign n2416 = /* CARRY 16 18  1 */ (1'b0 & n2142) | ((1'b0 | n2142) & n3168);
assign n3145 = /* CARRY  1 17  0 */ (n126 & 1'b0) | ((n126 | 1'b0) & n4702);
assign n2001 = /* CARRY 13 19  1 */ (1'b0 & n1836) | ((1'b0 | n1836) & n3171);
assign n3146 = /* CARRY  3 13  0 */ (1'b0 & n589) | ((1'b0 | n589) & n4730);
assign n798  = /* CARRY  4 21  1 */ (1'b0 & n630) | ((1'b0 | n630) & n3102);
assign n571  = /* CARRY  3  9  2 */ (n568 & n409) | ((n568 | n409) & n570);
assign n2276 = /* CARRY 15 16  1 */ (n1624 & 1'b0) | ((n1624 | 1'b0) & n3172);
assign n3029 = /* CARRY 22 14  5 */ (n8 & n3021) | ((n8 | n3021) & n3173);
assign n3147 = /* CARRY  8 17  0 */ (1'b0 & n1034) | ((1'b0 | n1034) & n4763);
assign n3148 = /* CARRY 17 19  4 */ (1'b0 & n8) | ((1'b0 | n8) & n2578);
assign n809  = /* CARRY  5  6  1 */ (n8 & n410) | ((n8 | n410) & n3103);
assign n3149 = /* CARRY 11  1  6 */ (n1534 & 1'b0) | ((n1534 | 1'b0) & n3176);
assign n3150 = /* CARRY  9 18  3 */ (n918 & 1'b0) | ((n918 | 1'b0) & n3105);
assign n3151 = /* CARRY 10 18  6 */ (n177 & 1'b0) | ((n177 | 1'b0) & n3106);
assign n3152 = /* CARRY 15 18  0 */ (n1997 & 1'b0) | ((n1997 | 1'b0) & n4817);
assign n420  = /* CARRY  2  9  1 */ (n208 & 1'b0) | ((n208 | 1'b0) & n3107);
assign n3153 = /* CARRY  3 13  3 */ (1'b0 & n433) | ((1'b0 | n433) & n3179);
assign n3154 = /* CARRY 13  2  0 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1862);
assign n2164 = /* CARRY 14 23  3 */ (n1845 & n2026) | ((n1845 | n2026) & n2163);
assign n2288 = /* CARRY 15 19  1 */ (n8 & n1987) | ((n8 | n1987) & n3180);
assign n2614 = /* CARRY 18  6  4 */ (n2468 & 1'b0) | ((n2468 | 1'b0) & n2613);
assign n800  = /* CARRY  4 21  4 */ (n621 & 1'b0) | ((n621 | 1'b0) & n3181);
assign n2930 = /* CARRY 21  5  0 */ (n2776 & n8) | ((n2776 | n8) & n2924);
assign n2425 = /* CARRY 16 19  3 */ (n2280 & 1'b0) | ((n2280 | 1'b0) & n3108);
assign n3155 = /* CARRY  7 18  0 */ (1'b0 & n1034) | ((1'b0 | n1034) & n4856);
assign n3156 = /* CARRY  8 17  3 */ (1'b0 & n918) | ((1'b0 | n918) & n3183);
assign n2580 = /* CARRY 17 19  7 */ (n2293 & 1'b0) | ((n2293 | 1'b0) & n3184);
assign n3157 = /* CARRY 23  2  0 */ (n3011 & 1'b0) | ((n3011 | 1'b0) & n4871);
assign n3048 = /* CARRY 23  3  1 */ (n8 & n2896) | ((n8 | n2896) & n3185);
assign n3158 = /* CARRY 12 22  0 */ (n1846 & 1'b0) | ((n1846 | 1'b0) & n4892);
assign n3159 = /* CARRY  9 18  6 */ (1'b0 & n913) | ((1'b0 | n913) & n3186);
assign n2948 = /* CARRY 21  8  1 */ (1'b0 & n2804) | ((1'b0 | n2804) & n3111);
assign n2147 = /* CARRY 14 19  0 */ (n1966 & n2007) | ((n1966 | n2007) & n4925);
assign n2920 = /* CARRY 21  4  3 */ (n8 & n2912) | ((n8 | n2912) & n2919);
assign n2282 = /* CARRY 15 18  3 */ (n1992 & n8) | ((n1992 | n8) & n3188);
assign n3160 = /* CARRY  8 19  3 */ (1'b0 & n1047) | ((1'b0 | n1047) & n3112);
assign n3161 = /* CARRY 12  3  0 */ (n1402 & 1'b0) | ((n1402 | 1'b0) & n4937);
assign n1862 = /* CARRY 13  1  7 */ (n1529 & 1'b0) | ((n1529 | 1'b0) & n3114);
assign n2569 = /* CARRY 17 18  1 */ (1'b0 & n2409) | ((1'b0 | n2409) & n3115);
assign n3162 = /* CARRY  7 16  1 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1051);
assign n2547 = /* CARRY 17 14  3 */ (1'b0 & n2392) | ((1'b0 | n2392) & n2546);
assign n2041 = /* CARRY 13 23  3 */ (n2033 & 1'b0) | ((n2033 | 1'b0) & n2040);
assign n2485 = /* CARRY 17  7  0 */ (1'b0 & n852) | ((1'b0 | n852) & n2477);
assign n2475 = /* CARRY 17  6  4 */ (1'b0 & n1125) | ((1'b0 | n1125) & n3116);
assign n1386 = /* CARRY  9 20  5 */ (n1189 & n8) | ((n1189 | n8) & n1385);
assign n1332 = /* CARRY  9 12  1 */ (n8 & n1322) | ((n8 | n1322) & n3117);
assign n3163 = /* CARRY 23  2  3 */ (1'b0 & n8) | ((1'b0 | n8) & n3044);
assign n3164 = /* CARRY 20  6  0 */ (1'b0 & n2621) | ((1'b0 | n2621) & n4981);
assign n1988 = /* CARRY 13 17  1 */ (1'b0 & n1978) | ((1'b0 | n1978) & n3190);
assign n1368 = /* CARRY  9 16  7 */ (n820 & 1'b0) | ((n820 | 1'b0) & n3118);
assign n2795 = /* CARRY 20  7  1 */ (n8 & n2790) | ((n8 | n2790) & n3191);
assign n1840 = /* CARRY 12 21  2 */ (n1834 & 1'b0) | ((n1834 | 1'b0) & n1839);
assign n788  = /* CARRY  4 19  0 */ (n477 & n8) | ((n477 | n8) & n781);
assign n2942 = /* CARRY 21  7  3 */ (1'b0 & n2690) | ((1'b0 | n2690) & n3120);
assign n3165 = /* CARRY  8 15  0 */ (n1034 & n1028) | ((n1034 | n1028) & n5035);
assign n2598 = /* CARRY 18  1  3 */ (n2448 & n8) | ((n2448 | n8) & n2597);
assign n3166 = /* CARRY  7 19  1 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1059);
assign n3167 = /* CARRY 12  1  6 */ (n1534 & 1'b0) | ((n1534 | 1'b0) & n3121);
assign n3168 = /* CARRY 16 18  0 */ (1'b0 & n1997) | ((1'b0 | n1997) & n5046);
assign n3169 = /* CARRY  8 19  6 */ (n920 & 1'b0) | ((n920 | 1'b0) & n3193);
assign n3170 = /* CARRY  7 20  2 */ (1'b0 & n921) | ((1'b0 | n921) & n3194);
assign n2572 = /* CARRY 17 18  4 */ (1'b0 & n2412) | ((1'b0 | n2412) & n2571);
assign n2510 = /* CARRY 17 10  0 */ (n2507 & n1622) | ((n2507 | n1622) & n5064);
assign n279  = /* CARRY  1 13  1 */ (1'b0 & n94) | ((1'b0 | n94) & n3122);
assign n3171 = /* CARRY 13 19  0 */ (n1822 & 1'b0) | ((n1822 | 1'b0) & n5073);
assign n2013 = /* CARRY 13 20  1 */ (n1836 & n8) | ((n1836 | n8) & n3196);
assign n995  = /* CARRY  7  8  5 */ (1'b0 & n869) | ((1'b0 | n869) & n994);
assign n622  = /* CARRY  3 18  1 */ (1'b0 & n312) | ((1'b0 | n312) & n3197);
assign n2477 = /* CARRY 17  6  7 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2476);
assign n2787 = /* CARRY 20  6  3 */ (n2679 & 1'b0) | ((n2679 | 1'b0) & n2786);
assign n3172 = /* CARRY 15 16  0 */ (1'b0 & n1790) | ((1'b0 | n1790) & n5098);
assign n3173 = /* CARRY 22 14  4 */ (1'b0 & n8) | ((1'b0 | n8) & n3028);
assign n3174 = /* CARRY 21  3  0 */ (n2901 & 1'b0) | ((n2901 | 1'b0) & n5117);
assign n781  = /* CARRY  4 18  7 */ (n620 & n8) | ((n620 | n8) & n3123);
assign n3175 = /* CARRY 21  7  6 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2943);
assign n3176 = /* CARRY 11  1  5 */ (1'b0 & n1532) | ((1'b0 | n1532) & n3124);
assign n3177 = /* CARRY  8 15  3 */ (n1020 & n918) | ((n1020 | n918) & n3200);
assign n3178 = /* CARRY 17 13  0 */ (1'b0 & n2257) | ((1'b0 | n2257) & n5145);
assign n2417 = /* CARRY 16 18  3 */ (1'b0 & n1992) | ((1'b0 | n1992) & n3201);
assign n3179 = /* CARRY  3 13  2 */ (n424 & n8) | ((n424 | n8) & n3128);
assign n3180 = /* CARRY 15 19  0 */ (1'b0 & n8) | ((1'b0 | n8) & n2284);
assign n3181 = /* CARRY  4 21  3 */ (1'b0 & n8) | ((1'b0 | n8) & n799);
assign n3182 = /* CARRY  3  9  4 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n572);
assign n3031 = /* CARRY 22 14  7 */ (n8 & 1'b0) | ((n8 | 1'b0) & n3030);
assign n3183 = /* CARRY  8 17  2 */ (n914 & 1'b0) | ((n914 | 1'b0) & n3130);
assign n3184 = /* CARRY 17 19  6 */ (1'b0 & n8) | ((1'b0 | n8) & n2579);
assign n3185 = /* CARRY 23  3  0 */ (1'b0 & n8) | ((1'b0 | n8) & n3047);
assign n3186 = /* CARRY  9 18  5 */ (1'b0 & n917) | ((1'b0 | n917) & n3132);
assign n3187 = /* CARRY  2 21  0 */ (1'b0 & n331) | ((1'b0 | n331) & n5251);
assign n2784 = /* CARRY 20  5  1 */ (1'b0 & n2674) | ((1'b0 | n2674) & n3206);
assign n3188 = /* CARRY 15 18  2 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2281);
assign n590  = /* CARRY  3 13  5 */ (n588 & 1'b0) | ((n588 | 1'b0) & n3207);
assign n2166 = /* CARRY 14 23  5 */ (n8 & n1847) | ((n8 | n1847) & n2165);
assign n2289 = /* CARRY 15 19  3 */ (n8 & n2280) | ((n8 | n2280) & n3208);
assign n802  = /* CARRY  4 21  6 */ (1'b0 & n477) | ((1'b0 | n477) & n801);
assign n2932 = /* CARRY 21  5  2 */ (n2926 & n8) | ((n2926 | n8) & n2931);
assign n3189 = /* CARRY  7 18  2 */ (1'b0 & n914) | ((1'b0 | n914) & n3209);
assign n1147 = /* CARRY  8  9  1 */ (n880 & 1'b0) | ((n880 | 1'b0) & n3211);
assign n3044 = /* CARRY 23  2  2 */ (n3005 & n8) | ((n3005 | n8) & n3043);
assign n3190 = /* CARRY 13 17  0 */ (n1980 & 1'b0) | ((n1980 | 1'b0) & n5316);
assign n3049 = /* CARRY 23  3  3 */ (n8 & n2897) | ((n8 | n2897) & n3213);
assign n3191 = /* CARRY 20  7  0 */ (1'b0 & n2794) | ((1'b0 | n2794) & n5327);
assign n1839 = /* CARRY 12 21  1 */ (n1831 & 1'b0) | ((n1831 | 1'b0) & n3135);
assign n2805 = /* CARRY 20  8  1 */ (n2804 & n8) | ((n2804 | n8) & n3214);
assign n1851 = /* CARRY 12 22  2 */ (1'b0 & n1843) | ((1'b0 | n1843) & n1850);
assign n555  = /* CARRY  3  8  1 */ (1'b0 & n53) | ((1'b0 | n53) & n3215);
assign n2949 = /* CARRY 21  8  3 */ (n2803 & 1'b0) | ((n2803 | 1'b0) & n3136);
assign n2597 = /* CARRY 18  1  2 */ (n8 & n2447) | ((n8 | n2447) & n2596);
assign n1602 = /* CARRY 11 11  1 */ (n1473 & n8) | ((n1473 | n8) & n3216);
assign n2149 = /* CARRY 14 19  2 */ (n1982 & n2006) | ((n1982 | n2006) & n2148);
assign n3192 = /* CARRY 15 15  0 */ (n212 & n2135) | ((n212 | n2135) & n5378);
assign n2922 = /* CARRY 21  4  5 */ (n8 & n2773) | ((n8 | n2773) & n2921);
assign n2283 = /* CARRY 15 18  5 */ (n1993 & n8) | ((n1993 | n8) & n3217);
assign n3193 = /* CARRY  8 19  5 */ (n909 & 1'b0) | ((n909 | 1'b0) & n3139);
assign n3194 = /* CARRY  7 20  1 */ (1'b0 & n1045) | ((1'b0 | n1045) & n3140);
assign n2571 = /* CARRY 17 18  3 */ (n2411 & 1'b0) | ((n2411 | 1'b0) & n2570);
assign n2549 = /* CARRY 17 14  5 */ (n2267 & 1'b0) | ((n2267 | 1'b0) & n2548);
assign n3195 = /* CARRY  7  9  0 */ (n875 & 1'b0) | ((n875 | 1'b0) & n5404);
assign n3196 = /* CARRY 13 20  0 */ (n1822 & 1'b0) | ((n1822 | 1'b0) & n5408);
assign n2043 = /* CARRY 13 23  5 */ (n2035 & 1'b0) | ((n2035 | 1'b0) & n2042);
assign n3197 = /* CARRY  3 18  0 */ (1'b0 & n309) | ((1'b0 | n309) & n5413);
assign n2476 = /* CARRY 17  6  6 */ (1'b0 & n1126) | ((1'b0 | n1126) & n3141);
assign n1388 = /* CARRY  9 20  7 */ (n907 & n8) | ((n907 | n8) & n1387);
assign n632  = /* CARRY  3 19  1 */ (n620 & 1'b0) | ((n620 | 1'b0) & n3221);
assign n2786 = /* CARRY 20  6  2 */ (1'b0 & n2678) | ((1'b0 | n2678) & n2785);
assign n2796 = /* CARRY 20  7  3 */ (n2690 & n8) | ((n2690 | n8) & n3223);
assign n3198 = /* CARRY  2  8  0 */ (n66 & 1'b0) | ((n66 | 1'b0) & n5448);
assign n3199 = /* CARRY  4 19  2 */ (n8 & 1'b0) | ((n8 | 1'b0) & n789);
assign n2943 = /* CARRY 21  7  5 */ (n2692 & 1'b0) | ((n2692 | 1'b0) & n3143);
assign n3200 = /* CARRY  8 15  2 */ (n1026 & n914) | ((n1026 | n914) & n3144);
assign n3201 = /* CARRY 16 18  2 */ (1'b0 & n8) | ((1'b0 | n8) & n2416);
assign n3202 = /* CARRY  7 20  4 */ (1'b0 & n919) | ((1'b0 | n919) & n3225);
assign n2002 = /* CARRY 13 19  2 */ (n1553 & 1'b0) | ((n1553 | 1'b0) & n2001);
assign n3203 = /* CARRY  1  6  0 */ (n214 & n209) | ((n214 | n209) & n5504);
assign n2015 = /* CARRY 13 20  3 */ (n8 & n1649) | ((n8 | n1649) & n2014);
assign n3030 = /* CARRY 22 14  6 */ (n2969 & n8) | ((n2969 | n8) & n3029);
assign n2904 = /* CARRY 21  3  2 */ (n2762 & n8) | ((n2762 | n8) & n2903);
assign n1536 = /* CARRY 11  1  7 */ (1'b0 & n1529) | ((1'b0 | n1529) & n3149);
assign n3204 = /* CARRY  7 15  0 */ (n1028 & n922) | ((n1028 | n922) & n5563);
assign n1378 = /* CARRY  9 19  0 */ (1'b0 & n923) | ((1'b0 | n923) & n1372);
assign n3205 = /* CARRY  8  7  1 */ (n873 & n990) | ((n873 | n990) & n3228);
assign n2538 = /* CARRY 17 13  2 */ (1'b0 & n2385) | ((1'b0 | n2385) & n2537);
assign n1516 = /* CARRY 10 18  7 */ (n175 & 1'b0) | ((n175 | 1'b0) & n3151);
assign n3206 = /* CARRY 20  5  0 */ (1'b0 & n2675) | ((1'b0 | n2675) & n5591);
assign n3207 = /* CARRY  3 13  4 */ (1'b0 & n444) | ((1'b0 | n444) & n3153);
assign n3208 = /* CARRY 15 19  2 */ (1'b0 & n8) | ((1'b0 | n8) & n2288);
assign n801  = /* CARRY  4 21  5 */ (n620 & 1'b0) | ((n620 | 1'b0) & n800);
assign n3209 = /* CARRY  7 18  1 */ (n1053 & 1'b0) | ((n1053 | 1'b0) & n3155);
assign n3210 = /* CARRY  8 17  4 */ (1'b0 & n915) | ((1'b0 | n915) & n3156);
assign n3211 = /* CARRY  8  9  0 */ (n812 & 1'b0) | ((n812 | 1'b0) & n5651);
assign n3212 = /* CARRY  9 22  0 */ (1'b0 & n1019) | ((1'b0 | n1019) & n5656);
assign n3213 = /* CARRY 23  3  2 */ (1'b0 & n8) | ((1'b0 | n8) & n3048);
assign n3214 = /* CARRY 20  8  0 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2798);
assign n1850 = /* CARRY 12 22  1 */ (1'b0 & n1528) | ((1'b0 | n1528) & n3158);
assign n1372 = /* CARRY  9 18  7 */ (n8 & n821) | ((n8 | n821) & n3159);
assign n3215 = /* CARRY  3  8  0 */ (1'b0 & n66) | ((1'b0 | n66) & n5695);
assign n3216 = /* CARRY 11 11  0 */ (1'b0 & n1474) | ((1'b0 | n1474) & n5705);
assign n2148 = /* CARRY 14 19  1 */ (n1956 & n2009) | ((n1956 | n2009) & n2147);
assign n3217 = /* CARRY 15 18  4 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2282);
assign n3218 = /* CARRY 12  3  1 */ (n8 & n1533) | ((n8 | n1533) & n3161);
assign n2934 = /* CARRY 21  5  4 */ (n8 & n2780) | ((n8 | n2780) & n2933);
assign n2548 = /* CARRY 17 14  4 */ (n2265 & 1'b0) | ((n2265 | 1'b0) & n2547);
assign n3219 = /* CARRY 17  7  1 */ (1'b0 & n8) | ((1'b0 | n8) & n2485);
assign n3220 = /* CARRY  7 18  4 */ (n915 & 1'b0) | ((n915 | 1'b0) & n3237);
assign n1149 = /* CARRY  8  9  3 */ (1'b0 & n876) | ((1'b0 | n876) & n1148);
assign n3221 = /* CARRY  3 19  0 */ (1'b0 & n621) | ((1'b0 | n621) & n5757);
assign n3045 = /* CARRY 23  2  4 */ (n8 & n2899) | ((n8 | n2899) & n3163);
assign n3222 = /* CARRY 13 17  2 */ (1'b0 & n8) | ((1'b0 | n8) & n1988);
assign n3223 = /* CARRY 20  7  2 */ (1'b0 & n8) | ((1'b0 | n8) & n2795);
assign n2806 = /* CARRY 20  8  3 */ (n8 & n2803) | ((n8 | n2803) & n3240);
assign n1853 = /* CARRY 12 22  4 */ (n1848 & 1'b0) | ((n1848 | 1'b0) & n1852);
assign n3224 = /* CARRY 12 14  0 */ (n1622 & 1'b0) | ((n1622 | 1'b0) & n5784);
assign n2599 = /* CARRY 18  1  4 */ (1'b0 & n8) | ((1'b0 | n8) & n2598);
assign n1603 = /* CARRY 11 11  3 */ (n1329 & n8) | ((n1329 | n8) & n3241);
assign n2151 = /* CARRY 14 19  4 */ (1'b0 & n1984) | ((1'b0 | n1984) & n2150);
assign n2924 = /* CARRY 21  4  7 */ (n8 & n2671) | ((n8 | n2671) & n2923);
assign n1214 = /* CARRY  8 19  7 */ (n8 & n820) | ((n8 | n820) & n3169);
assign n3225 = /* CARRY  7 20  3 */ (1'b0 & n1047) | ((1'b0 | n1047) & n3170);
assign n2511 = /* CARRY 17 10  1 */ (n1766 & n1617) | ((n1766 | n1617) & n2510);
assign n1003 = /* CARRY  7  9  2 */ (n8 & n997) | ((n8 | n997) & n1002);
assign n2014 = /* CARRY 13 20  2 */ (n1553 & n8) | ((n1553 | n8) & n2013);
assign n634  = /* CARRY  3 19  3 */ (n334 & 1'b0) | ((n334 | 1'b0) & n633);
assign n2788 = /* CARRY 20  6  4 */ (1'b0 & n2680) | ((1'b0 | n2680) & n2787);
assign n2903 = /* CARRY 21  3  1 */ (n2894 & n8) | ((n2894 | n8) & n3174);
assign n412  = /* CARRY  2  8  2 */ (1'b0 & n226) | ((1'b0 | n226) & n411);
assign n3226 = /* CARRY 13  1  1 */ (n1402 & 1'b0) | ((n1402 | 1'b0) & n3249);
assign n2944 = /* CARRY 21  7  7 */ (1'b0 & n2691) | ((1'b0 | n2691) & n3175);
assign n3227 = /* CARRY  8 15  4 */ (n1025 & n915) | ((n1025 | n915) & n3177);
assign n3228 = /* CARRY  8  7  0 */ (n982 & n812) | ((n982 | n812) & n5907);
assign n2537 = /* CARRY 17 13  1 */ (n2386 & 1'b0) | ((n2386 | 1'b0) & n3178);
assign n3229 = /* CARRY 16 18  4 */ (1'b0 & n8) | ((1'b0 | n8) & n2417);
assign n3230 = /* CARRY  7 20  6 */ (n920 & 1'b0) | ((n920 | 1'b0) & n3253);
assign n2004 = /* CARRY 13 19  4 */ (n1715 & 1'b0) | ((n1715 | 1'b0) & n2003);
assign n3231 = /* CARRY  1  6  2 */ (1'b0 & n48) | ((1'b0 | n48) & n3255);
assign n3232 = /* CARRY 12  1  0 */ (n1531 & 1'b0) | ((n1531 | 1'b0) & n5972);
assign n2906 = /* CARRY 21  3  4 */ (n2764 & n8) | ((n2764 | n8) & n2905);
assign n3233 = /* CARRY 23 12  0 */ (n2500 & 1'b0) | ((n2500 | 1'b0) & n5996);
assign n3234 = /* CARRY  7 15  2 */ (n921 & n1026) | ((n921 | n1026) & n3258);
assign n2540 = /* CARRY 17 13  4 */ (1'b0 & n2255) | ((1'b0 | n2255) & n2539);
assign n491  = /* CARRY  2 21  1 */ (n324 & 1'b0) | ((n324 | 1'b0) & n3187);
assign n1974 = /* CARRY 13 15  1 */ (n1787 & n1969) | ((n1787 | n1969) & n3262);
assign n3235 = /* CARRY  3 13  6 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n590);
assign n3236 = /* CARRY 15 19  4 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n2289);
assign n2933 = /* CARRY 21  5  3 */ (n2779 & n8) | ((n2779 | n8) & n2932);
assign n803  = /* CARRY  4 21  7 */ (1'b0 & n334) | ((1'b0 | n334) & n802);
assign n778  = /* CARRY  4 18  1 */ (n8 & n630) | ((n8 | n630) & n3264);
assign n3237 = /* CARRY  7 18  3 */ (1'b0 & n918) | ((1'b0 | n918) & n3189);
assign n3238 = /* CARRY  8 17  6 */ (n8 & n913) | ((n8 | n913) & n3265);
assign n1148 = /* CARRY  8  9  2 */ (1'b0 & n878) | ((1'b0 | n878) & n1147);
assign n1393 = /* CARRY  9 22  2 */ (1'b0 & n1189) | ((1'b0 | n1189) & n1392);
assign n332  = /* CARRY  1 20  1 */ (n146 & 1'b0) | ((n146 | 1'b0) & n3268);
assign n3239 = /* CARRY 10 19  0 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n1516);
assign n3050 = /* CARRY 23  3  4 */ (n8 & n2887) | ((n8 | n2887) & n3049);
assign n3240 = /* CARRY 20  8  2 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2805);
assign n1852 = /* CARRY 12 22  3 */ (1'b0 & n1845) | ((1'b0 | n1845) & n1851);
assign n556  = /* CARRY  3  8  2 */ (n226 & 1'b0) | ((n226 | 1'b0) & n555);
assign n3241 = /* CARRY 11 11  2 */ (1'b0 & n8) | ((1'b0 | n8) & n1602);
assign n2150 = /* CARRY 14 19  3 */ (n1983 & n2008) | ((n1983 | n2008) & n2149);
assign n3242 = /* CARRY 15 15  1 */ (n2136 & n1765) | ((n2136 | n1765) & n3192);
assign n2923 = /* CARRY 21  4  6 */ (n8 & n2774) | ((n8 | n2774) & n2922);
assign n3243 = /* CARRY 15 18  6 */ (n8 & 1'b0) | ((n8 | 1'b0) & n2283);
assign n3244 = /* CARRY 12  3  3 */ (n8 & n1530) | ((n8 | n1530) & n3271);
assign n3245 = /* CARRY 17 19  0 */ (1'b0 & n2427) | ((1'b0 | n2427) & n6136);
assign n1002 = /* CARRY  7  9  1 */ (n8 & n996) | ((n8 | n996) & n3195);
assign n3246 = /* CARRY 17  7  3 */ (1'b0 & n8) | ((1'b0 | n8) & n2486);
assign n633  = /* CARRY  3 19  2 */ (n477 & 1'b0) | ((n477 | 1'b0) & n632);
assign n3046 = /* CARRY 23  2  6 */ (n8 & n2891) | ((n8 | n2891) & n3276);
assign n3247 = /* CARRY 13 17  4 */ (1'b0 & n8) | ((1'b0 | n8) & n1989);
assign n3248 = /* CARRY 20  7  4 */ (1'b0 & n8) | ((1'b0 | n8) & n2796);
assign n1794 = /* CARRY 12 14  2 */ (1'b0 & n1618) | ((1'b0 | n1618) & n1793);
assign n411  = /* CARRY  2  8  1 */ (1'b0 & n53) | ((1'b0 | n53) & n3198);
assign n3249 = /* CARRY 13  1  0 */ (1'b0 & n1531) | ((1'b0 | n1531) & n6196);
assign n790  = /* CARRY  4 19  3 */ (n8 & n488) | ((n8 | n488) & n3199);
assign n3250 = /* CARRY 18  6  0 */ (1'b0 & n2481) | ((1'b0 | n2481) & n6202);
assign n3251 = /* CARRY  4 12  0 */ (n271 & 1'b0) | ((n271 | 1'b0) & n6212);
assign n3252 = /* CARRY  4 13  1 */ (n8 & n424) | ((n8 | n424) & n3279);
assign n3253 = /* CARRY  7 20  5 */ (1'b0 & n909) | ((1'b0 | n909) & n3202);
assign n3254 = /* CARRY  9 16  0 */ (n922 & 1'b0) | ((n922 | 1'b0) & n6244);
assign n2003 = /* CARRY 13 19  3 */ (1'b0 & n1649) | ((1'b0 | n1649) & n2002);
assign n3255 = /* CARRY  1  6  1 */ (n49 & n208) | ((n49 | n208) & n3203);
assign n2016 = /* CARRY 13 20  4 */ (n8 & n1715) | ((n8 | n1715) & n2015);
assign n3256 = /* CARRY  2 19  0 */ (n323 & 1'b0) | ((n323 | 1'b0) & n6268);
assign n229  = /* CARRY  1  7  1 */ (n49 & n63) | ((n49 | n63) & n228);
assign n2905 = /* CARRY 21  3  3 */ (n2763 & n8) | ((n2763 | n8) & n2904);
assign n3257 = /* CARRY 13  1  3 */ (1'b0 & n1535) | ((1'b0 | n1535) & n3056);
assign n3258 = /* CARRY  7 15  1 */ (n910 & n1045) | ((n910 | n1045) & n3204);
assign n3259 = /* CARRY  8 15  6 */ (n1022 & n913) | ((n1022 | n913) & n3057);
assign n3260 = /* CARRY  8  7  2 */ (n987 & n862) | ((n987 | n862) & n3205);
assign n2539 = /* CARRY 17 13  3 */ (n2387 & 1'b0) | ((n2387 | 1'b0) & n2538);
assign n3261 = /* CARRY 16 18  6 */ (1'b0 & n8) | ((1'b0 | n8) & n2418);
assign n2473 = /* CARRY 17  6  0 */ (n2196 & n1541) | ((n2196 | n1541) & n6336);
assign n1382 = /* CARRY  9 20  1 */ (n1044 & n8) | ((n1044 | n8) & n3058);
assign n3262 = /* CARRY 13 15  0 */ (n1971 & 1'b0) | ((n1971 | 1'b0) & n6346);
assign n3263 = /* CARRY  3 14  1 */ (1'b0 & n444) | ((1'b0 | n444) & n3060);
assign n216  = /* CARRY  1  6  4 */ (1'b0 & n215) | ((1'b0 | n215) & n3061);
assign n3264 = /* CARRY  4 18  0 */ (1'b0 & n642) | ((1'b0 | n642) & n6375);
assign n3265 = /* CARRY  8 17  5 */ (n8 & n917) | ((n8 | n917) & n3210);
assign n3266 = /* CARRY 12  1  2 */ (n1533 & 1'b0) | ((n1533 | 1'b0) & n3062);
assign n3267 = /* CARRY  5 11  0 */ (n733 & 1'b0) | ((n733 | 1'b0) & n6398);
assign n1392 = /* CARRY  9 22  1 */ (n1050 & 1'b0) | ((n1050 | 1'b0) & n3212);
assign n2908 = /* CARRY 21  3  6 */ (n8 & n2766) | ((n8 | n2766) & n2907);
assign n3268 = /* CARRY  1 20  0 */ (1'b0 & n149) | ((1'b0 | n149) & n6409);
assign n336  = /* CARRY  1 21  1 */ (n152 & 1'b0) | ((n152 | 1'b0) & n3064);
assign n3269 = /* CARRY  7 15  4 */ (n919 & n1025) | ((n919 | n1025) & n3065);
assign n616  = /* CARRY  3 17  1 */ (1'b0 & n614) | ((1'b0 | n614) & n3068);
assign n1976 = /* CARRY 13 15  3 */ (n1802 & n1801) | ((n1802 | n1801) & n1975);
assign n3270 = /* CARRY 22 14  0 */ (1'b0 & n2976) | ((1'b0 | n2976) & n6450);
assign n3271 = /* CARRY 12  3  2 */ (n1535 & n8) | ((n1535 | n8) & n3218);
assign n3272 = /* CARRY  2  6  0 */ (1'b0 & n6) | ((1'b0 | n6) & n6465);
assign n2935 = /* CARRY 21  5  5 */ (n2929 & n8) | ((n2929 | n8) & n2934);
assign n779  = /* CARRY  4 18  3 */ (n777 & n8) | ((n777 | n8) & n3070);
assign n3273 = /* CARRY 11  1  1 */ (1'b0 & n1402) | ((1'b0 | n1402) & n3071);
assign n3274 = /* CARRY  7 18  5 */ (1'b0 & n917) | ((1'b0 | n917) & n3220);
assign n2486 = /* CARRY 17  7  2 */ (n1868 & 1'b0) | ((n1868 | 1'b0) & n3219);
assign n1150 = /* CARRY  8  9  4 */ (n989 & 1'b0) | ((n989 | 1'b0) & n1149);
assign n3275 = /* CARRY 10 18  1 */ (1'b0 & n189) | ((1'b0 | n189) & n3072);
assign n1395 = /* CARRY  9 22  4 */ (n907 & 1'b0) | ((n907 | 1'b0) & n1394);
assign n3276 = /* CARRY 23  2  5 */ (1'b0 & n8) | ((1'b0 | n8) & n3045);
assign n1989 = /* CARRY 13 17  3 */ (1'b0 & n1812) | ((1'b0 | n1812) & n3222);
assign n3277 = /* CARRY 20  8  4 */ (1'b0 & 1'b0) | ((1'b0 | 1'b0) & n2806);
assign n1854 = /* CARRY 12 22  5 */ (n1847 & 1'b0) | ((n1847 | 1'b0) & n1853);
assign n1793 = /* CARRY 12 14  1 */ (1'b0 & n1617) | ((1'b0 | n1617) & n3224);
assign n3278 = /* CARRY  2 17  0 */ (n316 & 1'b0) | ((n316 | 1'b0) & n6533);
assign n2759 = /* CARRY 20  1  1 */ (1'b0 & n2595) | ((1'b0 | n2595) & n3074);
assign n3279 = /* CARRY  4 13  0 */ (1'b0 & n430) | ((1'b0 | n430) & n6557);
assign n1070 = /* CARRY  7 21  0 */ (1'b0 & n911) | ((1'b0 | n911) & n1065);
assign n3280 = /* CARRY 12  3  5 */ (n1534 & 1'b0) | ((n1534 | 1'b0) & n3075);
assign n3281 = /* CARRY 17 19  2 */ (1'b0 & n8) | ((1'b0 | n8) & n2577);
assign n1371 = /* CARRY  9 17  0 */ (1'b0 & n911) | ((1'b0 | n911) & n1368);
assign n1004 = /* CARRY  7  9  3 */ (n998 & n8) | ((n998 | n8) & n1003);
assign n228  = /* CARRY  1  7  0 */ (n214 & n60) | ((n214 | n60) & n6606);
assign n635  = /* CARRY  3 19  4 */ (n488 & 1'b0) | ((n488 | 1'b0) & n634);
assign n2789 = /* CARRY 20  6  5 */ (1'b0 & n2681) | ((1'b0 | n2681) & n2788);
assign n3282 = /* CARRY 13 17  6 */ (1'b0 & n8) | ((1'b0 | n8) & n1990);
assign n3283 = /* CARRY  1  8  1 */ (n231 & n46) | ((n231 | n46) & n3079);
assign n3284 = /* CARRY 20  7  6 */ (1'b0 & n8) | ((1'b0 | n8) & n2797);
/* FF 13  1  2 */ assign n3285 = n3286;
/* FF  2  8  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n227 <= 1'b0; else if (n70) n227 <= n3287;
/* FF  4 19  5 */ assign n627 = n3288;
/* FF 14 22  5 */ assign n2025 = n3289;
/* FF 14 14  1 */ assign n1960 = n3290;
/* FF  3  7  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n44 <= 1'b0; else if (n224) n44 <= n3291;
/* FF 11 10  7 */ always @(posedge io_13_31_1) if (n4) n1462 <= 1'b0 ? 1'b0 : n3292;
/* FF 12  6  5 */ assign n1561 = n3293;
/* FF 15 13  4 */ assign n2102 = n3294;
/* FF  5 16  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n764 <= 1'b0; else if (n80) n764 <= n3295;
/* FF  4 20  6 */ assign n489 = n3296;
/* FF  4 12  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n579 <= 1'b0; else if (n432) n579 <= n3297;
/* FF 14 15  2 */ assign n1779 = n3298;
/* FF  8 16  1 */ assign n1049 = n3299;
/* FF  2  4  5 */ assign n196 = n3300;
/* FF 22  4  6 */ assign n2914 = n3301;
/* FF 14 18  7 */ always @(posedge io_13_31_1) if (n1513) n1997 <= n1 ? 1'b0 : n3302;
/* FF 11  2  2 */ assign n1399 = n3303;
/* FF  8 15  5 */ assign n3304 = n3305;
/* FF 15 14  5 */ assign n2104 = n3306;
/* FF 15  6  1 */ assign n2055 = n3307;
/* FF  5  9  0 */ always @(posedge io_13_31_1) if (n4) n714 <= 1'b0 ? 1'b0 : n3308;
/* FF 24 13  4 */ always @(posedge io_13_31_1) if (1'b1) n3052 <= n2395 ? 1'b0 : n3309;
/* FF 12  2  7 */ assign n1535 = n3310;
/* FF  5  8  4 */ always @(posedge io_13_31_1) if (n4) n706 <= 1'b0 ? 1'b0 : n3311;
/* FF 16 19  1 */ assign n3312 = n3313;
/* FF  4  4  3 */ assign n522 = n3314;
/* FF 11  3  3 */ assign n956 = n3315;
/* FF 16 18  5 */ assign n3316 = n3317;
/* FF  1 18  0 */ assign n130 = n3318;
/* FF 20 22  4 */ assign n2594 = n3319;
/* FF  9 20  0 */ assign n3320 = n3321;
/* FF  5  1  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n650 <= 1'b0; else if (n656) n650 <= n3323;
/* FF  7 20  7 */ assign n3324 = n3325;
/* FF 17  9  4 */ assign n2360 = n3326;
/* FF  7 12  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n887 <= 1'b0; else if (n818) n887 <= n3327;
/* FF  8  8  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n876 <= 1'b0; else if (n877) n876 <= n3328;
/* FF  5  4  6 */ assign n676 = n3329;
/* FF 16 11  2 */ always @(posedge io_13_31_1) if (n2076) n2231 <= 1'b0 ? 1'b0 : n3330;
/* FF 16 14  7 */ assign n1766 = n3331;
/* FF 17 10  5 */ assign n2369 = n3332;
/* FF  7 13  4 */ assign n898 = n3333;
/* FF 17  2  1 */ always @(posedge io_13_31_1) if (n2324) n2306 <= 1'b0 ? 1'b0 : n3334;
/* FF  7  5  0 */ assign n699 = n3335;
/* FF  5  5  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n680 <= 1'b0; else if (n524) n680 <= n3336;
/* FF  9 16  2 */ assign n3337 = n3338;
/* FF  4  1  6 */ assign n498 = n3339;
/* FF 14  3  4 */ assign n1872 = n3340;
/* FF  8  4  3 */ assign n656 = n3341;
/* FF 16  7  4 */ assign n2200 = n3342;
/* FF 13 19  5 */ assign n1820 = n3343;
/* FF 20 18  5 */ assign n2732 = n3344;
/* FF  3 14  0 */ assign n3345 = n3346;
/* FF  1 14  7 */ assign n111 = n3348;
/* FF  1  6  3 */ assign n3349 = n3350;
/* FF 10 12  4 */ assign n1324 = n3351;
/* FF  9  8  3 */ always @(posedge io_13_31_1) if (n4) n1130 <= 1'b0 ? 1'b0 : n3352;
/* FF 13 20  6 */ assign n1825 = n3353;
/* FF  2 18  1 */ assign n310 = n3354;
/* FF 21 22  5 */ assign n2881 = n3355;
/* FF 11 17  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1469 <= 1'b0; else if (n762) n1469 <= n3356;
/* FF 18 16  0 */ always @(posedge io_13_31_1) if (n2011) n2551 <= 1'b0 ? 1'b0 : n3357;
/* FF  3 18  6 */ assign n463 = n3358;
/* FF 10  5  1 */ assign n1264 = n3359;
/* FF  9  1  0 */ assign n1076 = n3360;
/* FF  2 19  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n320 <= 1'b0; else if (n322) n320 <= n3361;
/* FF  7  1  7 */ assign n828 = n3362;
/* FF  3 15  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n438 <= 1'b0; else if (1'b1) n438 <= n3363;
/* FF 11 18  1 */ always @(posedge io_13_31_1) if (1'b1) n1504 <= 1'b0 ? 1'b0 : n3364;
/* FF 11 21  6 */ assign n1525 = n3365;
/* FF 12 17  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1171 <= 1'b0; else if (1'b1) n1171 <= n3366;
/* FF 12  9  0 */ assign n1583 = n3367;
/* FF  3 10  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n63 <= 1'b0; else if (n576) n63 <= n3368;
/* FF 22 12  0 */ always @(posedge io_13_31_1) if (n2137) n2956 <= n3 ? 1'b0 : n3369;
/* FF  3  2  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n349 <= 1'b0; else if (n500) n349 <= n3370;
/* FF 18 11  6 */ always @(posedge io_13_31_1) if (n2137) n2518 <= n3 ? 1'b0 : n3371;
/* FF 15 16  5 */ assign n2136 = n3372;
/* FF  8 18  0 */ assign n3373 = n3374;
/* FF 11 13  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1465 <= 1'b0; else if (n1461) n1465 <= n3375;
/* FF 18 12  7 */ assign n2390 = n3376;
/* FF 11  5  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1418 <= 1'b0; else if (n1279) n1418 <= n3377;
/* FF 18  4  3 */ always @(posedge io_13_31_1) if (n2603) n2453 <= 1'b0 ? 1'b0 : n3378;
/* FF 12  1  1 */ assign n3379 = n3380;
/* FF  5 19  3 */ assign n784 = n3381;
/* FF  4 15  2 */ assign n602 = n3382;
/* FF 12  4  6 */ assign n1349 = n3383;
/* FF  8 19  1 */ assign n3384 = n3385;
/* FF  2  7  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n221 <= 1'b0; else if (n224) n221 <= n3386;
/* FF 22  7  6 */ always @(posedge io_13_31_1) if (n2694) n2692 <= n1 ? 1'b0 : n3387;
/* FF  3  3  3 */ assign n358 = n3388;
/* FF 21  3  5 */ always @(posedge io_13_31_1) if (n2902) n2765 <= n7 ? 1'b0 : n3389;
/* FF 14 21  7 */ assign n1981 = n3390;
/* FF 11  6  4 */ assign n1122 = n3391;
/* FF 15 17  5 */ assign n2134 = n3392;
/* FF 15  9  1 */ assign n2078 = n3393;
/* FF  5 12  0 */ always @(posedge io_13_31_1) if (n4) n738 <= 1'b0 ? 1'b0 : n3394;
/* FF 17 21  5 */ assign n2296 = n3395;
/* FF 12  5  7 */ assign n1552 = n3396;
/* FF 14 14  4 */ assign n1961 = n3397;
/* FF 14  6  0 */ assign n1894 = n3398;
/* FF  1 21  0 */ assign n3399 = n3400;
/* FF 23 12  1 */ always @(posedge io_13_31_1) if (n2826) n2809 <= n2957 ? 1'b0 : n3402;
/* FF  8 14  7 */ assign n1042 = n3403;
/* FF 20 17  0 */ assign n2724 = n3404;
/* FF  7 15  3 */ assign n3405 = n3406;
/* FF  5  7  6 */ assign n696 = n3407;
/* FF  9 19  3 */ assign n1210 = n3408;
/* FF  4  3  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n515 <= 1'b0; else if (n509) n515 <= n3409;
/* FF  8  7  4 */ assign n3410 = n3411;
/* FF 16  9  3 */ assign n2217 = n3412;
/* FF 20 21  6 */ assign n2590 = n3413;
/* FF 17 13  5 */ always @(posedge io_13_31_1) if (n2536) n2256 <= n1 ? 1'b0 : n3414;
/* FF 17  5  1 */ always @(posedge io_13_31_1) if (n2456) n2335 <= 1'b0 ? 1'b0 : n3415;
/* FF 20 13  2 */ always @(posedge io_13_31_1) if (n2663) n2708 <= 1'b0 ? 1'b0 : n3416;
/* FF  7  8  0 */ assign n3417 = n3418;
/* FF  5  8  7 */ always @(posedge io_13_31_1) if (n4) n709 <= 1'b0 ? 1'b0 : n3420;
/* FF 18 18  0 */ always @(posedge io_13_31_1) if (n2563) n2561 <= 1'b0 ? 1'b0 : n3421;
/* FF  4  4  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n381 <= 1'b0; else if (n198) n381 <= n3422;
/* FF  7 11  5 */ always @(posedge io_13_31_1) if (n4) n884 <= 1'b0 ? 1'b0 : n3423;
/* FF 13 23  1 */ assign n1855 = n3424;
/* FF 16 10  4 */ assign n2225 = n3425;
/* FF 13 22  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1846 <= 1'b0; else if (n1666) n1846 <= n3426;
/* FF 17  6  2 */ assign n3427 = n3428;
/* FF 14  2  7 */ assign n1867 = n3429;
/* FF  3 17  0 */ assign n3430 = n3431;
/* FF 10 16  0 */ always @(posedge io_13_31_1) if (n4) n1361 <= 1'b0 ? 1'b0 : n3433;
/* FF  1 17  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n126 <= 1'b0; else if (n118) n126 <= n3434;
/* FF 17  9  7 */ assign n2362 = n3435;
/* FF  1  9  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n66 <= 1'b0; else if (n70) n66 <= n3436;
/* FF  7  4  2 */ assign n842 = n3437;
/* FF  9 11  3 */ assign n1161 = n3438;
/* FF 16  3  1 */ assign n1529 = n3439;
/* FF 13 15  2 */ assign n1796 = n3440;
/* FF  7  3  6 */ assign n838 = n3441;
/* FF 10 11  7 */ always @(posedge io_13_31_1) if (n4) n1317 <= 1'b0 ? 1'b0 : n3442;
/* FF 13 18  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1650 <= 1'b0; else if (n1967) n1650 <= n3443;
/* FF  3 21  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n486 <= 1'b0; else if (1'b1) n486 <= n3444;
/* FF 10  8  1 */ assign n1283 = n3445;
/* FF 22 22  3 */ assign n3003 = n3446;
/* FF  9  7  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n208 <= 1'b0; else if (n877) n208 <= n3447;
/* FF 13 11  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1751 <= 1'b0; else if (n734) n1751 <= n3448;
/* FF 21 21  7 */ assign n2875 = n3449;
/* FF  3 14  3 */ assign n436 = n3450;
/* FF 11 16  2 */ always @(posedge io_13_31_1) if (n4) n1498 <= 1'b0 ? 1'b0 : n3451;
/* FF 12 12  0 */ assign n3452 = n3453;
/* FF 22 15  0 */ assign n3455 = n3456;
/* FF  3 13  7 */ assign n433 = n3457;
/* FF 10 12  7 */ assign n1327 = n3458;
/* FF 10  4  3 */ assign n1260 = n3459;
/* FF  9  8  6 */ always @(posedge io_13_31_1) if (n4) n1133 <= 1'b0 ? 1'b0 : n3460;
/* FF  2 18  4 */ assign n313 = n3461;
/* FF 21 14  4 */ always @(posedge io_13_31_1) if (n2842) n2833 <= 1'b0 ? 1'b0 : n3462;
/* FF 11 17  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1359 <= 1'b0; else if (n762) n1359 <= n3463;
/* FF  8 21  0 */ assign n1066 = n3464;
/* FF 13  3  5 */ assign n840 = n3465;
/* FF 18  7  3 */ always @(posedge io_13_31_1) if (n2076) n2479 <= 1'b0 ? 1'b0 : n3466;
/* FF 15 20  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1649 <= 1'b0; else if (n1815) n1649 <= n3467;
/* FF 15 12  2 */ assign n1778 = n3468;
/* FF  4 18  2 */ assign n617 = n3469;
/* FF  2 10  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n199 <= 1'b0; else if (1'b1) n199 <= n3470;
/* FF  5 18  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n630 <= 1'b0; else if (n474) n630 <= n3471;
/* FF  2  2  1 */ assign n168 = n3472;
/* FF 21  6  5 */ always @(posedge io_13_31_1) if (n2686) n2194 <= 1'b0 ? 1'b0 : n3473;
/* FF 14 16  3 */ assign n1979 = n3474;
/* FF 11  1  0 */ assign n3475 = n3476;
/* FF  5 15  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n757 <= 1'b0; else if (n451) n757 <= n3478;
/* FF  3  2  6 */ assign n352 = n3479;
/* FF 23 15  2 */ assign n3032 = n3480;
/* FF 11  4  5 */ assign n1413 = n3481;
/* FF 12  8  7 */ assign n1582 = n3482;
/* FF  2  3  2 */ assign n182 = n3483;
/* FF 24 14  5 */ always @(posedge io_13_31_1) if (n2819) n2818 <= n2841 ? 1'b1 : n3484;
/* FF  4 14  4 */ assign n588 = n3485;
/* FF 14  9  0 */ assign n1913 = n3486;
/* FF 11  5  6 */ assign n983 = n3487;
/* FF  8 17  7 */ assign n3488 = n3489;
/* FF 17  8  2 */ assign n2349 = n3490;
/* FF 10 18  0 */ assign n3491 = n3492;
/* FF  9 22  3 */ assign n1230 = n3494;
/* FF 17 11  7 */ assign n2378 = n3495;
/* FF  4  6  5 */ assign n539 = n3496;
/* FF  7 14  6 */ assign n906 = n3497;
/* FF  8 10  4 */ always @(posedge io_13_31_1) if (n4) n1009 <= 1'b0 ? 1'b0 : n3498;
/* FF  8  2  0 */ assign n518 = n3499;
/* FF  1 20  2 */ assign n144 = n3500;
/* FF 14  4  6 */ assign n1565 = n3501;
/* FF 10 19  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n277 <= 1'b0; else if (1'b1) n277 <= n3502;
/* FF  5  3  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n380 <= 1'b0; else if (n198) n380 <= n3503;
/* FF 23  3  5 */ always @(posedge io_13_31_1) if (1'b1) n3010 <= n2888 ? 1'b0 : n3504;
/* FF  9 15  0 */ assign n1190 = n3505;
/* FF 17  4  4 */ always @(posedge io_13_31_1) if (n2316) n2329 <= 1'b0 ? 1'b0 : n3506;
/* FF  8  3  1 */ assign n949 = n3507;
/* FF 16 13  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1938 <= 1'b0; else if (n735) n1938 <= n3508;
/* FF  4  2  7 */ assign n508 = n3509;
/* FF 16  5  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1914 <= 1'b0; else if (n1869) n1914 <= n3510;
/* FF 14  5  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1889 <= 1'b0; else if (n1433) n1889 <= n3511;
/* FF 18 22  1 */ assign n2587 = n3512;
/* FF  1 12  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) io_4_31_0 <= 1'b1; else if (1'b1) io_4_31_0 <= n3513;
/* FF  7 15  6 */ assign n3514 = n3515;
/* FF  7  7  2 */ assign n855 = n3516;
/* FF 16  6  1 */ assign n2185 = n3517;
/* FF 10 14  7 */ always @(posedge io_13_31_1) if (n4) n1348 <= 1'b0 ? 1'b0 : n3518;
/* FF  9 10  6 */ always @(posedge io_13_31_1) if (n4) n1157 <= 1'b0 ? 1'b0 : n3519;
/* FF 16  9  6 */ assign n2219 = n3520;
/* FF  1  5  0 */ always @(posedge io_13_31_1) if (n201) n36 <= n42 ? 1'b0 : n3521;
/* FF  3 16  2 */ assign n447 = n3522;
/* FF 20  1  0 */ assign n3523 = n3524;
/* FF 12 15  1 */ always @(posedge io_13_31_1) if (n1180) n1629 <= n1 ? 1'b0 : n3526;
/* FF 20  4  5 */ assign n2603 = n3527;
/* FF 13 14  4 */ assign n1786 = n3528;
/* FF 22 13  2 */ always @(posedge io_13_31_1) if (n2663) n2959 <= 1'b0 ? 1'b0 : n3529;
/* FF  3 17  3 */ assign n453 = n3530;
/* FF  1  9  6 */ assign n68 = n3531;
/* FF 15 23  1 */ always @(posedge io_13_31_1) if (n2157) n2159 <= 1'b0 ? 1'b0 : n3532;
/* FF 20  5  6 */ assign n2363 = n3533;
/* FF  9 11  6 */ assign n1164 = n3534;
/* FF 12 19  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1648 <= 1'b0; else if (n1815) n1648 <= n3535;
/* FF 18 10  4 */ always @(posedge io_13_31_1) if (n2120) n2374 <= 1'b0 ? 1'b0 : n3536;
/* FF  9  3  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1095 <= 1'b0; else if (n851) n1095 <= n3537;
/* FF 12 11  3 */ assign n1564 = n3538;
/* FF 18  2  0 */ always @(posedge io_13_31_1) if (n2456) n2443 <= 1'b0 ? 1'b0 : n3539;
/* FF 13  7  1 */ always @(posedge io_13_31_1) if (n4) n1167 <= 1'b0 ? 1'b0 : n3540;
/* FF 21 17  4 */ assign n2850 = n3541;
/* FF 11 20  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1520 <= 1'b0; else if (n1515) n1520 <= n3542;
/* FF  2 13  6 */ assign n275 = n3543;
/* FF 13  6  5 */ assign n1712 = n3544;
/* FF  3  1  0 */ assign n338 = n3545;
/* FF 22 14  2 */ always @(posedge io_13_31_1) if (1'b1) n2966 <= n3025 ? 1'b0 : n3546;
/* FF 15 15  2 */ assign n3547 = n3548;
/* FF  3  4  5 */ assign n368 = n3549;
/* FF 15 18  7 */ assign n3550 = n3551;
/* FF 12  3  4 */ assign n3552 = n3553;
/* FF  5 13  2 */ assign n578 = n3554;
/* FF  4 17  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n316 <= 1'b1; else if (n317) n316 <= n3555;
/* FF  4  9  1 */ always @(posedge io_13_31_1) if (n4) n557 <= 1'b0 ? 1'b0 : n3556;
/* FF  3  5  6 */ assign n379 = n3557;
/* FF 16 23  3 */ always @(posedge io_13_31_1) if (n2300) n2299 <= 1'b0 ? 1'b0 : n3558;
/* FF 17 19  1 */ assign n3559 = n3560;
/* FF 11  7  5 */ assign n1432 = n3561;
/* FF 15 11  4 */ assign n2098 = n3562;
/* FF  2  6  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n176 <= 1'b0; else if (n217) n176 <= n3563;
/* FF  5 14  3 */ assign n754 = n3564;
/* FF 14 20  4 */ always @(posedge io_13_31_1) if (n1838) n2009 <= n2155 ? 1'b0 : n3565;
/* FF  8 21  3 */ assign n1068 = n3566;
/* FF 14 12  0 */ assign n1941 = n3567;
/* FF 21  5  7 */ assign n2783 = n3568;
/* FF 17 20  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2156 <= 1'b0; else if (n2023) n2156 <= n3569;
/* FF 11  8  6 */ always @(posedge io_13_31_1) if (n4) n1441 <= 1'b0 ? 1'b0 : n3570;
/* FF 15 12  5 */ assign n2108 = n3571;
/* FF 15  4  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1904 <= 1'b0; else if (n1547) n1904 <= n3572;
/* FF 23 14  4 */ always @(posedge io_13_31_1) if (1'b1) n3022 <= 1'b0 ? 1'b0 : n3573;
/* FF  4 10  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n573 <= 1'b0; else if (n576) n573 <= n3574;
/* FF 14 13  1 */ assign n1949 = n3575;
/* FF 22  2  5 */ always @(posedge io_13_31_1) if (1'b1) n2891 <= 1'b0 ? 1'b0 : n3576;
/* FF  2  2  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n171 <= 1'b0; else if (n178) n171 <= n3577;
/* FF 16 24  3 */ assign n2301 = n3578;
/* FF  7 17  6 */ assign n917 = n3579;
/* FF 14 16  6 */ assign n1973 = n3580;
/* FF 11  1  3 */ assign n3581 = n3582;
/* FF  8 13  4 */ assign n1027 = n3583;
/* FF  8  5  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n968 <= 1'b0; else if (n663) n968 <= n3584;
/* FF 23  7  1 */ always @(posedge io_13_31_1) if (n2676) n2621 <= n1 ? 1'b0 : n3585;
/* FF  9 18  0 */ assign n3586 = n3587;
/* FF  7 18  7 */ assign n3589 = n3590;
/* FF 17  7  4 */ assign n3591 = n3592;
/* FF  7 10  3 */ always @(posedge io_13_31_1) if (n4) n879 <= 1'b0 ? 1'b0 : n3593;
/* FF  9 21  5 */ assign n1224 = n3594;
/* FF  8  6  1 */ assign n977 = n3595;
/* FF 16  8  0 */ assign n2205 = n3596;
/* FF 20 20  3 */ assign n2743 = n3597;
/* FF 14  8  7 */ assign n1922 = n3598;
/* FF  8  9  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1000 <= 1'b0; else if (n877) n1000 <= n3599;
/* FF 17  8  5 */ always @(posedge io_13_31_1) if (n2344) n2352 <= 1'b0 ? 1'b0 : n3600;
/* FF 10 18  3 */ assign n3601 = n3602;
/* FF  9 22  6 */ assign n1232 = n3603;
/* FF  5  2  5 */ assign n661 = n3604;
/* FF 23  2  7 */ assign n3008 = n3605;
/* FF  9 14  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1144 <= 1'b0; else if (n762) n1144 <= n3606;
/* FF 16 12  6 */ assign n2237 = n3607;
/* FF 16  4  2 */ always @(posedge io_13_31_1) if (n2324) n2174 <= 1'b0 ? 1'b0 : n3608;
/* FF  1  8  0 */ assign n3609 = n3610;
/* FF 13 17  5 */ assign n3612 = n3613;
/* FF  8  1  7 */ assign n940 = n3614;
/* FF 12 18  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1641 <= 1'b0; else if (1'b1) n1641 <= n3615;
/* FF 20  7  5 */ assign n3616 = n3617;
/* FF 10 10  4 */ always @(posedge io_13_31_1) if (n4) n1306 <= 1'b0 ? 1'b0 : n3618;
/* FF 10  2  0 */ assign n1244 = n3619;
/* FF  9  6  3 */ assign n1118 = n3620;
/* FF 22 16  2 */ assign n2978 = n3621;
/* FF 13  9  0 */ assign n1742 = n3622;
/* FF  2 16  1 */ assign n293 = n3623;
/* FF  3 20  3 */ assign n479 = n3624;
/* FF 21 20  5 */ assign n2865 = n3625;
/* FF 21 12  1 */ always @(posedge io_13_31_1) if (n2663) n2812 <= 1'b0 ? 1'b0 : n3626;
/* FF  1 12  6 */ assign n88 = n3627;
/* FF  1  4  2 */ always @(posedge io_13_31_1) if (n201) n29 <= n42 ? 1'b0 : n3628;
/* FF 20  8  6 */ always @(posedge io_13_31_1) if (1'b1) n15 <= 1'b0 ? 1'b0 : n3629;
/* FF 12 22  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1665 <= 1'b0; else if (n1666) n1665 <= n3630;
/* FF 18 13  4 */ always @(posedge io_13_31_1) if (n2137) n2532 <= n3 ? 1'b0 : n3631;
/* FF 12 14  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1619 <= 1'b0; else if (n1630) n1619 <= n3632;
/* FF 18  5  0 */ assign n2457 = n3633;
/* FF 22 17  3 */ assign n2736 = n3634;
/* FF  2 17  2 */ assign n299 = n3635;
/* FF 13 10  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1730 <= 1'b0; else if (n734) n1730 <= n3636;
/* FF  9  2  5 */ assign n1088 = n3637;
/* FF 14 23  0 */ assign n3638 = n3639;
/* FF 21 16  7 */ always @(posedge io_13_31_1) if (n2852) n2847 <= 1'b0 ? 1'b0 : n3641;
/* FF 20  1  3 */ always @(posedge io_13_31_1) if (n2600) n2448 <= n2758 ? 1'b0 : n3642;
/* FF 10  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1253 <= 1'b0; else if (n851) n1253 <= n3643;
/* FF 18  6  1 */ always @(posedge io_13_31_1) if (n2602) n2465 <= n1 ? 1'b0 : n3644;
/* FF 12  7  0 */ assign n1567 = n3645;
/* FF 21 13  1 */ assign n3646 = n3647;
/* FF 18  9  6 */ assign n2497 = n3648;
/* FF 12  6  4 */ assign n1560 = n3649;
/* FF  5 16  2 */ assign n763 = n3650;
/* FF 11 19  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1477 <= 1'b1; else if (1'b1) n1477 <= n3651;
/* FF  4 20  5 */ assign n639 = n3652;
/* FF  4 12  1 */ assign n3653 = n3654;
/* FF 13  5  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1698 <= 1'b0; else if (n1279) n1698 <= n3655;
/* FF 14 15  1 */ assign n1969 = n3656;
/* FF  8 16  0 */ assign n3657 = n3658;
/* FF  2  4  4 */ always @(posedge io_13_31_1) if (n201) n195 <= n42 ? 1'b0 : n3659;
/* FF  3  8  6 */ assign n408 = n3660;
/* FF 17 22  1 */ always @(posedge io_13_31_1) if (n2160) n2433 <= 1'b0 ? 1'b0 : n3661;
/* FF 18  2  3 */ always @(posedge io_13_31_1) if (n2456) n2445 <= 1'b0 ? 1'b0 : n3662;
/* FF  5 17  3 */ assign n770 = n3663;
/* FF 15  6  0 */ always @(posedge io_13_31_1) if (n2191) n1416 <= 1'b0 ? 1'b0 : n3664;
/* FF  4 13  2 */ assign n3665 = n3666;
/* FF 12  2  6 */ assign n1533 = n3667;
/* FF  2  5  5 */ assign n206 = n3668;
/* FF 16 19  0 */ assign n2285 = n3669;
/* FF  4 16  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n605 <= 1'b0; else if (1'b1) n605 <= n3670;
/* FF  3  1  3 */ assign n341 = n3671;
/* FF 11 11  6 */ assign n1179 = n3672;
/* FF 11  3  2 */ assign n1404 = n3673;
/* FF 15 15  5 */ assign n2130 = n3674;
/* FF 14 11  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1891 <= 1'b0; else if (n734) n1891 <= n3675;
/* FF 14 19  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1966 <= 1'b0; else if (n1527) n1966 <= n3676;
/* FF 15  7  1 */ assign n2059 = n3677;
/* FF  5 10  0 */ always @(posedge io_13_31_1) if (n4) n723 <= 1'b0 ? 1'b0 : n3678;
/* FF  7 21  2 */ assign n925 = n3679;
/* FF 12  3  7 */ assign n1540 = n3680;
/* FF 22  5  5 */ always @(posedge io_13_31_1) if (n2456) n2617 <= 1'b0 ? 1'b0 : n3681;
/* FF  5 13  5 */ always @(posedge io_13_31_1) if (n4) n746 <= 1'b0 ? 1'b0 : n3682;
/* FF  4  9  4 */ always @(posedge io_13_31_1) if (n4) n560 <= 1'b0 ? 1'b0 : n3683;
/* FF  8  8  0 */ assign n987 = n3684;
/* FF 17 11  0 */ assign n3685 = n3686;
/* FF 17 10  4 */ assign n2368 = n3688;
/* FF  7 13  3 */ always @(posedge io_13_31_1) if (n4) n897 <= 1'b0 ? 1'b0 : n3689;
/* FF 15  2  7 */ assign n2048 = n3690;
/* FF  5  5  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n678 <= 1'b0; else if (n524) n678 <= n3691;
/* FF  9 16  1 */ assign n3692 = n3693;
/* FF  4  1  5 */ assign n497 = n3694;
/* FF 14  3  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1703 <= 1'b0; else if (n1690) n1703 <= n3695;
/* FF  8  4  2 */ assign n963 = n3696;
/* FF 16 15  7 */ always @(posedge io_13_31_1) if (n2268) n2264 <= 1'b0 ? 1'b0 : n3697;
/* FF 20 18  4 */ assign n2731 = n3698;
/* FF 17  3  1 */ assign n2318 = n3699;
/* FF  7  6  0 */ assign n532 = n3700;
/* FF  9 17  2 */ always @(posedge io_13_31_1) if (1'b1) n1200 <= 1'b0 ? 1'b0 : n3701;
/* FF  7  9  5 */ assign n874 = n3702;
/* FF  8  5  3 */ assign n663 = n3703;
/* FF 13 20  5 */ assign n1826 = n3704;
/* FF 20 11  1 */ always @(posedge io_13_31_1) if (n2137) n2696 <= n3 ? 1'b0 : n3705;
/* FF 10 14  0 */ always @(posedge io_13_31_1) if (n4) n1341 <= 1'b0 ? 1'b0 : n3706;
/* FF 18 24  3 */ always @(posedge io_13_31_1) if (n2591) n2567 <= 1'b0 ? 1'b0 : n3707;
/* FF 17  7  7 */ assign n2344 = n3708;
/* FF  3 18  5 */ assign n462 = n3709;
/* FF 16  8  3 */ assign n2208 = n3710;
/* FF  2 19  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n319 <= 1'b0; else if (n322) n319 <= n3711;
/* FF  7  1  6 */ assign n827 = n3712;
/* FF 13 13  2 */ assign n1772 = n3713;
/* FF 18 17  0 */ always @(posedge io_13_31_1) if (n2559) n2557 <= 1'b0 ? 1'b0 : n3714;
/* FF  1  7  2 */ assign n47 = n3715;
/* FF 13 16  7 */ assign n1801 = n3716;
/* FF  3 19  6 */ assign n472 = n3717;
/* FF 20  3  2 */ always @(posedge io_13_31_1) if (1'b1) n233 <= 1'b0 ? 1'b0 : n3718;
/* FF 11 21  5 */ assign n1524 = n3719;
/* FF 12 17  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1495 <= 1'b0; else if (1'b1) n1495 <= n3720;
/* FF 20  6  7 */ assign n2602 = n3721;
/* FF  2 20  2 */ assign n328 = n3722;
/* FF 10  9  6 */ always @(posedge io_13_31_1) if (n4) n1299 <= 1'b0 ? 1'b0 : n3723;
/* FF  9  5  5 */ assign n1112 = n3724;
/* FF  1  8  3 */ assign n54 = n3725;
/* FF 21 19  7 */ assign n2861 = n3726;
/* FF  3 11  1 */ assign n424 = n3727;
/* FF 11 14  2 */ assign n762 = n3728;
/* FF 12 18  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1643 <= 1'b0; else if (1'b1) n1643 <= n3729;
/* FF 12 10  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1548 <= 1'b0; else if (n1430) n1548 <= n3730;
/* FF 10 10  7 */ always @(posedge io_13_31_1) if (n4) n1309 <= 1'b0 ? 1'b0 : n3731;
/* FF 10  2  3 */ assign n1245 = n3732;
/* FF 18 12  6 */ always @(posedge io_13_31_1) if (n2137) n2527 <= n3 ? 1'b0 : n3733;
/* FF  9  6  6 */ always @(posedge io_13_31_1) if (n4) n1119 <= 1'b0 ? 1'b0 : n3734;
/* FF 18  4  2 */ always @(posedge io_13_31_1) if (n2603) n2452 <= 1'b0 ? 1'b0 : n3735;
/* FF 22 16  5 */ assign n2980 = n3736;
/* FF 22  8  1 */ assign n2945 = n3737;
/* FF 21 12  4 */ always @(posedge io_13_31_1) if (n2663) n2815 <= 1'b0 ? 1'b0 : n3738;
/* FF 21  4  0 */ always @(posedge io_13_31_1) if (n2902) n2768 <= n7 ? 1'b0 : n3739;
/* FF  8 19  0 */ assign n3740 = n3741;
/* FF  3  3  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n357 <= 1'b0; else if (n198) n357 <= n3743;
/* FF 18 13  7 */ always @(posedge io_13_31_1) if (n2137) n2535 <= n3 ? 1'b0 : n3744;
/* FF 18  5  3 */ always @(posedge io_13_31_1) if (n2456) n2460 <= 1'b0 ? 1'b0 : n3745;
/* FF  5 20  3 */ assign n793 = n3746;
/* FF 17 21  4 */ assign n2423 = n3747;
/* FF 12  5  6 */ assign n1551 = n3748;
/* FF  8 20  1 */ assign n1060 = n3749;
/* FF 13  1  4 */ assign n3750 = n3751;
/* FF  2  8  5 */ assign n214 = n3752;
/* FF  4 19  7 */ assign n629 = n3753;
/* FF 14 14  3 */ assign n1957 = n3754;
/* FF 15 10  1 */ assign n2086 = n3755;
/* FF 12  6  7 */ assign n1279 = n3756;
/* FF 15 13  6 */ assign n2119 = n3757;
/* FF  5 16  5 */ assign n766 = n3758;
/* FF  4 12  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n581 <= 1'b0; else if (n432) n581 <= n3759;
/* FF 14 15  4 */ assign n1970 = n3760;
/* FF  2  4  7 */ assign n197 = n3761;
/* FF 23 13  1 */ assign n2842 = n3762;
/* FF 17 14  0 */ assign n3763 = n3764;
/* FF 11  2  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1396 <= 1'b0; else if (n1120) n1396 <= n3766;
/* FF  8 15  7 */ assign n3767 = n3768;
/* FF  8  7  3 */ assign n3769 = n3770;
/* FF 15  6  3 */ always @(posedge io_13_31_1) if (n2191) n1126 <= 1'b0 ? 1'b0 : n3771;
/* FF  5  8  6 */ assign n708 = n3772;
/* FF 13 23  0 */ assign n3773 = n3774;
/* FF 16 18  7 */ assign n3776 = n3777;
/* FF 16 10  3 */ assign n2224 = n3778;
/* FF 17  6  1 */ assign n1726 = n3779;
/* FF 14  2  6 */ assign n1408 = n3780;
/* FF  9 20  2 */ assign n1206 = n3781;
/* FF  5  1  3 */ assign n652 = n3782;
/* FF 17  9  6 */ always @(posedge io_13_31_1) if (n1591) n2346 <= 1'b0 ? 1'b0 : n3783;
/* FF 18 19  0 */ always @(posedge io_13_31_1) if (n2575) n2573 <= 1'b0 ? 1'b0 : n3784;
/* FF  7 12  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n889 <= 1'b0; else if (n818) n889 <= n3785;
/* FF  7  4  1 */ assign n843 = n3786;
/* FF  8  8  3 */ assign n988 = n3787;
/* FF 16 11  4 */ assign n2233 = n3788;
/* FF 16  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1555 <= 1'b0; else if (n1690) n1555 <= n3789;
/* FF 20 14  1 */ assign n3790 = n3791;
/* FF 17 10  7 */ always @(posedge io_13_31_1) if (n2213) n2370 <= 1'b0 ? 1'b0 : n3792;
/* FF 17  2  3 */ always @(posedge io_13_31_1) if (n2324) n2308 <= 1'b0 ? 1'b0 : n3793;
/* FF  3 21  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n485 <= 1'b0; else if (1'b1) n485 <= n3794;
/* FF  7  5  2 */ always @(posedge io_13_31_1) if (n4) n810 <= 1'b0 ? 1'b0 : n3795;
/* FF  9 16  4 */ assign n3796 = n3797;
/* FF 12 20  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1653 <= 1'b0; else if (n1654) n1653 <= n3798;
/* FF 14  3  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1554 <= 1'b0; else if (n1690) n1554 <= n3799;
/* FF 16  7  6 */ always @(posedge io_13_31_1) if (n2093) n2202 <= 1'b0 ? 1'b0 : n3800;
/* FF 13 19  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1715 <= 1'b0; else if (n1815) n1715 <= n3801;
/* FF  3 14  2 */ assign n3802 = n3803;
/* FF  1  6  5 */ assign n43 = n3804;
/* FF 10 12  6 */ assign n1326 = n3805;
/* FF 10  4  2 */ assign n1259 = n3806;
/* FF  9  8  5 */ assign n1132 = n3807;
/* FF  2 18  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n312 <= 1'b0; else if (n310) n312 <= n3808;
/* FF 13 12  4 */ assign n1761 = n3809;
/* FF 13  4  0 */ assign n1681 = n3810;
/* FF 21 14  3 */ always @(posedge io_13_31_1) if (n2842) n2832 <= 1'b0 ? 1'b0 : n3811;
/* FF 11 17  2 */ assign n1505 = n3812;
/* FF 12 13  0 */ assign n1610 = n3813;
/* FF 20  2  4 */ assign n2449 = n3814;
/* FF 18  7  2 */ always @(posedge io_13_31_1) if (n2076) n2478 <= 1'b0 ? 1'b0 : n3815;
/* FF 22 19  5 */ assign n2986 = n3816;
/* FF  2 19  4 */ assign n321 = n3817;
/* FF  2 11  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n251 <= 1'b0; else if (1'b1) n251 <= n3818;
/* FF 21 15  4 */ assign n2840 = n3819;
/* FF 11 18  3 */ assign n1510 = n3820;
/* FF 21  7  0 */ assign n3821 = n3822;
/* FF  8 22  0 */ assign n1072 = n3824;
/* FF 18  8  3 */ assign n2120 = n3825;
/* FF 12  9  2 */ assign n1585 = n3826;
/* FF  3  2  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n351 <= 1'b0; else if (n500) n351 <= n3827;
/* FF 12  8  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1576 <= 1'b0; else if (n1430) n1576 <= n3828;
/* FF 15 16  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1624 <= 1'b0; else if (n1811) n1624 <= n3829;
/* FF  2  3  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n181 <= 1'b0; else if (n17) n181 <= n3830;
/* FF  4 14  3 */ assign n593 = n3831;
/* FF 14 17  3 */ assign n1985 = n3832;
/* FF  8 18  2 */ assign n1053 = n3833;
/* FF 18  1  0 */ assign n3834 = n3835;
/* FF 17 17  1 */ always @(posedge io_13_31_1) if (1'b1) n2405 <= 1'b0 ? 1'b0 : n3837;
/* FF 11  5  5 */ assign n1420 = n3838;
/* FF 12  1  3 */ assign n3839 = n3840;
/* FF  5 19  5 */ assign n474 = n3841;
/* FF  5 11  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n731 <= 1'b0; else if (n128) n731 <= n3842;
/* FF  4 15  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n586 <= 1'b0; else if (n451) n586 <= n3843;
/* FF  4  7  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n542 <= 1'b0; else if (n532) n542 <= n3844;
/* FF  2  7  7 */ assign n223 = n3845;
/* FF 14 10  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1934 <= 1'b0; else if (n734) n1934 <= n3846;
/* FF  3  3  5 */ assign n360 = n3847;
/* FF 21  3  7 */ always @(posedge io_13_31_1) if (n2902) n2767 <= n7 ? 1'b0 : n3848;
/* FF 11  6  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1428 <= 1'b0; else if (n1426) n1428 <= n3849;
/* FF 15  9  3 */ always @(posedge io_13_31_1) if (n2213) n2080 <= 1'b0 ? 1'b0 : n3850;
/* FF  5 12  2 */ assign n739 = n3851;
/* FF  4  8  1 */ assign n548 = n3852;
/* FF 14  6  2 */ assign n1896 = n3853;
/* FF  8  3  0 */ assign n948 = n3854;
/* FF  1 21  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n153 <= 1'b0; else if (n80) n153 <= n3855;
/* FF 15  1  4 */ assign n1688 = n3856;
/* FF  7 15  5 */ assign n3857 = n3858;
/* FF  7  7  1 */ assign n854 = n3859;
/* FF  9 19  5 */ assign n1211 = n3860;
/* FF  4  3  7 */ assign n517 = n3861;
/* FF 16  6  0 */ assign n2184 = n3862;
/* FF  8  7  6 */ assign n981 = n3863;
/* FF 16  9  5 */ assign n2218 = n3864;
/* FF 17 13  7 */ always @(posedge io_13_31_1) if (n2536) n2257 <= n1 ? 1'b0 : n3865;
/* FF 17  5  3 */ always @(posedge io_13_31_1) if (n2456) n2337 <= 1'b0 ? 1'b0 : n3866;
/* FF 20 13  4 */ always @(posedge io_13_31_1) if (n2663) n2710 <= 1'b0 ? 1'b0 : n3867;
/* FF  7  8  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n866 <= 1'b0; else if (1'b1) n866 <= n3868;
/* FF 18 18  2 */ assign n2563 = n3869;
/* FF 16 10  6 */ assign n2227 = n3870;
/* FF 13 22  7 */ assign n1666 = n3871;
/* FF 13 14  3 */ assign n1785 = n3872;
/* FF  3 17  2 */ assign n133 = n3873;
/* FF 18 19  3 */ assign n3 = n3874;
/* FF  1  9  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n67 <= 1'b0; else if (n70) n67 <= n3875;
/* FF 20  5  5 */ always @(posedge io_13_31_1) if (n2472) n2675 <= n2471 ? 1'b0 : n3876;
/* FF  9 11  5 */ assign n1163 = n3877;
/* FF 13 15  4 */ assign n1797 = n3878;
/* FF 13  7  0 */ assign n1719 = n3879;
/* FF  1  2  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n10 <= 1'b0; else if (n17) n10 <= n3880;
/* FF 10  8  3 */ always @(posedge io_13_31_1) if (n4) n1285 <= 1'b0 ? 1'b0 : n3881;
/* FF 12 20  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1652 <= 1'b0; else if (n1654) n1652 <= n3882;
/* FF  9  4  2 */ assign n1102 = n3883;
/* FF 22 14  1 */ assign n2965 = n3884;
/* FF  2 14  0 */ assign n267 = n3885;
/* FF 13  8  1 */ assign n1733 = n3886;
/* FF  9  7  7 */ assign n1124 = n3887;
/* FF 13 11  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1454 <= 1'b0; else if (n734) n1454 <= n3888;
/* FF 10  1  0 */ assign n1234 = n3889;
/* FF 11 16  4 */ always @(posedge io_13_31_1) if (n4) n1499 <= 1'b0 ? 1'b0 : n3890;
/* FF 12 12  2 */ assign n1605 = n3891;
/* FF 22 15  2 */ assign n3892 = n3893;
/* FF  3  5  5 */ assign n378 = n3894;
/* FF 10  4  5 */ assign n974 = n3895;
/* FF 15 19  7 */ assign n2011 = n3896;
/* FF 22 18  7 */ assign n2991 = n3897;
/* FF  2  6  1 */ assign n3898 = n3899;
/* FF  5 14  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n266 <= 1'b0; else if (1'b1) n266 <= n3900;
/* FF 21 14  6 */ assign n2835 = n3901;
/* FF 11  9  1 */ always @(posedge io_13_31_1) if (n4) n1447 <= 1'b0 ? 1'b0 : n3902;
/* FF  8 21  2 */ assign n1067 = n3903;
/* FF 13  3  7 */ assign n1677 = n3904;
/* FF  3  6  6 */ assign n383 = n3905;
/* FF 17 20  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2292 <= 1'b0; else if (n2023) n2292 <= n3906;
/* FF 11  8  5 */ always @(posedge io_13_31_1) if (n4) n1440 <= 1'b0 ? 1'b0 : n3907;
/* FF 18  7  5 */ always @(posedge io_13_31_1) if (n2076) n2480 <= 1'b0 ? 1'b0 : n3908;
/* FF 15 12  4 */ assign n2107 = n3909;
/* FF 15  4  0 */ assign n1869 = n3910;
/* FF  4 18  4 */ assign n618 = n3911;
/* FF  4 10  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n565 <= 1'b0; else if (n576) n565 <= n3912;
/* FF  8 22  3 */ assign n1074 = n3913;
/* FF  2 10  7 */ assign n248 = n3914;
/* FF 14 13  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1789 <= 1'b0; else if (n735) n1789 <= n3915;
/* FF 22  2  4 */ always @(posedge io_13_31_1) if (1'b1) n2890 <= 1'b0 ? 1'b0 : n3916;
/* FF  2  2  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n170 <= 1'b0; else if (n178) n170 <= n3917;
/* FF 21  6  7 */ always @(posedge io_13_31_1) if (n2686) n2192 <= 1'b0 ? 1'b0 : n3918;
/* FF 11  1  2 */ assign n3919 = n3920;
/* FF  5 15  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n759 <= 1'b0; else if (n451) n759 <= n3921;
/* FF 17 24  7 */ assign n2438 = n3922;
/* FF 17 16  3 */ always @(posedge io_13_31_1) if (n2268) n2399 <= 1'b0 ? 1'b0 : n3923;
/* FF 11  4  7 */ assign n1415 = n3924;
/* FF  4 11  1 */ assign n270 = n3925;
/* FF 22  3  5 */ assign n2898 = n3926;
/* FF  2  3  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n184 <= 1'b0; else if (n17) n184 <= n3927;
/* FF  4 14  6 */ assign n595 = n3928;
/* FF  7 18  6 */ assign n3929 = n3930;
/* FF 14 17  6 */ always @(posedge io_13_31_1) if (1'b1) n1986 <= 1'b0 ? 1'b0 : n3931;
/* FF 14  9  2 */ always @(posedge io_13_31_1) if (n1739) n1928 <= 1'b0 ? 1'b0 : n3932;
/* FF 15  5  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1893 <= 1'b0; else if (n1869) n1893 <= n3933;
/* FF  8  6  0 */ assign n698 = n3934;
/* FF 20 20  2 */ always @(posedge io_13_31_1) if (n2738) n2742 <= 1'b0 ? 1'b0 : n3935;
/* FF  8  9  5 */ assign n985 = n3936;
/* FF 17  8  4 */ assign n2351 = n3937;
/* FF 10 18  2 */ assign n3938 = n3939;
/* FF  9 22  5 */ assign n1227 = n3940;
/* FF  5  2  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n389 <= 1'b0; else if (n509) n389 <= n3941;
/* FF  9 14  1 */ assign n1183 = n3942;
/* FF  4  6  7 */ assign n535 = n3943;
/* FF  8 10  6 */ assign n1010 = n3944;
/* FF  8  2  2 */ assign n942 = n3945;
/* FF  1 20  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n146 <= 1'b0; else if (n147) n146 <= n3946;
/* FF 16 12  5 */ assign n2243 = n3947;
/* FF 10 19  3 */ assign n1374 = n3948;
/* FF  5  3  5 */ assign n668 = n3949;
/* FF  9 15  2 */ assign n1191 = n3950;
/* FF 18 21  2 */ assign n2584 = n3951;
/* FF 17  4  6 */ always @(posedge io_13_31_1) if (n2316) n2331 <= 1'b0 ? 1'b0 : n3952;
/* FF 23  3  7 */ always @(posedge io_13_31_1) if (1'b1) n3011 <= n2888 ? 1'b0 : n3953;
/* FF 16 13  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2067 <= 1'b0; else if (n735) n2067 <= n3954;
/* FF 16  5  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2179 <= 1'b0; else if (n1869) n2179 <= n3955;
/* FF  3 20  2 */ assign n478 = n3956;
/* FF 20  9  1 */ always @(posedge io_13_31_1) if (n2093) n2229 <= 1'b0 ? 1'b0 : n3957;
/* FF 18 22  3 */ always @(posedge io_13_31_1) if (n2582) n2589 <= 1'b0 ? 1'b0 : n3958;
/* FF  1 12  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n87 <= 1'b0; else if (1'b1) n87 <= n3959;
/* FF  7  7  4 */ assign n857 = n3960;
/* FF 12 22  6 */ assign n1664 = n3961;
/* FF 22 17  2 */ always @(posedge io_13_31_1) if (n2737) n2984 <= 1'b0 ? 1'b0 : n3962;
/* FF  2 17  1 */ assign n3963 = n3964;
/* FF 13 10  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1753 <= 1'b0; else if (n734) n1753 <= n3965;
/* FF 10  6  5 */ assign n984 = n3966;
/* FF  9  2  4 */ assign n1087 = n3967;
/* FF  3 16  4 */ assign n448 = n3968;
/* FF 20  1  2 */ always @(posedge io_13_31_1) if (n2600) n2447 <= n2758 ? 1'b0 : n3969;
/* FF 12 15  3 */ assign n1181 = n3970;
/* FF 20  4  7 */ assign n2672 = n3971;
/* FF 10  7  6 */ always @(posedge io_13_31_1) if (n4) n1277 <= 1'b0 ? 1'b0 : n3972;
/* FF 21 13  0 */ assign n3973 = n3974;
/* FF 24 21  1 */ always @(posedge io_13_31_1) if (n2995) n3042 <= 1'b0 ? 1'b0 : n3976;
/* FF  4 21  0 */ assign n3977 = n3978;
/* FF 13 14  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1632 <= 1'b0; else if (n604) n1632 <= n3980;
/* FF  2 21  7 */ assign n150 = n3981;
/* FF 22 13  4 */ assign n2663 = n3982;
/* FF  3 17  5 */ assign n112 = n3983;
/* FF  3  9  1 */ assign n414 = n3984;
/* FF 11 19  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1508 <= 1'b0; else if (1'b1) n1508 <= n3985;
/* FF 18 10  6 */ assign n2507 = n3986;
/* FF  9  3  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n966 <= 1'b0; else if (n851) n966 <= n3987;
/* FF 18  2  2 */ assign n2333 = n3988;
/* FF 21 17  6 */ assign n2852 = n3989;
/* FF 21  9  2 */ always @(posedge io_13_31_1) if (1'b1) n175 <= 1'b0 ? 1'b0 : n3990;
/* FF 11 12  1 */ assign n1472 = n3991;
/* FF 13  6  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1702 <= 1'b0; else if (n1433) n1702 <= n3992;
/* FF  2  5  4 */ assign n205 = n3993;
/* FF  3  1  2 */ assign n340 = n3994;
/* FF 14 19  6 */ assign n1998 = n3995;
/* FF 15 15  4 */ assign n2121 = n3996;
/* FF  3  4  7 */ assign n370 = n3997;
/* FF 15  7  0 */ assign n1915 = n3998;
/* FF  7 21  1 */ assign n924 = n3999;
/* FF 12  3  6 */ assign n4000 = n4001;
/* FF 22  5  4 */ assign n2929 = n4002;
/* FF  5 13  4 */ assign n745 = n4003;
/* FF  4 17  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n315 <= 1'b0; else if (n317) n315 <= n4004;
/* FF  4  9  3 */ assign n559 = n4005;
/* FF 15  8  1 */ always @(posedge io_13_31_1) if (n1591) n2069 <= 1'b0 ? 1'b0 : n4006;
/* FF 17 19  3 */ assign n4007 = n4008;
/* FF 11  7  7 */ assign n1187 = n4009;
/* FF 15 11  6 */ assign n2100 = n4010;
/* FF  2  6  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n51 <= 1'b0; else if (n217) n51 <= n4011;
/* FF  5 14  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n296 <= 1'b0; else if (1'b1) n296 <= n4012;
/* FF 14 12  2 */ assign n1943 = n4013;
/* FF 17 12  0 */ always @(posedge io_13_31_1) if (n2137) n2380 <= n3 ? 1'b0 : n4014;
/* FF 15  4  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1903 <= 1'b0; else if (n1547) n1903 <= n4015;
/* FF 23 14  6 */ always @(posedge io_13_31_1) if (1'b1) n3024 <= 1'b0 ? 1'b0 : n4016;
/* FF  5  6  0 */ assign n4017 = n4018;
/* FF 15  3  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1689 <= 1'b0; else if (n1547) n1689 <= n4020;
/* FF 22  2  7 */ assign n2893 = n4021;
/* FF 16 16  1 */ assign n2271 = n4022;
/* FF  9 17  1 */ assign n1199 = n4023;
/* FF 13 21  0 */ assign n1830 = n4024;
/* FF  7  9  4 */ assign n864 = n4025;
/* FF  8 13  6 */ assign n1029 = n4026;
/* FF  8  5  2 */ assign n958 = n4027;
/* FF 20 11  0 */ always @(posedge io_13_31_1) if (n2137) n2695 <= n3 ? 1'b0 : n4028;
/* FF  9 18  2 */ assign n4029 = n4030;
/* FF 17  7  6 */ assign n1739 = n4031;
/* FF  7 10  5 */ assign n576 = n4032;
/* FF  7  2  1 */ assign n830 = n4033;
/* FF  9 21  7 */ assign n1226 = n4034;
/* FF  8  6  3 */ assign n978 = n4035;
/* FF  1 16  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n119 <= 1'b0; else if (n127) n119 <= n4036;
/* FF 16  8  2 */ always @(posedge io_13_31_1) if (n2344) n2207 <= 1'b0 ? 1'b0 : n4037;
/* FF 20 20  5 */ assign n2744 = n4038;
/* FF 20 12  1 */ assign n2704 = n4039;
/* FF 10 15  0 */ always @(posedge io_13_31_1) if (n4) n1352 <= 1'b0 ? 1'b0 : n4040;
/* FF 17  8  7 */ always @(posedge io_13_31_1) if (n2344) n2354 <= 1'b0 ? 1'b0 : n4041;
/* FF 10 18  5 */ assign n4042 = n4043;
/* FF  3 19  5 */ assign n471 = n4044;
/* FF  5  2  7 */ assign n662 = n4045;
/* FF  9 14  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1046 <= 1'b0; else if (n762) n1046 <= n4046;
/* FF  2 20  1 */ assign n160 = n4047;
/* FF  1  8  2 */ assign n4048 = n4049;
/* FF 13 17  7 */ assign n4050 = n4051;
/* FF  3 11  0 */ assign n17 = n4052;
/* FF  1 11  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n78 <= 1'b1; else if (n245) n78 <= n4053;
/* FF 12 18  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1642 <= 1'b0; else if (1'b1) n1642 <= n4054;
/* FF 20  7  7 */ assign n4055 = n4056;
/* FF 10 10  6 */ assign n1308 = n4057;
/* FF 10  2  2 */ assign n1243 = n4058;
/* FF  9  6  5 */ assign n1116 = n4059;
/* FF 22 16  4 */ assign n2971 = n4060;
/* FF  2 16  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n294 <= 1'b0; else if (n127) n294 <= n4061;
/* FF  3 20  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n334 <= 1'b0; else if (n629) n334 <= n4062;
/* FF 13  9  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1718 <= 1'b0; else if (n734) n1718 <= n4063;
/* FF  3 12  1 */ assign n431 = n4064;
/* FF 22  8  0 */ assign n2066 = n4065;
/* FF 21 20  7 */ assign n2867 = n4066;
/* FF 21 12  3 */ assign n2814 = n4067;
/* FF  1  4  4 */ assign n31 = n4068;
/* FF 18 13  6 */ always @(posedge io_13_31_1) if (n2137) n2534 <= n3 ? 1'b0 : n4069;
/* FF 12 14  5 */ assign n1621 = n4070;
/* FF 18  5  2 */ always @(posedge io_13_31_1) if (n2456) n2459 <= 1'b0 ? 1'b0 : n4071;
/* FF  2 17  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n132 <= 1'b0; else if (1'b1) n132 <= n4072;
/* FF 13 10  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1706 <= 1'b0; else if (n734) n1706 <= n4073;
/* FF  2  9  0 */ assign n4074 = n4075;
/* FF  9  2  7 */ assign n1090 = n4077;
/* FF 11 15  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1488 <= 1'b0; else if (1'b1) n1488 <= n4078;
/* FF 14 23  2 */ assign n2032 = n4079;
/* FF  8 20  0 */ assign n4080 = n4081;
/* FF 10  3  2 */ assign n1251 = n4082;
/* FF 18  6  3 */ always @(posedge io_13_31_1) if (n2602) n2467 <= n1 ? 1'b0 : n4083;
/* FF  3  7  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n401 <= 1'b0; else if (n224) n401 <= n4084;
/* FF 21 13  3 */ always @(posedge io_13_31_1) if (n2819) n2821 <= n2823 ? 1'b0 : n4085;
/* FF 12  6  6 */ assign n1562 = n4086;
/* FF  5 16  4 */ assign n765 = n4087;
/* FF  4 20  7 */ assign n640 = n4088;
/* FF 23 22  0 */ always @(posedge io_13_31_1) if (n3003) n2755 <= 1'b0 ? 1'b0 : n4089;
/* FF  4 12  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n580 <= 1'b0; else if (n432) n580 <= n4090;
/* FF 14 15  3 */ assign n1478 = n4091;
/* FF  8 16  2 */ assign n922 = n4092;
/* FF  2  4  6 */ always @(posedge io_13_31_1) if (n201) n191 <= n42 ? 1'b0 : n4093;
/* FF 22  4  7 */ assign n2915 = n4094;
/* FF 15 14  6 */ assign n2123 = n4095;
/* FF  5 17  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n772 <= 1'b0; else if (1'b1) n772 <= n4096;
/* FF 15  6  2 */ assign n2056 = n4097;
/* FF  2  1  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n161 <= 1'b0; else if (n178) n161 <= n4098;
/* FF  5  9  1 */ always @(posedge io_13_31_1) if (n4) n715 <= 1'b0 ? 1'b0 : n4099;
/* FF  4 13  4 */ assign n4100 = n4101;
/* FF  4  5  0 */ assign n526 = n4102;
/* FF  2  5  7 */ assign n207 = n4103;
/* FF 16 19  2 */ assign n2286 = n4104;
/* FF 11  3  4 */ assign n1402 = n4105;
/* FF 14 11  5 */ assign n1940 = n4106;
/* FF 15  7  3 */ assign n2061 = n4107;
/* FF 20 22  5 */ assign n2753 = n4108;
/* FF 22  5  7 */ assign n2472 = n4109;
/* FF  5  1  2 */ assign n651 = n4110;
/* FF  8  8  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n812 <= 1'b0; else if (n877) n812 <= n4111;
/* FF  5  4  7 */ assign n677 = n4112;
/* FF 16 11  3 */ assign n2232 = n4113;
/* FF 20 14  0 */ assign n4114 = n4115;
/* FF 17 10  6 */ assign n2364 = n4117;
/* FF  7 13  5 */ always @(posedge io_13_31_1) if (n4) n899 <= 1'b0 ? 1'b0 : n4118;
/* FF 17  2  2 */ always @(posedge io_13_31_1) if (n2324) n2307 <= 1'b0 ? 1'b0 : n4119;
/* FF  7  5  1 */ assign n848 = n4120;
/* FF  9 16  3 */ assign n4121 = n4122;
/* FF  1 19  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n135 <= 1'b0; else if (n140) n135 <= n4123;
/* FF  4  1  7 */ assign n499 = n4124;
/* FF 20 15  1 */ always @(posedge io_13_31_1) if (n2722) n2721 <= 1'b0 ? 1'b0 : n4125;
/* FF 14  3  5 */ assign n1873 = n4126;
/* FF  8  4  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n964 <= 1'b0; else if (n663) n964 <= n4127;
/* FF 16  7  5 */ assign n2201 = n4128;
/* FF 20 18  6 */ assign n2733 = n4129;
/* FF 17  3  3 */ always @(posedge io_13_31_1) if (n2324) n2319 <= 1'b0 ? 1'b0 : n4130;
/* FF  7  6  2 */ always @(posedge io_13_31_1) if (n4) n710 <= 1'b0 ? 1'b0 : n4131;
/* FF 10 13  1 */ assign n1334 = n4132;
/* FF  9 17  4 */ always @(posedge io_13_31_1) if (1'b1) n1202 <= 1'b0 ? 1'b0 : n4133;
/* FF  9  9  0 */ assign n1136 = n4134;
/* FF  7  9  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n90 <= 1'b0; else if (1'b1) n90 <= n4135;
/* FF 13 20  7 */ always @(posedge io_13_31_1) if (n1838) n1829 <= 1'b0 ? 1'b0 : n4136;
/* FF 13 12  3 */ assign n1760 = n4137;
/* FF 20 11  3 */ always @(posedge io_13_31_1) if (n2137) n2698 <= n3 ? 1'b0 : n4138;
/* FF 18 16  1 */ always @(posedge io_13_31_1) if (n2011) n2552 <= 1'b0 ? 1'b0 : n4139;
/* FF 20 10  7 */ always @(posedge io_13_31_1) if (n2112) n2631 <= 1'b0 ? 1'b0 : n4140;
/* FF  3 18  7 */ assign n464 = n4141;
/* FF 22 20  0 */ assign n8 = n4142;
/* FF  9  1  1 */ assign n1077 = n4143;
/* FF  2 19  3 */ assign n306 = n4144;
/* FF 13 13  4 */ always @(posedge io_13_31_1) if (1'b1) n1774 <= 1'b0 ? 1'b0 : n4145;
/* FF 22 19  4 */ assign n2993 = n4146;
/* FF  3 15  1 */ assign n439 = n4147;
/* FF 21 15  3 */ always @(posedge io_13_31_1) if (n2828) n2839 <= 1'b0 ? 1'b0 : n4148;
/* FF 11 18  2 */ always @(posedge io_13_31_1) if (1'b1) n1509 <= 1'b0 ? 1'b0 : n4149;
/* FF  1  7  4 */ assign n48 = n4150;
/* FF 12 17  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1637 <= 1'b0; else if (1'b1) n1637 <= n4151;
/* FF 18  8  2 */ assign n1591 = n4152;
/* FF  2 20  4 */ assign n158 = n4153;
/* FF 12  9  1 */ assign n1584 = n4154;
/* FF 22 12  1 */ assign n2826 = n4155;
/* FF  2 12  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n70 <= 1'b0; else if (1'b1) n70 <= n4156;
/* FF 18 11  7 */ always @(posedge io_13_31_1) if (n2137) n2519 <= n3 ? 1'b0 : n4157;
/* FF 21  8  0 */ assign n2799 = n4158;
/* FF  9  5  7 */ assign n1114 = n4159;
/* FF  3 11  3 */ assign n102 = n4160;
/* FF 11 14  4 */ always @(posedge io_13_31_1) if (n1180) n1482 <= n1 ? 1'b0 : n4161;
/* FF 12 10  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1577 <= 1'b0; else if (n1430) n1577 <= n4162;
/* FF 10  2  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1247 <= 1'b0; else if (n979) n1247 <= n4163;
/* FF 22 16  7 */ assign n2982 = n4164;
/* FF  5 19  4 */ assign n785 = n4165;
/* FF 22  8  3 */ always @(posedge io_13_31_1) if (1'b1) n2946 <= n2802 ? 1'b0 : n4166;
/* FF 21 12  6 */ assign n2817 = n4167;
/* FF 21  4  2 */ always @(posedge io_13_31_1) if (n2902) n2770 <= n7 ? 1'b0 : n4168;
/* FF  4 15  3 */ assign n603 = n4169;
/* FF  8 19  2 */ assign n4170 = n4171;
/* FF  2  7  6 */ assign n222 = n4172;
/* FF  3  3  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n359 <= 1'b0; else if (n198) n359 <= n4173;
/* FF 11  6  5 */ assign n1425 = n4174;
/* FF 18  5  5 */ always @(posedge io_13_31_1) if (n2456) n2462 <= 1'b0 ? 1'b0 : n4175;
/* FF  5 20  5 */ assign n795 = n4176;
/* FF 15  9  2 */ assign n2079 = n4177;
/* FF 23 20  7 */ always @(posedge io_13_31_1) if (n2997) n3034 <= 1'b0 ? 1'b0 : n4178;
/* FF  5 12  1 */ assign n735 = n4179;
/* FF 17 21  6 */ assign n2431 = n4180;
/* FF  4  8  0 */ assign n4181 = n4182;
/* FF  8 20  3 */ assign n1062 = n4184;
/* FF  2  8  7 */ assign n231 = n4185;
/* FF 13  1  6 */ assign n4186 = n4187;
/* FF 16 22  2 */ assign n2294 = n4188;
/* FF 17 18  0 */ assign n4189 = n4190;
/* FF 14 14  5 */ assign n1962 = n4192;
/* FF 14  6  1 */ assign n1895 = n4193;
/* FF 15 10  3 */ always @(posedge io_13_31_1) if (n1591) n2087 <= 1'b0 ? 1'b0 : n4194;
/* FF 23 12  2 */ always @(posedge io_13_31_1) if (n2826) n2509 <= n2957 ? 1'b0 : n4195;
/* FF  7 16  0 */ assign n4196 = n4197;
/* FF  5 16  7 */ assign n767 = n4198;
/* FF  4 12  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n271 <= 1'b0; else if (n432) n271 <= n4199;
/* FF 14 15  6 */ assign n1781 = n4200;
/* FF 17 14  2 */ always @(posedge io_13_31_1) if (n2396) n2391 <= n1 ? 1'b0 : n4201;
/* FF  8  7  5 */ assign n4202 = n4203;
/* FF 17 13  6 */ always @(posedge io_13_31_1) if (n2536) n2388 <= n1 ? 1'b0 : n4204;
/* FF 20 21  7 */ assign n2750 = n4205;
/* FF 20 13  3 */ always @(posedge io_13_31_1) if (n2663) n2709 <= 1'b0 ? 1'b0 : n4206;
/* FF  7  8  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n865 <= 1'b0; else if (1'b1) n865 <= n4207;
/* FF 14  7  1 */ assign n1906 = n4208;
/* FF  4  4  7 */ assign n523 = n4209;
/* FF  7 11  6 */ assign n631 = n4210;
/* FF 13 23  2 */ assign n1856 = n4211;
/* FF 16 10  5 */ always @(posedge io_13_31_1) if (n2112) n2226 <= 1'b0 ? 1'b0 : n4212;
/* FF 17  6  3 */ assign n2065 = n4213;
/* FF 16  2  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1884 <= 1'b0; else if (n1552) n1884 <= n4214;
/* FF  9 20  4 */ assign n1216 = n4215;
/* FF  5  1  5 */ assign n654 = n4216;
/* FF  9 12  0 */ assign n4217 = n4218;
/* FF 18 19  2 */ assign n2568 = n4220;
/* FF  7 12  7 */ assign n890 = n4221;
/* FF  8  8  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n878 <= 1'b0; else if (n877) n878 <= n4222;
/* FF  7  4  3 */ assign n844 = n4223;
/* FF 16 11  6 */ assign n2235 = n4224;
/* FF 16  3  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1678 <= 1'b0; else if (n1690) n1678 <= n4225;
/* FF 20 14  3 */ assign n2715 = n4226;
/* FF 17  2  5 */ assign n2310 = n4227;
/* FF  3 21  7 */ assign n487 = n4228;
/* FF  1  2  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n9 <= 1'b0; else if (n17) n9 <= n4229;
/* FF  9 16  6 */ assign n4230 = n4231;
/* FF 13  8  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n212 <= 1'b0; else if (n1860) n212 <= n4232;
/* FF 13 11  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1705 <= 1'b0; else if (n734) n1705 <= n4233;
/* FF  3 14  4 */ assign n92 = n4234;
/* FF  1  6  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n16 <= 1'b0; else if (n17) n16 <= n4235;
/* FF 12 12  1 */ assign n1604 = n4236;
/* FF 22 15  1 */ assign n2972 = n4237;
/* FF  2 15  0 */ assign n286 = n4238;
/* FF 10  4  4 */ assign n1258 = n4239;
/* FF  9  8  7 */ always @(posedge io_13_31_1) if (n4) n1134 <= 1'b0 ? 1'b0 : n4240;
/* FF 21 11  0 */ always @(posedge io_13_31_1) if (n2213) n2365 <= 1'b0 ? 1'b0 : n4241;
/* FF 22 18  6 */ always @(posedge io_13_31_1) if (n2989) n2990 <= 1'b0 ? 1'b0 : n4242;
/* FF  1  3  1 */ assign n19 = n4243;
/* FF  2 18  5 */ assign n307 = n4244;
/* FF 13 12  6 */ assign n1475 = n4245;
/* FF 13  4  2 */ assign n1682 = n4246;
/* FF 21 14  5 */ assign n2834 = n4247;
/* FF 11  9  0 */ always @(posedge io_13_31_1) if (n4) n1446 <= 1'b0 ? 1'b0 : n4248;
/* FF 12 13  2 */ assign n1612 = n4249;
/* FF 20  2  6 */ always @(posedge io_13_31_1) if (n2324) n2669 <= 1'b0 ? 1'b0 : n4250;
/* FF 10  5  5 */ assign n1265 = n4251;
/* FF  3  6  5 */ assign n387 = n4252;
/* FF 24 19  0 */ always @(posedge io_13_31_1) if (n2868) n3055 <= 1'b0 ? 1'b0 : n4253;
/* FF  9  1  4 */ assign n1079 = n4254;
/* FF 15 20  7 */ assign n1815 = n4255;
/* FF 22 19  7 */ assign n2992 = n4256;
/* FF 22 11  3 */ always @(posedge io_13_31_1) if (n2955) n1608 <= 1'b0 ? 1'b0 : n4257;
/* FF  2 11  2 */ assign n253 = n4258;
/* FF 21  7  2 */ assign n2791 = n4259;
/* FF 11 10  1 */ assign n1456 = n4260;
/* FF  8 22  2 */ always @(posedge io_13_31_1) if (1'b1) n1073 <= 1'b0 ? 1'b0 : n4261;
/* FF 18  8  5 */ always @(posedge io_13_31_1) if (n2120) n2489 <= 1'b0 ? 1'b0 : n4262;
/* FF  3  2  7 */ assign n353 = n4263;
/* FF  5 15  1 */ assign n758 = n4264;
/* FF 17 16  2 */ always @(posedge io_13_31_1) if (n2268) n2398 <= 1'b0 ? 1'b0 : n4265;
/* FF  4 11  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n577 <= 1'b0; else if (1'b1) n577 <= n4266;
/* FF 22  3  4 */ always @(posedge io_13_31_1) if (1'b1) n2897 <= n2757 ? 1'b0 : n4267;
/* FF  2  3  3 */ assign n183 = n4268;
/* FF  4 14  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n594 <= 1'b0; else if (1'b1) n594 <= n4269;
/* FF 14 17  5 */ assign n1967 = n4270;
/* FF  8 18  4 */ assign n1055 = n4271;
/* FF 14  9  1 */ always @(posedge io_13_31_1) if (n1739) n1927 <= 1'b0 ? 1'b0 : n4272;
/* FF 17 17  3 */ always @(posedge io_13_31_1) if (1'b1) n2404 <= 1'b0 ? 1'b0 : n4273;
/* FF 11  5  7 */ assign n1421 = n4274;
/* FF  7 19  0 */ assign n4275 = n4276;
/* FF 12  1  5 */ assign n4277 = n4278;
/* FF  5 19  7 */ assign n787 = n4279;
/* FF  5 11  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n732 <= 1'b0; else if (n128) n732 <= n4280;
/* FF  4 15  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n450 <= 1'b0; else if (n451) n450 <= n4281;
/* FF  4  7  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n545 <= 1'b0; else if (n532) n545 <= n4282;
/* FF 14 10  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1925 <= 1'b0; else if (n734) n1925 <= n4283;
/* FF  8 11  1 */ always @(posedge io_13_31_1) if (n4) n1013 <= 1'b0 ? 1'b0 : n4284;
/* FF 15  9  5 */ assign n2082 = n4285;
/* FF  1 20  3 */ assign n145 = n4286;
/* FF  5  4  0 */ assign n672 = n4287;
/* FF 10 19  2 */ assign n930 = n4288;
/* FF  5  3  4 */ assign n667 = n4289;
/* FF 16 14  1 */ assign n2253 = n4290;
/* FF 14  6  4 */ assign n1898 = n4291;
/* FF  8  3  2 */ assign n950 = n4292;
/* FF 16 13  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2204 <= 1'b0; else if (n735) n2204 <= n4293;
/* FF  1 13  0 */ assign n4294 = n4295;
/* FF 20 17  4 */ always @(posedge io_13_31_1) if (n2566) n2725 <= 1'b0 ? 1'b0 : n4297;
/* FF 20  9  0 */ assign n2093 = n4298;
/* FF 18 22  2 */ assign n2588 = n4299;
/* FF  7 15  7 */ assign n4300 = n4301;
/* FF  7  7  3 */ always @(posedge io_13_31_1) if (n4) n856 <= 1'b0 ? 1'b0 : n4302;
/* FF  9 19  7 */ assign n1213 = n4303;
/* FF 16  6  2 */ assign n2186 = n4304;
/* FF 16  9  7 */ assign n2220 = n4305;
/* FF 20 13  6 */ always @(posedge io_13_31_1) if (n2663) n2712 <= 1'b0 ? 1'b0 : n4306;
/* FF  7  8  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n868 <= 1'b0; else if (1'b1) n868 <= n4307;
/* FF 20 10  0 */ assign n2213 = n4308;
/* FF  2 21  6 */ assign n333 = n4309;
/* FF 13 14  5 */ assign n1787 = n4310;
/* FF  3 17  4 */ assign n363 = n4311;
/* FF  3  9  0 */ assign n4312 = n4313;
/* FF 18 19  5 */ assign n2574 = n4315;
/* FF 20  5  7 */ assign n2471 = n4316;
/* FF  9 11  7 */ always @(posedge io_13_31_1) if (n4) n1165 <= 1'b0 ? 1'b0 : n4317;
/* FF  4 22  0 */ assign n641 = n4318;
/* FF  9  3  3 */ assign n1093 = n4319;
/* FF 13 15  6 */ always @(posedge io_13_31_1) if (1'b1) n1799 <= 1'b0 ? 1'b0 : n4320;
/* FF 13  7  2 */ assign n1720 = n4321;
/* FF 21 17  5 */ assign n2851 = n4322;
/* FF  3 10  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n60 <= 1'b0; else if (n576) n60 <= n4323;
/* FF 11 20  4 */ assign n1515 = n4324;
/* FF 11 12  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1329 <= 1'b0; else if (n102) n1329 <= n4325;
/* FF  1  2  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n12 <= 1'b0; else if (n17) n12 <= n4326;
/* FF 18 11  0 */ always @(posedge io_13_31_1) if (n2137) n2512 <= n3 ? 1'b0 : n4327;
/* FF 10  8  5 */ assign n1287 = n4328;
/* FF  9  4  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1104 <= 1'b0; else if (n840) n1104 <= n4329;
/* FF 22 22  7 */ assign n2593 = n4330;
/* FF 22 14  3 */ assign n2967 = n4331;
/* FF  2 14  2 */ assign n281 = n4332;
/* FF 21 18  6 */ assign n2666 = n4333;
/* FF 21 10  2 */ always @(posedge io_13_31_1) if (n2137) n2807 <= n3 ? 1'b1 : n4334;
/* FF 11 16  6 */ assign n1501 = n4335;
/* FF 12 12  4 */ assign n1606 = n4336;
/* FF 18  3  1 */ always @(posedge io_13_31_1) if (n2191) n1868 <= 1'b0 ? 1'b0 : n4337;
/* FF 12  4  0 */ assign n1422 = n4338;
/* FF  3  5  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n213 <= 1'b0; else if (n532) n213 <= n4339;
/* FF 15  8  0 */ assign n2068 = n4340;
/* FF 22  7  0 */ always @(posedge io_13_31_1) if (n2694) n2794 <= n1 ? 1'b0 : n4341;
/* FF 15 11  5 */ always @(posedge io_13_31_1) if (n2112) n2099 <= 1'b0 ? 1'b0 : n4342;
/* FF  2  6  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n200 <= 1'b0; else if (n217) n200 <= n4343;
/* FF  5 14  4 */ assign n755 = n4344;
/* FF  8 21  4 */ assign n1069 = n4345;
/* FF 17 20  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2426 <= 1'b0; else if (n2023) n2426 <= n4346;
/* FF 11  8  7 */ always @(posedge io_13_31_1) if (n4) n1442 <= 1'b0 ? 1'b0 : n4347;
/* FF 15 12  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1754 <= 1'b0; else if (n735) n1754 <= n4348;
/* FF 15  4  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1699 <= 1'b0; else if (n1547) n1699 <= n4349;
/* FF  4 18  6 */ assign n619 = n4350;
/* FF  4 10  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n568 <= 1'b0; else if (n576) n568 <= n4351;
/* FF 14 13  2 */ assign n1950 = n4352;
/* FF  8 14  1 */ assign n1036 = n4353;
/* FF  2  2  5 */ assign n172 = n4354;
/* FF 22  2  6 */ always @(posedge io_13_31_1) if (1'b1) n2892 <= 1'b0 ? 1'b0 : n4355;
/* FF 16 16  0 */ always @(posedge io_13_31_1) if (1'b1) n2270 <= 1'b0 ? 1'b0 : n4356;
/* FF 14 16  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1980 <= 1'b0; else if (n1967) n1980 <= n4357;
/* FF 11  1  4 */ assign n4358 = n4359;
/* FF  5 15  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n610 <= 1'b0; else if (n451) n610 <= n4360;
/* FF 23 15  6 */ always @(posedge io_13_31_1) if (n2982) n3033 <= 1'b0 ? 1'b0 : n4361;
/* FF  5  7  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n695 <= 1'b0; else if (n532) n695 <= n4362;
/* FF 23  7  2 */ assign n2676 = n4363;
/* FF 24  3  0 */ always @(posedge io_13_31_1) if (n2902) n2894 <= n7 ? 1'b0 : n4364;
/* FF 22  3  7 */ assign n2900 = n4365;
/* FF  9 18  1 */ assign n4366 = n4367;
/* FF 16 17  1 */ always @(posedge io_13_31_1) if (n2273) n1645 <= n1 ? 1'b0 : n4368;
/* FF 14  9  4 */ always @(posedge io_13_31_1) if (n1739) n1597 <= 1'b0 ? 1'b0 : n4369;
/* FF  8  6  2 */ assign n976 = n4370;
/* FF  1 16  0 */ assign n4371 = n4372;
/* FF 20 20  4 */ assign n2738 = n4374;
/* FF  8  9  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n880 <= 1'b0; else if (n877) n880 <= n4375;
/* FF 20 12  0 */ assign n2703 = n4376;
/* FF 17  8  6 */ always @(posedge io_13_31_1) if (n2344) n2353 <= 1'b0 ? 1'b0 : n4377;
/* FF 10 18  4 */ assign n4378 = n4379;
/* FF  9 22  7 */ assign n1233 = n4380;
/* FF  5  2  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n658 <= 1'b0; else if (n509) n658 <= n4381;
/* FF  9 14  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1184 <= 1'b0; else if (n762) n1184 <= n4382;
/* FF  1 17  1 */ assign n4383 = n4384;
/* FF  8  2  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n944 <= 1'b0; else if (n840) n944 <= n4385;
/* FF  1 20  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n148 <= 1'b0; else if (n147) n148 <= n4386;
/* FF 16 12  7 */ always @(posedge io_13_31_1) if (n2120) n2244 <= 1'b0 ? 1'b0 : n4387;
/* FF 16  4  3 */ always @(posedge io_13_31_1) if (n2324) n2175 <= 1'b0 ? 1'b0 : n4388;
/* FF 10 19  5 */ assign n1376 = n4389;
/* FF  7  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n834 <= 1'b0; else if (n663) n834 <= n4390;
/* FF 10 11  1 */ always @(posedge io_13_31_1) if (n4) n1311 <= 1'b0 ? 1'b0 : n4391;
/* FF  5  3  7 */ assign n670 = n4392;
/* FF  9 15  4 */ assign n1193 = n4393;
/* FF 16  5  4 */ assign n1563 = n4394;
/* FF 17  1  2 */ assign n2304 = n4395;
/* FF  3 20  4 */ assign n466 = n4396;
/* FF  3 12  0 */ assign n430 = n4397;
/* FF  1 12  7 */ assign n89 = n4398;
/* FF 18 14  1 */ always @(posedge io_13_31_1) if (n2137) n2542 <= n3 ? 1'b0 : n4399;
/* FF  1  4  3 */ always @(posedge io_13_31_1) if (n201) n30 <= n42 ? 1'b0 : n4400;
/* FF 21 21  1 */ assign n2871 = n4401;
/* FF 12 14  4 */ assign n1620 = n4402;
/* FF 22 17  4 */ assign n2985 = n4403;
/* FF  2 17  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n300 <= 1'b0; else if (1'b1) n300 <= n4404;
/* FF 13 10  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1752 <= 1'b0; else if (n734) n1752 <= n4405;
/* FF  3 13  1 */ assign n4406 = n4407;
/* FF  9  2  6 */ assign n1089 = n4408;
/* FF  1  5  4 */ always @(posedge io_13_31_1) if (n201) n26 <= n42 ? 1'b0 : n4409;
/* FF 11 15  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1487 <= 1'b0; else if (1'b1) n1487 <= n4410;
/* FF 14 23  1 */ assign n2031 = n4411;
/* FF  3 16  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n304 <= 1'b0; else if (1'b1) n304 <= n4412;
/* FF 20  1  4 */ always @(posedge io_13_31_1) if (n2600) n2595 <= n2758 ? 1'b0 : n4413;
/* FF 10  3  1 */ assign n1252 = n4414;
/* FF 12 15  5 */ assign n4 = n4415;
/* FF 18  6  2 */ always @(posedge io_13_31_1) if (n2602) n2466 <= n1 ? 1'b0 : n4416;
/* FF 12  7  1 */ assign n1568 = n4417;
/* FF 21 13  2 */ always @(posedge io_13_31_1) if (n2819) n2820 <= n2823 ? 1'b0 : n4418;
/* FF  4 21  2 */ assign n645 = n4419;
/* FF 18  9  7 */ assign n2498 = n4420;
/* FF 15 20  0 */ assign n2152 = n4421;
/* FF  3  9  3 */ assign n416 = n4422;
/* FF  3  8  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n409 <= 1'b0; else if (n71) n409 <= n4423;
/* FF  9  3  6 */ assign n1094 = n4424;
/* FF  5 17  4 */ assign n771 = n4425;
/* FF  4 13  3 */ assign n4426 = n4427;
/* FF 11 12  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1473 <= 1'b0; else if (n102) n1473 <= n4428;
/* FF  2  5  6 */ always @(posedge io_13_31_1) if (n201) n35 <= n42 ? 1'b0 : n4429;
/* FF  3  1  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n342 <= 1'b0; else if (n500) n342 <= n4430;
/* FF 11 11  7 */ assign n892 = n4431;
/* FF 23 18  1 */ always @(posedge io_13_31_1) if (n2987) n3039 <= 1'b0 ? 1'b0 : n4432;
/* FF 14 11  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1933 <= 1'b0; else if (n734) n1933 <= n4433;
/* FF 15 15  6 */ always @(posedge io_13_31_1) if (n1180) n2131 <= n1 ? 1'b1 : n4434;
/* FF 15  7  2 */ assign n2060 = n4435;
/* FF  5 10  1 */ always @(posedge io_13_31_1) if (n4) n724 <= 1'b0 ? 1'b0 : n4436;
/* FF  7 21  3 */ assign n926 = n4437;
/* FF  8 17  1 */ assign n4438 = n4439;
/* FF 22  5  6 */ assign n2916 = n4440;
/* FF  5 13  6 */ assign n747 = n4441;
/* FF 21  1  5 */ assign n2757 = n4442;
/* FF  4  9  5 */ always @(posedge io_13_31_1) if (n4) n561 <= 1'b0 ? 1'b0 : n4443;
/* FF 15  8  3 */ assign n2071 = n4444;
/* FF 16 23  7 */ assign n2300 = n4445;
/* FF 17 19  5 */ assign n4446 = n4447;
/* FF 17 11  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2375 <= 1'b0; else if (n1764) n2375 <= n4448;
/* FF  7 14  0 */ assign n818 = n4449;
/* FF  2  6  6 */ assign n210 = n4450;
/* FF 14 12  4 */ assign n1945 = n4451;
/* FF 14  4  0 */ assign n1875 = n4452;
/* FF  1 19  0 */ assign n4453 = n4454;
/* FF  8 12  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1022 <= 1'b1; else if (n1166) n1022 <= n4456;
/* FF 10 21  4 */ assign n1389 = n4457;
/* FF 10 13  0 */ assign n1333 = n4458;
/* FF  9 17  3 */ assign n1201 = n4459;
/* FF 13 21  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1832 <= 1'b0; else if (n1830) n1832 <= n4460;
/* FF  7  9  6 */ assign n875 = n4461;
/* FF  8  5  4 */ assign n970 = n4462;
/* FF 21 23  1 */ always @(posedge io_13_31_1) if (n2879) n2878 <= 1'b0 ? 1'b0 : n4463;
/* FF 20 19  6 */ always @(posedge io_13_31_1) if (n2745) n2667 <= 1'b0 ? 1'b0 : n4464;
/* FF 20 11  2 */ always @(posedge io_13_31_1) if (n2137) n2697 <= n3 ? 1'b0 : n4465;
/* FF 10 14  1 */ assign n1342 = n4466;
/* FF 18 24  4 */ assign n2591 = n4467;
/* FF  9 18  4 */ assign n4468 = n4469;
/* FF  9 10  0 */ always @(posedge io_13_31_1) if (n4) n1151 <= 1'b0 ? 1'b0 : n4470;
/* FF 16  8  4 */ assign n2209 = n4471;
/* FF 13 13  3 */ always @(posedge io_13_31_1) if (1'b1) n1773 <= 1'b0 ? 1'b0 : n4472;
/* FF 20 12  3 */ assign n2664 = n4473;
/* FF  3 19  7 */ assign n473 = n4474;
/* FF 16  1  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n79 <= 1'b1; else if (1'b1) n79 <= n4475;
/* FF  2 20  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n318 <= 1'b0; else if (1'b1) n318 <= n4476;
/* FF 10  9  7 */ assign n1300 = n4477;
/* FF  9  5  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1113 <= 1'b0; else if (n840) n1113 <= n4478;
/* FF  1  8  4 */ assign n55 = n4479;
/* FF  3 11  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n425 <= 1'b1; else if (n70) n425 <= n4480;
/* FF 11 14  3 */ assign n1481 = n4481;
/* FF 12 18  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1644 <= 1'b0; else if (1'b1) n1644 <= n4482;
/* FF 12 10  1 */ assign n816 = n4483;
/* FF  2 13  0 */ assign n225 = n4484;
/* FF 10  2  4 */ assign n1246 = n4485;
/* FF  9  6  7 */ assign n891 = n4486;
/* FF 22 16  6 */ assign n2981 = n4487;
/* FF  2 16  5 */ assign n127 = n4488;
/* FF 13  9  4 */ assign n1745 = n4489;
/* FF 22  8  2 */ assign n2623 = n4490;
/* FF  3 12  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n45 <= 1'b1; else if (n98) n45 <= n4491;
/* FF 21 12  5 */ always @(posedge io_13_31_1) if (n2663) n2816 <= 1'b0 ? 1'b0 : n4492;
/* FF 21  4  1 */ always @(posedge io_13_31_1) if (n2902) n2769 <= n7 ? 1'b0 : n4493;
/* FF  1  4  6 */ always @(posedge io_13_31_1) if (n201) n33 <= n42 ? 1'b0 : n4494;
/* FF 15 18  1 */ assign n4495 = n4496;
/* FF 12 14  7 */ assign n1623 = n4497;
/* FF 18  5  4 */ always @(posedge io_13_31_1) if (n2456) n2461 <= 1'b0 ? 1'b0 : n4498;
/* FF  5 20  4 */ assign n794 = n4499;
/* FF  2  9  2 */ assign n239 = n4500;
/* FF 13  2  1 */ assign n1532 = n4501;
/* FF 11 15  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1490 <= 1'b0; else if (1'b1) n1490 <= n4502;
/* FF 14 23  4 */ assign n2034 = n4503;
/* FF  8 20  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1061 <= 1'b0; else if (n1062) n1061 <= n4504;
/* FF  2  8  6 */ assign n71 = n4505;
/* FF 13  1  5 */ assign n4506 = n4507;
/* FF 18  6  5 */ always @(posedge io_13_31_1) if (n2602) n2469 <= n1 ? 1'b0 : n4508;
/* FF 15 10  2 */ assign n1594 = n4509;
/* FF 21  5  1 */ always @(posedge io_13_31_1) if (n2902) n2777 <= n7 ? 1'b0 : n4510;
/* FF 15 13  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1965 <= 1'b0; else if (n735) n1965 <= n4511;
/* FF  5 16  6 */ assign n611 = n4512;
/* FF  4 12  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n582 <= 1'b0; else if (n432) n582 <= n4513;
/* FF 14 15  5 */ assign n1971 = n4514;
/* FF  8 16  4 */ assign n1045 = n4515;
/* FF 17 22  5 */ assign n2434 = n4516;
/* FF 23 13  2 */ always @(posedge io_13_31_1) if (n2842) n3017 <= 1'b0 ? 1'b0 : n4517;
/* FF 17 14  1 */ always @(posedge io_13_31_1) if (n2396) n2266 <= n1 ? 1'b0 : n4518;
/* FF 11  2  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1401 <= 1'b0; else if (n1120) n1401 <= n4519;
/* FF  7 17  0 */ assign n914 = n4520;
/* FF  5 17  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n773 <= 1'b0; else if (1'b1) n773 <= n4521;
/* FF 15  6  4 */ always @(posedge io_13_31_1) if (n2191) n1125 <= 1'b0 ? 1'b0 : n4522;
/* FF  2  1  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n162 <= 1'b0; else if (n178) n162 <= n4523;
/* FF  5  9  3 */ always @(posedge io_13_31_1) if (n4) n717 <= 1'b0 ? 1'b0 : n4524;
/* FF  4 13  6 */ assign n584 = n4525;
/* FF  4  5  2 */ assign n528 = n4526;
/* FF 14  7  0 */ assign n1905 = n4527;
/* FF 16 19  4 */ always @(posedge io_13_31_1) if (n1513) n2279 <= n1 ? 1'b0 : n4528;
/* FF 17 15  2 */ assign n2396 = n4529;
/* FF 11  3  6 */ assign n1406 = n4530;
/* FF 14 11  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1453 <= 1'b0; else if (n734) n1453 <= n4531;
/* FF 15  7  5 */ always @(posedge io_13_31_1) if (n1739) n1923 <= 1'b0 ? 1'b0 : n4532;
/* FF 20 22  7 */ assign n2727 = n4533;
/* FF 14  8  1 */ assign n1918 = n4534;
/* FF  9 20  3 */ assign n1215 = n4535;
/* FF  5  1  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n653 <= 1'b0; else if (n656) n653 <= n4536;
/* FF  7 12  6 */ assign n749 = n4537;
/* FF  8  8  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n989 <= 1'b0; else if (n877) n989 <= n4538;
/* FF 16 11  5 */ assign n2234 = n4539;
/* FF 23  2  1 */ assign n4540 = n4541;
/* FF 20 14  2 */ assign n2714 = n4542;
/* FF 10 17  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1369 <= 1'b0; else if (n1502) n1369 <= n4543;
/* FF  9 13  0 */ always @(posedge io_13_31_1) if (n4) n1172 <= 1'b0 ? 1'b0 : n4544;
/* FF  7 13  7 */ always @(posedge io_13_31_1) if (n4) n901 <= 1'b0 ? 1'b0 : n4545;
/* FF 17  2  4 */ always @(posedge io_13_31_1) if (n2324) n2309 <= 1'b0 ? 1'b0 : n4546;
/* FF  7  5  3 */ always @(posedge io_13_31_1) if (n4) n849 <= 1'b0 ? 1'b0 : n4547;
/* FF  8  1  1 */ assign n934 = n4548;
/* FF  9 16  5 */ assign n4549 = n4550;
/* FF  1 19  3 */ assign n137 = n4551;
/* FF 14  3  7 */ assign n1874 = n4552;
/* FF  8  4  6 */ assign n965 = n4553;
/* FF 16  7  7 */ assign n2203 = n4554;
/* FF 12 21  0 */ assign n4555 = n4556;
/* FF 17  3  5 */ assign n2321 = n4558;
/* FF 10 21  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1367 <= 1'b1; else if (1'b1) n1367 <= n4559;
/* FF 10 13  3 */ always @(posedge io_13_31_1) if (n4) n1336 <= 1'b0 ? 1'b0 : n4560;
/* FF  9 17  6 */ assign n911 = n4561;
/* FF  9  9  2 */ assign n1138 = n4562;
/* FF 21 23  4 */ assign n2879 = n4563;
/* FF  1  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n18 <= 1'b0; else if (n17) n18 <= n4564;
/* FF 13 12  5 */ assign n1762 = n4565;
/* FF 13  4  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1679 <= 1'b0; else if (n1433) n1679 <= n4566;
/* FF 18 16  3 */ always @(posedge io_13_31_1) if (n2011) n2553 <= 1'b0 ? 1'b0 : n4567;
/* FF 12 13  1 */ always @(posedge io_13_31_1) if (n4) n1611 <= 1'b0 ? 1'b0 : n4568;
/* FF 10  5  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1257 <= 1'b0; else if (n979) n1257 <= n4569;
/* FF  9  1  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1078 <= 1'b0; else if (n851) n1078 <= n4570;
/* FF  2 19  5 */ assign n322 = n4571;
/* FF 13 13  6 */ always @(posedge io_13_31_1) if (1'b1) n1776 <= 1'b0 ? 1'b0 : n4572;
/* FF 22 11  2 */ assign n2955 = n4573;
/* FF  2 11  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n252 <= 1'b0; else if (1'b1) n252 <= n4574;
/* FF  3 15  3 */ assign n441 = n4575;
/* FF 22 19  6 */ assign n2747 = n4576;
/* FF 21 15  5 */ assign n2841 = n4577;
/* FF 21  7  1 */ always @(posedge io_13_31_1) if (n2694) n2790 <= n1 ? 1'b0 : n4578;
/* FF  1  7  6 */ assign n50 = n4579;
/* FF 11 10  0 */ always @(posedge io_13_31_1) if (n4) n1455 <= 1'b0 ? 1'b0 : n4580;
/* FF 12 17  7 */ assign n1638 = n4581;
/* FF 18  8  4 */ assign n2076 = n4582;
/* FF  2 20  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n329 <= 1'b0; else if (1'b1) n329 <= n4583;
/* FF 12  9  3 */ assign n1586 = n4584;
/* FF  2 12  2 */ assign n260 = n4585;
/* FF 13  5  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1694 <= 1'b0; else if (n1279) n1694 <= n4586;
/* FF 21  8  2 */ assign n2800 = n4587;
/* FF 14 18  0 */ always @(posedge io_13_31_1) if (n1513) n1992 <= n1 ? 1'b0 : n4588;
/* FF 11 14  6 */ assign n1484 = n4589;
/* FF 18  1  1 */ assign n2439 = n4590;
/* FF  8 18  3 */ assign n1054 = n4591;
/* FF 12  2  0 */ assign n1537 = n4592;
/* FF 17 17  2 */ always @(posedge io_13_31_1) if (1'b1) n2403 <= 1'b0 ? 1'b0 : n4593;
/* FF 12  1  4 */ assign n4594 = n4595;
/* FF  5 19  6 */ assign n786 = n4596;
/* FF 22  8  5 */ assign n2936 = n4597;
/* FF  5 11  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n730 <= 1'b0; else if (n128) n730 <= n4598;
/* FF 21  4  4 */ always @(posedge io_13_31_1) if (n2902) n2772 <= n7 ? 1'b0 : n4599;
/* FF  4 15  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n587 <= 1'b0; else if (n451) n587 <= n4600;
/* FF  4  7  1 */ assign n59 = n4601;
/* FF  8 19  4 */ assign n4602 = n4603;
/* FF 14 10  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1892 <= 1'b0; else if (n734) n1892 <= n4604;
/* FF  8 11  0 */ always @(posedge io_13_31_1) if (n4) n1012 <= 1'b0 ? 1'b0 : n4605;
/* FF 11  6  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1429 <= 1'b0; else if (n1426) n1429 <= n4606;
/* FF  7 20  0 */ assign n4607 = n4608;
/* FF  5 20  7 */ assign n796 = n4610;
/* FF 15  9  4 */ assign n2081 = n4611;
/* FF  5 12  3 */ assign n736 = n4612;
/* FF  4  8  2 */ assign n549 = n4613;
/* FF 16 14  0 */ assign n2252 = n4614;
/* FF 17 18  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2410 <= 1'b0; else if (n2011) n2410 <= n4615;
/* FF 14 14  7 */ assign n1964 = n4616;
/* FF 15 10  5 */ assign n2089 = n4617;
/* FF 14  6  3 */ assign n1897 = n4618;
/* FF 15  2  1 */ assign n2044 = n4619;
/* FF  1 21  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n154 <= 1'b0; else if (n80) n154 <= n4620;
/* FF  5  5  0 */ assign n681 = n4621;
/* FF  7 16  2 */ assign n913 = n4622;
/* FF 16 15  1 */ always @(posedge io_13_31_1) if (n2268) n2259 <= 1'b0 ? 1'b0 : n4623;
/* FF  9 19  6 */ assign n1212 = n4624;
/* FF  1 14  0 */ assign n105 = n4625;
/* FF 10 20  1 */ assign n1379 = n4626;
/* FF  8  7  7 */ assign n982 = n4627;
/* FF 17  5  4 */ always @(posedge io_13_31_1) if (n2456) n2338 <= 1'b0 ? 1'b0 : n4628;
/* FF 20 13  5 */ always @(posedge io_13_31_1) if (n2663) n2711 <= 1'b0 ? 1'b0 : n4629;
/* FF  7  8  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n867 <= 1'b0; else if (1'b1) n867 <= n4630;
/* FF 13 23  4 */ assign n1858 = n4631;
/* FF 16 10  7 */ assign n2228 = n4632;
/* FF 17  6  5 */ assign n2193 = n4633;
/* FF 16  2  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2053 <= 1'b0; else if (n1552) n2053 <= n4634;
/* FF 10 16  3 */ always @(posedge io_13_31_1) if (n4) n1363 <= 1'b0 ? 1'b0 : n4635;
/* FF  9 20  6 */ assign n1218 = n4636;
/* FF  5  1  7 */ assign n655 = n4637;
/* FF  9 12  2 */ assign n902 = n4638;
/* FF  7  4  5 */ assign n845 = n4639;
/* FF 13 15  5 */ assign n1798 = n4640;
/* FF 20 14  5 */ always @(posedge io_13_31_1) if (n2137) n2717 <= n3 ? 1'b0 : n4641;
/* FF 20  6  1 */ always @(posedge io_13_31_1) if (n2676) n2677 <= n1 ? 1'b0 : n4642;
/* FF 10  9  0 */ always @(posedge io_13_31_1) if (n4) n1293 <= 1'b0 ? 1'b0 : n4643;
/* FF  1 10  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n74 <= 1'b1; else if (n70) n74 <= n4644;
/* FF 17  2  7 */ always @(posedge io_13_31_1) if (n2324) n2312 <= 1'b0 ? 1'b0 : n4645;
/* FF  1  2  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n11 <= 1'b0; else if (n17) n11 <= n4646;
/* FF 10  8  4 */ always @(posedge io_13_31_1) if (n4) n1286 <= 1'b0 ? 1'b0 : n4647;
/* FF  9  4  3 */ assign n1103 = n4648;
/* FF  2 14  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n280 <= 1'b0; else if (n269) n280 <= n4649;
/* FF 13  8  2 */ assign n1729 = n4650;
/* FF 18 12  0 */ always @(posedge io_13_31_1) if (n2137) n2521 <= n3 ? 1'b0 : n4651;
/* FF 13 11  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1593 <= 1'b0; else if (n734) n1593 <= n4652;
/* FF 11 16  5 */ assign n1500 = n4653;
/* FF 10  1  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1235 <= 1'b0; else if (n1120) n1235 <= n4654;
/* FF 12 12  3 */ assign n1601 = n4655;
/* FF 22 15  3 */ always @(posedge io_13_31_1) if (1'b1) n2973 <= n3025 ? 1'b0 : n4656;
/* FF  2 15  2 */ assign n276 = n4657;
/* FF 10  4  6 */ assign n1261 = n4658;
/* FF  1  3  3 */ assign n21 = n4659;
/* FF  2 18  7 */ assign n314 = n4660;
/* FF 14 21  0 */ assign n2018 = n4661;
/* FF 13  4  4 */ assign n1684 = n4662;
/* FF 21 14  7 */ always @(posedge io_13_31_1) if (n2842) n2836 <= 1'b0 ? 1'b0 : n4663;
/* FF 11 17  6 */ assign n1506 = n4664;
/* FF 11  9  2 */ assign n1448 = n4665;
/* FF 12 13  4 */ always @(posedge io_13_31_1) if (n4) n1319 <= 1'b0 ? 1'b0 : n4666;
/* FF 12  5  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1435 <= 1'b0; else if (n1426) n1435 <= n4667;
/* FF  3  6  7 */ assign n388 = n4668;
/* FF 10  5  7 */ assign n1266 = n4669;
/* FF  4 19  1 */ assign n624 = n4670;
/* FF  9  1  6 */ assign n1081 = n4671;
/* FF 14 22  1 */ assign n2027 = n4672;
/* FF  2 11  4 */ assign n61 = n4673;
/* FF  4 18  5 */ assign n4674 = n4675;
/* FF 21  7  4 */ assign n2792 = n4676;
/* FF  8 14  0 */ assign n1035 = n4677;
/* FF 18  8  7 */ always @(posedge io_13_31_1) if (n2120) n2491 <= 1'b0 ? 1'b0 : n4678;
/* FF  5 15  3 */ assign n760 = n4679;
/* FF 17 16  4 */ assign n2400 = n4680;
/* FF  4 11  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n264 <= 1'b0; else if (1'b1) n264 <= n4681;
/* FF  8 15  1 */ assign n4682 = n4683;
/* FF  2  3  5 */ assign n185 = n4684;
/* FF 22  3  6 */ always @(posedge io_13_31_1) if (1'b1) n2899 <= n2757 ? 1'b1 : n4685;
/* FF  4 14  7 */ assign n596 = n4686;
/* FF 16 17  0 */ assign n2277 = n4687;
/* FF  8 18  6 */ assign n1034 = n4688;
/* FF 14  9  3 */ always @(posedge io_13_31_1) if (n1739) n1929 <= 1'b0 ? 1'b0 : n4689;
/* FF 15  5  1 */ assign n1902 = n4690;
/* FF  5  8  0 */ always @(posedge io_13_31_1) if (n4) n702 <= 1'b0 ? 1'b0 : n4691;
/* FF 17 17  5 */ always @(posedge io_13_31_1) if (1'b1) n2407 <= 1'b0 ? 1'b0 : n4692;
/* FF 12  1  7 */ assign n4693 = n4694;
/* FF 16 18  1 */ always @(posedge io_13_31_1) if (n1513) n2142 <= n1 ? 1'b0 : n4695;
/* FF  4  7  4 */ assign n232 = n4696;
/* FF 14 10  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1926 <= 1'b0; else if (n734) n1926 <= n4697;
/* FF 14  2  0 */ assign n1550 = n4698;
/* FF 16 21  6 */ always @(posedge io_13_31_1) if (n2038) n2291 <= 1'b0 ? 1'b0 : n4699;
/* FF  1 17  0 */ assign n4700 = n4701;
/* FF 23  8  1 */ always @(posedge io_13_31_1) if (1'b1) n3015 <= 1'b0 ? 1'b0 : n4703;
/* FF 17  9  0 */ always @(posedge io_13_31_1) if (n1591) n2356 <= 1'b0 ? 1'b0 : n4704;
/* FF  8 10  7 */ always @(posedge io_13_31_1) if (n4) n1011 <= 1'b0 ? 1'b0 : n4705;
/* FF  8  2  3 */ assign n943 = n4706;
/* FF  1 20  5 */ assign n147 = n4707;
/* FF 10 19  4 */ assign n1375 = n4708;
/* FF 10 11  0 */ always @(posedge io_13_31_1) if (n4) n1310 <= 1'b0 ? 1'b0 : n4709;
/* FF  5  3  6 */ assign n669 = n4710;
/* FF  9 15  3 */ always @(posedge io_13_31_1) if (n4) n1192 <= 1'b0 ? 1'b0 : n4711;
/* FF 17  4  7 */ always @(posedge io_13_31_1) if (n2316) n2332 <= 1'b0 ? 1'b0 : n4712;
/* FF 13 18  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1651 <= 1'b0; else if (n1967) n1651 <= n4713;
/* FF  8  3  4 */ assign n952 = n4714;
/* FF  1 21  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n156 <= 1'b0; else if (n80) n156 <= n4715;
/* FF 16 13  7 */ assign n2122 = n4716;
/* FF 16  5  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1700 <= 1'b0; else if (n1869) n1700 <= n4717;
/* FF  1 13  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n95 <= 1'b0; else if (n105) n95 <= n4718;
/* FF 17  1  1 */ assign n2303 = n4719;
/* FF 20  9  2 */ always @(posedge io_13_31_1) if (n2093) n2372 <= 1'b0 ? 1'b0 : n4720;
/* FF 18 22  4 */ assign n2582 = n4721;
/* FF 18 14  0 */ assign n2133 = n4722;
/* FF 13 19  1 */ assign n1816 = n4723;
/* FF  7  7  5 */ assign n858 = n4724;
/* FF 21 21  0 */ always @(posedge io_13_31_1) if (n2873) n2870 <= 1'b0 ? 1'b0 : n4725;
/* FF 16  6  4 */ assign n2187 = n4726;
/* FF 10 12  0 */ assign n1320 = n4727;
/* FF  3 13  0 */ assign n4728 = n4729;
/* FF 17  5  7 */ always @(posedge io_13_31_1) if (n2456) n2190 <= 1'b0 ? 1'b0 : n4731;
/* FF  1  5  3 */ assign n37 = n4732;
/* FF  3 16  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n303 <= 1'b0; else if (1'b1) n303 <= n4733;
/* FF 18 18  6 */ assign n2564 = n4734;
/* FF 12 15  4 */ assign n1630 = n4735;
/* FF 10  7  7 */ always @(posedge io_13_31_1) if (n4) n1278 <= 1'b0 ? 1'b0 : n4736;
/* FF  4 21  1 */ assign n4737 = n4738;
/* FF 16  2  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1931 <= 1'b0; else if (n1552) n1931 <= n4739;
/* FF 13 14  7 */ assign n1788 = n4740;
/* FF  3 17  6 */ assign n454 = n4741;
/* FF  3  9  2 */ assign n415 = n4742;
/* FF 18 10  7 */ always @(posedge io_13_31_1) if (n2120) n2508 <= 1'b0 ? 1'b0 : n4743;
/* FF  9  3  5 */ assign n1096 = n4744;
/* FF 12 11  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1598 <= 1'b0; else if (n734) n1598 <= n4745;
/* FF 13  7  4 */ assign n1722 = n4746;
/* FF 21 17  7 */ always @(posedge io_13_31_1) if (n2735) n2853 <= 1'b0 ? 1'b0 : n4747;
/* FF 11 20  6 */ assign n1390 = n4748;
/* FF  1  2  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n13 <= 1'b0; else if (n17) n13 <= n4749;
/* FF 12  8  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1271 <= 1'b0; else if (n1430) n1271 <= n4750;
/* FF 15 16  1 */ assign n4751 = n4752;
/* FF 10  8  7 */ assign n1289 = n4753;
/* FF  9  4  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1105 <= 1'b0; else if (n840) n1105 <= n4754;
/* FF 22 14  5 */ assign n4755 = n4756;
/* FF  2 14  4 */ assign n269 = n4757;
/* FF 22  6  1 */ always @(posedge io_13_31_1) if (1'b1) n354 <= 1'b0 ? 1'b0 : n4758;
/* FF 11 13  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n819 <= 1'b0; else if (n1461) n819 <= n4759;
/* FF 21  2  0 */ assign n2761 = n4760;
/* FF  8 17  0 */ assign n4761 = n4762;
/* FF 23 19  1 */ assign n2877 = n4764;
/* FF 12  4  2 */ assign n1539 = n4765;
/* FF 15  8  2 */ assign n2070 = n4766;
/* FF 22  7  2 */ always @(posedge io_13_31_1) if (n2694) n2690 <= n1 ? 1'b0 : n4767;
/* FF 17 19  4 */ assign n2421 = n4768;
/* FF 15 11  7 */ always @(posedge io_13_31_1) if (n2112) n2101 <= 1'b0 ? 1'b0 : n4769;
/* FF  2  6  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n52 <= 1'b0; else if (n217) n52 <= n4770;
/* FF  5 14  6 */ assign n604 = n4771;
/* FF  8 21  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n932 <= 1'b0; else if (n1068) n932 <= n4772;
/* FF 14 12  3 */ assign n1944 = n4773;
/* FF 17 20  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2427 <= 1'b0; else if (n2023) n2427 <= n4774;
/* FF 17 12  1 */ assign n2191 = n4775;
/* FF 15  4  4 */ assign n2050 = n4776;
/* FF 23 14  7 */ assign n2819 = n4777;
/* FF  5  6  1 */ assign n686 = n4778;
/* FF 14 13  4 */ assign n1952 = n4779;
/* FF  4  2  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n501 <= 1'b0; else if (n509) n501 <= n4780;
/* FF  8 14  3 */ assign n1038 = n4781;
/* FF  2  2  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n174 <= 1'b0; else if (n178) n174 <= n4782;
/* FF 14  5  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1885 <= 1'b0; else if (n1433) n1885 <= n4783;
/* FF 16 16  2 */ always @(posedge io_13_31_1) if (1'b1) n2272 <= 1'b0 ? 1'b0 : n4784;
/* FF 13 21  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1831 <= 1'b0; else if (n1830) n1831 <= n4785;
/* FF  8 13  7 */ assign n1030 = n4786;
/* FF 11  1  6 */ assign n4787 = n4788;
/* FF  5  7  2 */ assign n372 = n4789;
/* FF  4  3  1 */ assign n511 = n4790;
/* FF  9 18  3 */ assign n4791 = n4792;
/* FF 16 17  3 */ assign n2278 = n4793;
/* FF  7  2  2 */ assign n831 = n4794;
/* FF  8  6  4 */ assign n712 = n4795;
/* FF  1 16  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n120 <= 1'b0; else if (n127) n120 <= n4796;
/* FF 20 20  6 */ assign n2745 = n4797;
/* FF 10 15  1 */ always @(posedge io_13_31_1) if (n4) n1353 <= 1'b0 ? 1'b0 : n4798;
/* FF 13 22  1 */ assign n1842 = n4799;
/* FF 10 18  6 */ assign n4800 = n4801;
/* FF  9 14  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1185 <= 1'b0; else if (n762) n1185 <= n4802;
/* FF  8  2  6 */ assign n361 = n4803;
/* FF 16  4  5 */ always @(posedge io_13_31_1) if (n2324) n2176 <= 1'b0 ? 1'b0 : n4804;
/* FF 12 19  0 */ assign n1646 = n4805;
/* FF  7  3  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n835 <= 1'b0; else if (n663) n835 <= n4806;
/* FF 10 11  3 */ assign n1313 = n4807;
/* FF 16  5  6 */ assign n2180 = n4808;
/* FF  2 16  4 */ assign n295 = n4809;
/* FF  3 20  6 */ assign n480 = n4810;
/* FF 13  9  3 */ assign n1744 = n4811;
/* FF  3 12  2 */ assign n432 = n4812;
/* FF 18 14  3 */ assign n2536 = n4813;
/* FF  1  4  5 */ assign n32 = n4814;
/* FF 15 18  0 */ assign n4815 = n4816;
/* FF 12 14  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1622 <= 1'b0; else if (n1630) n1622 <= n4818;
/* FF 22 17  6 */ assign n2737 = n4819;
/* FF  2 17  5 */ assign n257 = n4820;
/* FF 13 10  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1434 <= 1'b0; else if (n734) n1434 <= n4821;
/* FF  2  9  1 */ assign n238 = n4822;
/* FF  3 13  3 */ assign n4823 = n4824;
/* FF 13  2  0 */ assign n1423 = n4825;
/* FF 11 15  2 */ assign n1489 = n4826;
/* FF  1  5  6 */ assign n39 = n4827;
/* FF 14 23  3 */ assign n2033 = n4828;
/* FF 15 19  1 */ assign n4829 = n4830;
/* FF 10  3  3 */ assign n959 = n4831;
/* FF 12 15  7 */ always @(posedge io_13_31_1) if (n1180) n1366 <= n1 ? 1'b0 : n4832;
/* FF 18  6  4 */ always @(posedge io_13_31_1) if (n2602) n2468 <= n1 ? 1'b0 : n4833;
/* FF 12  7  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1570 <= 1'b0; else if (n1279) n1570 <= n4834;
/* FF 13  3  1 */ assign n1672 = n4835;
/* FF 21 13  4 */ assign n2822 = n4836;
/* FF  4 21  4 */ assign n4837 = n4838;
/* FF 21  5  0 */ always @(posedge io_13_31_1) if (n2902) n2776 <= n7 ? 1'b0 : n4839;
/* FF  8 16  3 */ assign n920 = n4840;
/* FF 21  6  1 */ always @(posedge io_13_31_1) if (n2686) n2601 <= 1'b0 ? 1'b0 : n4841;
/* FF 18  2  6 */ always @(posedge io_13_31_1) if (n2456) n2171 <= 1'b0 ? 1'b0 : n4842;
/* FF 15 14  7 */ assign n2127 = n4843;
/* FF  5  9  2 */ always @(posedge io_13_31_1) if (n4) n716 <= 1'b0 ? 1'b0 : n4844;
/* FF  4 13  5 */ assign n585 = n4845;
/* FF 11  4  1 */ assign n1411 = n4846;
/* FF  4  5  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n527 <= 1'b0; else if (n524) n527 <= n4847;
/* FF  3  1  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n344 <= 1'b0; else if (n500) n344 <= n4848;
/* FF 16 19  3 */ assign n4849 = n4850;
/* FF 17 15  1 */ assign n2138 = n4851;
/* FF 11  3  5 */ assign n1405 = n4852;
/* FF 14 11  6 */ assign n1764 = n4853;
/* FF  7 18  0 */ assign n4854 = n4855;
/* FF 15  7  4 */ assign n2062 = n4857;
/* FF 23 17  7 */ assign n2856 = n4858;
/* FF  5 10  3 */ assign n726 = n4859;
/* FF  7 21  5 */ assign n927 = n4860;
/* FF  8 17  3 */ assign n4861 = n4862;
/* FF 14  8  0 */ assign n1917 = n4863;
/* FF  4  9  7 */ assign n563 = n4864;
/* FF 15  8  5 */ assign n2073 = n4865;
/* FF 17 19  7 */ assign n4866 = n4867;
/* FF 17 11  3 */ assign n2376 = n4868;
/* FF 23  2  0 */ assign n4869 = n4870;
/* FF  4  6  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n537 <= 1'b0; else if (n532) n537 <= n4872;
/* FF  7 14  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n904 <= 1'b0; else if (1'b1) n904 <= n4873;
/* FF 16 20  3 */ assign n2022 = n4874;
/* FF  7 13  6 */ always @(posedge io_13_31_1) if (n4) n900 <= 1'b0 ? 1'b0 : n4875;
/* FF 14 12  6 */ assign n1947 = n4876;
/* FF 14  4  2 */ assign n1878 = n4877;
/* FF  8  1  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n933 <= 1'b0; else if (n656) n933 <= n4878;
/* FF  1 19  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n136 <= 1'b0; else if (n140) n136 <= n4879;
/* FF 23  3  1 */ assign n4880 = n4881;
/* FF  8  4  5 */ assign n947 = n4882;
/* FF 20 18  7 */ assign n2734 = n4883;
/* FF 17  3  4 */ always @(posedge io_13_31_1) if (n2324) n2320 <= 1'b0 ? 1'b0 : n4884;
/* FF 10 13  2 */ always @(posedge io_13_31_1) if (n4) n1335 <= 1'b0 ? 1'b0 : n4885;
/* FF  9 17  5 */ assign n1203 = n4886;
/* FF  9  9  1 */ always @(posedge io_13_31_1) if (n4) n1137 <= 1'b0 ? 1'b0 : n4887;
/* FF 13 21  4 */ assign n1527 = n4888;
/* FF  8  5  6 */ assign n808 = n4889;
/* FF 12 22  0 */ assign n4890 = n4891;
/* FF 20 11  4 */ always @(posedge io_13_31_1) if (n2137) n2699 <= n3 ? 1'b0 : n4893;
/* FF 10 14  3 */ always @(posedge io_13_31_1) if (n4) n1344 <= 1'b0 ? 1'b0 : n4894;
/* FF  9 18  6 */ assign n4895 = n4896;
/* FF  9 10  2 */ assign n1153 = n4897;
/* FF 22 20  1 */ always @(posedge io_13_31_1) if (n2998) n2996 <= 1'b0 ? 1'b0 : n4898;
/* FF  7  2  5 */ assign n832 = n4899;
/* FF 21 16  0 */ assign n2843 = n4900;
/* FF 16  8  6 */ assign n2211 = n4901;
/* FF 13 13  5 */ always @(posedge io_13_31_1) if (1'b1) n1775 <= 1'b0 ? 1'b0 : n4902;
/* FF  3 15  2 */ assign n440 = n4903;
/* FF 20  4  1 */ assign n2670 = n4904;
/* FF 18 17  3 */ assign n2559 = n4905;
/* FF  1  7  5 */ assign n49 = n4906;
/* FF 12 17  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1609 <= 1'b0; else if (1'b1) n1609 <= n4907;
/* FF  2 20  5 */ assign n159 = n4908;
/* FF 22 12  2 */ assign n2957 = n4909;
/* FF  2 12  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n261 <= 1'b0; else if (1'b1) n261 <= n4910;
/* FF 13  5  0 */ assign n1693 = n4911;
/* FF 21  8  1 */ assign n4912 = n4913;
/* FF  1  8  6 */ assign n57 = n4914;
/* FF 11 14  5 */ assign n1483 = n4915;
/* FF 12 18  7 */ assign n1639 = n4916;
/* FF  2 13  2 */ assign n274 = n4917;
/* FF 13  6  1 */ assign n1708 = n4918;
/* FF 10  2  6 */ assign n1098 = n4919;
/* FF  4 16  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n455 <= 1'b0; else if (1'b1) n455 <= n4920;
/* FF  2 16  7 */ assign n291 = n4921;
/* FF 13  9  6 */ assign n1747 = n4922;
/* FF 14 19  0 */ assign n4923 = n4924;
/* FF  3 12  5 */ assign n428 = n4926;
/* FF 21 12  7 */ always @(posedge io_13_31_1) if (n2663) n2810 <= 1'b0 ? 1'b0 : n4927;
/* FF 22  8  4 */ assign n2940 = n4928;
/* FF  3  4  1 */ assign n364 = n4929;
/* FF 21  4  3 */ always @(posedge io_13_31_1) if (n2902) n2771 <= n7 ? 1'b0 : n4930;
/* FF 15 18  3 */ assign n4931 = n4932;
/* FF  8 19  3 */ assign n4933 = n4934;
/* FF 12  3  0 */ assign n4935 = n4936;
/* FF 18  5  6 */ always @(posedge io_13_31_1) if (n2456) n2463 <= 1'b0 ? 1'b0 : n4938;
/* FF  5 20  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n620 <= 1'b0; else if (n629) n620 <= n4939;
/* FF 17 21  7 */ assign n2432 = n4940;
/* FF 11 15  5 */ assign n1492 = n4941;
/* FF 11  7  1 */ assign n1430 = n4942;
/* FF  8 20  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1043 <= 1'b0; else if (n1062) n1043 <= n4943;
/* FF 13  1  7 */ assign n4944 = n4945;
/* FF 17 18  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2409 <= 1'b0; else if (n2011) n2409 <= n4946;
/* FF 14 14  6 */ assign n1963 = n4947;
/* FF 15 10  4 */ assign n2088 = n4948;
/* FF 15  2  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1883 <= 1'b0; else if (n1552) n1883 <= n4949;
/* FF  7 16  1 */ assign n912 = n4950;
/* FF 16 15  0 */ always @(posedge io_13_31_1) if (n2268) n2258 <= 1'b0 ? 1'b0 : n4951;
/* FF 14 15  7 */ assign n1972 = n4952;
/* FF  8 16  6 */ assign n921 = n4953;
/* FF 15  3  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1595 <= 1'b0; else if (n1547) n1595 <= n4954;
/* FF 17 14  3 */ always @(posedge io_13_31_1) if (n2396) n2392 <= n1 ? 1'b0 : n4955;
/* FF  7 17  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n614 <= 1'b0; else if (n916) n614 <= n4956;
/* FF 15  6  6 */ assign n2057 = n4957;
/* FF  2  1  4 */ assign n163 = n4958;
/* FF  5  9  5 */ always @(posedge io_13_31_1) if (n4) n719 <= 1'b0 ? 1'b0 : n4959;
/* FF  4  5  4 */ assign n525 = n4960;
/* FF 14  7  2 */ assign n1907 = n4961;
/* FF 16 19  6 */ always @(posedge io_13_31_1) if (n1513) n2280 <= n1 ? 1'b0 : n4962;
/* FF 13 23  3 */ assign n1857 = n4963;
/* FF 17  7  0 */ assign n4964 = n4965;
/* FF  1 18  5 */ assign n118 = n4966;
/* FF 17  6  4 */ assign n4967 = n4968;
/* FF 10 16  2 */ assign n1362 = n4969;
/* FF  9 20  5 */ assign n1217 = n4970;
/* FF  9 12  1 */ assign n1024 = n4971;
/* FF 13 16  0 */ assign n1802 = n4972;
/* FF  7  4  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n371 <= 1'b0; else if (n224) n371 <= n4973;
/* FF  8  8  6 */ assign n990 = n4974;
/* FF 16 11  7 */ always @(posedge io_13_31_1) if (n2076) n2236 <= 1'b0 ? 1'b0 : n4975;
/* FF 23  2  3 */ assign n3006 = n4976;
/* FF 16  3  3 */ assign n1534 = n4977;
/* FF 20 14  4 */ always @(posedge io_13_31_1) if (n2137) n2716 <= n3 ? 1'b0 : n4978;
/* FF 20  6  0 */ assign n4979 = n4980;
/* FF  9 13  2 */ always @(posedge io_13_31_1) if (n4) n1174 <= 1'b0 ? 1'b0 : n4982;
/* FF 17  2  6 */ assign n2311 = n4983;
/* FF 22 23  1 */ assign n3004 = n4984;
/* FF 13 17  1 */ assign n4985 = n4986;
/* FF  7  5  5 */ assign n850 = n4987;
/* FF  8  1  3 */ assign n936 = n4988;
/* FF  9 16  7 */ assign n4989 = n4990;
/* FF 20 15  5 */ assign n2722 = n4991;
/* FF 20  7  1 */ assign n4992 = n4993;
/* FF 10 10  0 */ always @(posedge io_13_31_1) if (n4) n1302 <= 1'b0 ? 1'b0 : n4994;
/* FF 18 20  3 */ always @(posedge io_13_31_1) if (n1837) n2581 <= 1'b0 ? 1'b0 : n4995;
/* FF 12 21  2 */ assign n1656 = n4996;
/* FF 17  3  7 */ always @(posedge io_13_31_1) if (n2324) n2323 <= 1'b0 ? 1'b0 : n4997;
/* FF  3 14  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n80 <= 1'b0; else if (1'b1) n80 <= n4998;
/* FF 10 13  5 */ always @(posedge io_13_31_1) if (n4) n1331 <= 1'b0 ? 1'b0 : n4999;
/* FF  9  9  4 */ always @(posedge io_13_31_1) if (n4) n1140 <= 1'b0 ? 1'b0 : n5000;
/* FF  2 15  1 */ assign n287 = n5001;
/* FF 18 13  0 */ always @(posedge io_13_31_1) if (n2137) n2528 <= n3 ? 1'b0 : n5002;
/* FF  1  3  2 */ assign n20 = n5003;
/* FF 13 12  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1763 <= 1'b0; else if (n755) n1763 <= n5004;
/* FF  2 18  6 */ assign n305 = n5005;
/* FF 13  4  3 */ assign n1683 = n5006;
/* FF 11 17  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1479 <= 1'b0; else if (n762) n1479 <= n5007;
/* FF 18 16  5 */ always @(posedge io_13_31_1) if (n2011) n2555 <= 1'b0 ? 1'b0 : n5008;
/* FF 12 13  3 */ always @(posedge io_13_31_1) if (n4) n1470 <= 1'b0 ? 1'b0 : n5009;
/* FF  4 19  0 */ assign n623 = n5010;
/* FF  9  1  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1080 <= 1'b0; else if (n851) n1080 <= n5011;
/* FF  2 19  7 */ assign n134 = n5012;
/* FF 14 22  0 */ assign n2026 = n5013;
/* FF 22 11  4 */ assign n2250 = n5014;
/* FF  2 11  3 */ assign n254 = n5015;
/* FF  3 15  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n442 <= 1'b0; else if (1'b1) n442 <= n5016;
/* FF  3  7  1 */ assign n397 = n5017;
/* FF 11 18  6 */ always @(posedge io_13_31_1) if (1'b1) n1512 <= 1'b0 ? 1'b0 : n5018;
/* FF 21  7  3 */ assign n5019 = n5020;
/* FF 11 10  2 */ assign n1457 = n5021;
/* FF 12  6  0 */ assign n1292 = n5022;
/* FF 24 20  2 */ always @(posedge io_13_31_1) if (n2876) n2999 <= 1'b0 ? 1'b0 : n5023;
/* FF  4 20  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n488 <= 1'b0; else if (n629) n488 <= n5024;
/* FF 18  8  6 */ always @(posedge io_13_31_1) if (n2120) n2490 <= 1'b0 ? 1'b0 : n5025;
/* FF 12  9  5 */ assign n1588 = n5026;
/* FF  2 12  4 */ assign n262 = n5027;
/* FF 13  5  3 */ assign n1574 = n5028;
/* FF 22  4  1 */ assign n2910 = n5029;
/* FF  2  4  0 */ always @(posedge io_13_31_1) if (n201) n192 <= n42 ? 1'b0 : n5030;
/* FF 21  8  4 */ always @(posedge io_13_31_1) if (n2694) n2801 <= n1 ? 1'b0 : n5031;
/* FF 14 18  2 */ assign n1994 = n5032;
/* FF  8 15  0 */ assign n5033 = n5034;
/* FF 18  1  3 */ assign n2441 = n5036;
/* FF  8 18  5 */ assign n1056 = n5037;
/* FF 17 17  4 */ always @(posedge io_13_31_1) if (1'b1) n2406 <= 1'b0 ? 1'b0 : n5038;
/* FF  7 19  1 */ assign n822 = n5039;
/* FF 12  1  6 */ assign n5040 = n5041;
/* FF  5 11  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n583 <= 1'b0; else if (n128) n583 <= n5042;
/* FF  4 15  7 */ assign n589 = n5043;
/* FF 16 18  0 */ assign n5044 = n5045;
/* FF 23 17  0 */ always @(posedge io_13_31_1) if (n2985) n3038 <= 1'b0 ? 1'b0 : n5047;
/* FF  4  7  3 */ assign n543 = n5048;
/* FF  8 19  6 */ assign n5049 = n5050;
/* FF 14 10  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1463 <= 1'b0; else if (n734) n1463 <= n5051;
/* FF  8 11  2 */ always @(posedge io_13_31_1) if (n4) n1014 <= 1'b0 ? 1'b0 : n5052;
/* FF  7 20  2 */ assign n5053 = n5054;
/* FF 15  9  6 */ assign n2083 = n5055;
/* FF  5 12  5 */ assign n737 = n5056;
/* FF  5  4  1 */ assign n673 = n5057;
/* FF  4  8  4 */ always @(posedge io_13_31_1) if (n4) n551 <= 1'b0 ? 1'b0 : n5058;
/* FF 16 22  6 */ always @(posedge io_13_31_1) if (n2294) n2295 <= 1'b0 ? 1'b0 : n5059;
/* FF 16 14  2 */ always @(posedge io_13_31_1) if (1'b1) n1807 <= n2253 ? 1'b0 : n5060;
/* FF 17 18  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2412 <= 1'b0; else if (n2011) n2412 <= n5061;
/* FF 17 10  0 */ assign n5062 = n5063;
/* FF 14  6  5 */ assign n1899 = n5065;
/* FF  8  3  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n951 <= 1'b0; else if (n840) n951 <= n5066;
/* FF  1 21  5 */ assign n155 = n5067;
/* FF 15  2  3 */ assign n2045 = n5068;
/* FF  1 13  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n94 <= 1'b0; else if (n105) n94 <= n5069;
/* FF 20 17  5 */ assign n2726 = n5070;
/* FF 13 19  0 */ assign n5071 = n5072;
/* FF 23 13  7 */ assign n3018 = n5074;
/* FF 16  6  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1731 <= 1'b0; else if (n1433) n1731 <= n5075;
/* FF 17  5  6 */ always @(posedge io_13_31_1) if (n2456) n2339 <= 1'b0 ? 1'b0 : n5076;
/* FF 20 13  7 */ always @(posedge io_13_31_1) if (n2663) n2713 <= 1'b0 ? 1'b0 : n5077;
/* FF 13 20  1 */ assign n5078 = n5079;
/* FF  7  8  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n869 <= 1'b0; else if (1'b1) n869 <= n5080;
/* FF 13 23  6 */ assign n1849 = n5081;
/* FF 20 10  1 */ assign n2112 = n5082;
/* FF  3 18  1 */ assign n459 = n5083;
/* FF 17  6  7 */ assign n2340 = n5084;
/* FF 16  2  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1716 <= 1'b0; else if (n1552) n1716 <= n5085;
/* FF  7  1  2 */ assign n824 = n5086;
/* FF  9 12  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1169 <= 1'b0; else if (n818) n1169 <= n5087;
/* FF  7  4  7 */ assign n847 = n5088;
/* FF  4 22  1 */ assign n481 = n5089;
/* FF 16  3  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1932 <= 1'b0; else if (n1690) n1932 <= n5090;
/* FF 11 21  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1521 <= 1'b0; else if (1'b1) n1521 <= n5091;
/* FF 13 15  7 */ always @(posedge io_13_31_1) if (1'b1) n1800 <= 1'b0 ? 1'b0 : n5092;
/* FF 13  7  3 */ assign n1721 = n5093;
/* FF 20  6  3 */ always @(posedge io_13_31_1) if (n2676) n2679 <= n1 ? 1'b0 : n5094;
/* FF 18 11  1 */ assign n2513 = n5095;
/* FF 15 16  0 */ assign n5096 = n5097;
/* FF 10  8  6 */ always @(posedge io_13_31_1) if (n4) n1288 <= 1'b0 ? 1'b0 : n5099;
/* FF  9  4  5 */ assign n1099 = n5100;
/* FF 22 14  4 */ assign n2968 = n5101;
/* FF  2 14  3 */ assign n282 = n5102;
/* FF 13  8  4 */ assign n1735 = n5103;
/* FF 10  1  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1237 <= 1'b0; else if (n1120) n1237 <= n5104;
/* FF 11 16  7 */ assign n1502 = n5105;
/* FF 12 12  5 */ always @(posedge io_13_31_1) if (n4) n1599 <= 1'b0 ? 1'b0 : n5106;
/* FF 18  3  2 */ always @(posedge io_13_31_1) if (n2191) n852 <= 1'b0 ? 1'b0 : n5107;
/* FF 22 15  5 */ assign n2975 = n5108;
/* FF  2 15  4 */ assign n289 = n5109;
/* FF 12  4  1 */ assign n1543 = n5110;
/* FF 22  7  1 */ assign n2694 = n5111;
/* FF  2  7  0 */ assign n217 = n5112;
/* FF 21 11  4 */ always @(posedge io_13_31_1) if (n2213) n2501 <= 1'b0 ? 1'b0 : n5113;
/* FF 24 18  3 */ always @(posedge io_13_31_1) if (n2862) n2994 <= 1'b0 ? 1'b0 : n5114;
/* FF 21  3  0 */ assign n5115 = n5116;
/* FF 15 17  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1822 <= 1'b0; else if (n1815) n1822 <= n5118;
/* FF 13  4  6 */ assign n1686 = n5119;
/* FF 17 21  0 */ assign n2428 = n5120;
/* FF 11  9  4 */ always @(posedge io_13_31_1) if (n4) n1449 <= 1'b0 ? 1'b0 : n5121;
/* FF  8 21  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1019 <= 1'b0; else if (n1068) n1019 <= n5122;
/* FF 12  5  2 */ assign n1318 = n5123;
/* FF 17 20  4 */ assign n2023 = n5124;
/* FF 15 12  7 */ assign n2109 = n5125;
/* FF  4 18  7 */ assign n5126 = n5127;
/* FF 21  7  6 */ assign n2793 = n5128;
/* FF  4 10  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n566 <= 1'b0; else if (n576) n566 <= n5129;
/* FF 14 13  3 */ assign n1951 = n5130;
/* FF  8 14  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1037 <= 1'b0; else if (n754) n1037 <= n5131;
/* FF  2  2  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n173 <= 1'b0; else if (n178) n173 <= n5132;
/* FF 11  1  5 */ assign n5133 = n5134;
/* FF  5 15  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n750 <= 1'b0; else if (n451) n750 <= n5135;
/* FF  5  7  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n692 <= 1'b0; else if (n532) n692 <= n5136;
/* FF 17 16  6 */ always @(posedge io_13_31_1) if (n2268) n2401 <= 1'b0 ? 1'b0 : n5137;
/* FF  4 11  4 */ assign n243 = n5138;
/* FF  4  3  0 */ assign n510 = n5139;
/* FF  8 15  3 */ assign n5140 = n5141;
/* FF  2  3  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n187 <= 1'b0; else if (n17) n187 <= n5142;
/* FF 17 13  0 */ assign n5143 = n5144;
/* FF 14  9  5 */ always @(posedge io_13_31_1) if (n1739) n1756 <= 1'b0 ? 1'b0 : n5146;
/* FF 15  5  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1877 <= 1'b0; else if (n1869) n1877 <= n5147;
/* FF  5  8  2 */ always @(posedge io_13_31_1) if (n4) n704 <= 1'b0 ? 1'b0 : n5148;
/* FF 17 17  7 */ always @(posedge io_13_31_1) if (1'b1) n2408 <= 1'b0 ? 1'b0 : n5149;
/* FF  7 19  4 */ assign n923 = n5150;
/* FF  4  4  1 */ assign n520 = n5151;
/* FF  7 11  0 */ always @(posedge io_13_31_1) if (n4) n881 <= 1'b0 ? 1'b0 : n5152;
/* FF  5 11  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n733 <= 1'b0; else if (n128) n733 <= n5153;
/* FF 16 18  3 */ assign n5154 = n5155;
/* FF  4  7  6 */ assign n544 = n5156;
/* FF 13 22  0 */ assign n1841 = n5157;
/* FF 14 10  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1936 <= 1'b0; else if (n734) n1936 <= n5158;
/* FF 14  2  2 */ assign n1863 = n5159;
/* FF  1 17  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n122 <= 1'b0; else if (n118) n122 <= n5160;
/* FF 17  9  2 */ assign n2358 = n5161;
/* FF  8  2  5 */ assign n945 = n5162;
/* FF  1 20  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n149 <= 1'b1; else if (n147) n149 <= n5163;
/* FF  7  3  1 */ assign n837 = n5164;
/* FF 10 11  2 */ always @(posedge io_13_31_1) if (n4) n1312 <= 1'b0 ? 1'b0 : n5165;
/* FF  9 15  5 */ always @(posedge io_13_31_1) if (n4) n1194 <= 1'b0 ? 1'b0 : n5166;
/* FF 13 18  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1812 <= 1'b0; else if (n1967) n1812 <= n5167;
/* FF  3 21  1 */ assign n335 = n5168;
/* FF  8  3  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n954 <= 1'b0; else if (n840) n954 <= n5169;
/* FF  1 13  4 */ assign n97 = n5170;
/* FF 17  1  3 */ assign n2305 = n5171;
/* FF 20  9  4 */ always @(posedge io_13_31_1) if (n2093) n2483 <= 1'b0 ? 1'b0 : n5172;
/* FF 18 14  2 */ always @(posedge io_13_31_1) if (n2137) n2543 <= n3 ? 1'b0 : n5173;
/* FF  9  7  0 */ assign n1123 = n5174;
/* FF  7  7  7 */ assign n860 = n5175;
/* FF 21 21  2 */ assign n2872 = n5176;
/* FF 16  6  6 */ assign n2188 = n5177;
/* FF  3 13  2 */ assign n5178 = n5179;
/* FF 10 12  2 */ assign n1322 = n5180;
/* FF  1  5  5 */ always @(posedge io_13_31_1) if (n201) n38 <= n42 ? 1'b0 : n5181;
/* FF 15 19  0 */ assign n2144 = n5182;
/* FF  3 16  7 */ assign n449 = n5183;
/* FF 21 22  3 */ always @(posedge io_13_31_1) if (n2881) n2880 <= 1'b0 ? 1'b0 : n5184;
/* FF 22 18  0 */ assign n2862 = n5185;
/* FF 12 15  6 */ always @(posedge io_13_31_1) if (n1180) n1631 <= n1 ? 1'b0 : n5186;
/* FF 12  7  2 */ assign n1569 = n5187;
/* FF 13  3  0 */ assign n1671 = n5188;
/* FF  4 21  3 */ assign n646 = n5189;
/* FF 18 15  2 */ always @(posedge io_13_31_1) if (n2402) n2550 <= 1'b0 ? 1'b0 : n5190;
/* FF 22 13  7 */ assign n2961 = n5191;
/* FF  3  9  4 */ assign n417 = n5192;
/* FF 11 19  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1514 <= 1'b0; else if (1'b1) n1514 <= n5193;
/* FF  2 10  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n244 <= 1'b1; else if (1'b1) n244 <= n5194;
/* FF  5 18  1 */ assign n774 = n5195;
/* FF  9  3  7 */ assign n1097 = n5196;
/* FF 21  6  0 */ always @(posedge io_13_31_1) if (n2686) n2197 <= 1'b0 ? 1'b0 : n5197;
/* FF 18  2  5 */ always @(posedge io_13_31_1) if (n2456) n2446 <= 1'b0 ? 1'b0 : n5198;
/* FF 13  7  6 */ assign n1724 = n5199;
/* FF  3  2  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n347 <= 1'b0; else if (n500) n347 <= n5200;
/* FF 11 12  4 */ assign n1471 = n5201;
/* FF 12  8  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1579 <= 1'b0; else if (n1430) n1579 <= n5202;
/* FF 11  4  0 */ assign n851 = n5203;
/* FF 15 16  3 */ assign n2135 = n5204;
/* FF  3  1  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n343 <= 1'b0; else if (n500) n343 <= n5205;
/* FF 22 14  7 */ assign n2970 = n5206;
/* FF 15 15  7 */ always @(posedge io_13_31_1) if (n1180) n2132 <= n1 ? 1'b1 : n5207;
/* FF  5 10  2 */ always @(posedge io_13_31_1) if (n4) n725 <= 1'b0 ? 1'b0 : n5208;
/* FF  7 21  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n151 <= 1'b0; else if (1'b1) n151 <= n5209;
/* FF 11  5  1 */ assign n975 = n5210;
/* FF  8 17  2 */ assign n5211 = n5212;
/* FF  5 13  7 */ assign n748 = n5213;
/* FF 23 19  3 */ always @(posedge io_13_31_1) if (n2993) n3040 <= 1'b0 ? 1'b0 : n5214;
/* FF  4  9  6 */ always @(posedge io_13_31_1) if (n4) n562 <= 1'b0 ? 1'b0 : n5215;
/* FF 15  8  4 */ always @(posedge io_13_31_1) if (n1591) n2072 <= 1'b0 ? 1'b0 : n5216;
/* FF 17 19  6 */ assign n2422 = n5217;
/* FF 17 11  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2341 <= 1'b0; else if (n1764) n2341 <= n5218;
/* FF  4  6  0 */ assign n533 = n5219;
/* FF  7 14  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n903 <= 1'b0; else if (1'b1) n903 <= n5220;
/* FF  2  6  7 */ assign n211 = n5221;
/* FF 16 20  2 */ assign n1838 = n5222;
/* FF 14 12  5 */ assign n1946 = n5223;
/* FF 14  4  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1876 <= 1'b0; else if (n1869) n1876 <= n5224;
/* FF 17 20  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2293 <= 1'b0; else if (n2023) n2293 <= n5225;
/* FF 17 12  3 */ always @(posedge io_13_31_1) if (n2137) n2381 <= n3 ? 1'b0 : n5226;
/* FF 23  3  0 */ assign n3012 = n5227;
/* FF 15  4  6 */ assign n1738 = n5228;
/* FF  5  6  3 */ always @(posedge io_13_31_1) if (n4) n688 <= 1'b0 ? 1'b0 : n5229;
/* FF 14 13  6 */ assign n1954 = n5230;
/* FF  4  2  2 */ assign n503 = n5231;
/* FF 14  5  2 */ assign n980 = n5232;
/* FF 16 16  4 */ assign n1823 = n5233;
/* FF 13 21  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1833 <= 1'b0; else if (n1830) n1833 <= n5234;
/* FF  8  5  5 */ assign n198 = n5235;
/* FF 24  3  4 */ always @(posedge io_13_31_1) if (n2902) n2901 <= n7 ? 1'b0 : n5236;
/* FF 10 14  2 */ assign n1343 = n5237;
/* FF  9 18  5 */ assign n5238 = n5239;
/* FF  9 10  1 */ always @(posedge io_13_31_1) if (n4) n1152 <= 1'b0 ? 1'b0 : n5240;
/* FF 16  9  1 */ assign n2215 = n5241;
/* FF  7  2  4 */ assign n805 = n5242;
/* FF  8  6  6 */ assign n679 = n5243;
/* FF 16  8  5 */ assign n2210 = n5244;
/* FF 10 15  3 */ assign n1354 = n5245;
/* FF 20  4  0 */ always @(posedge io_13_31_1) if (n2602) n2481 <= n1 ? 1'b0 : n5246;
/* FF 18 17  2 */ assign n2558 = n5247;
/* FF 13 22  3 */ assign n1844 = n5248;
/* FF  2 21  0 */ assign n5249 = n5250;
/* FF  9 14  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1186 <= 1'b0; else if (n762) n1186 <= n5252;
/* FF 20  5  1 */ assign n5253 = n5254;
/* FF 16  4  7 */ always @(posedge io_13_31_1) if (n2324) n2177 <= 1'b0 ? 1'b0 : n5255;
/* FF  1  8  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n56 <= 1'b0; else if (1'b1) n56 <= n5256;
/* FF  9 11  1 */ always @(posedge io_13_31_1) if (n4) n1159 <= 1'b0 ? 1'b0 : n5257;
/* FF  7  3  4 */ assign n671 = n5258;
/* FF 12 18  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1517 <= 1'b0; else if (1'b1) n1517 <= n5259;
/* FF  2 13  1 */ assign n273 = n5260;
/* FF 13  6  0 */ assign n1707 = n5261;
/* FF  2 16  6 */ assign n129 = n5262;
/* FF 13  9  5 */ assign n1746 = n5263;
/* FF  3 12  4 */ assign n427 = n5264;
/* FF  1  4  7 */ always @(posedge io_13_31_1) if (n201) n34 <= n42 ? 1'b0 : n5265;
/* FF 15 18  2 */ assign n2139 = n5266;
/* FF  4 17  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n456 <= 1'b0; else if (n317) n456 <= n5267;
/* FF  2 17  7 */ assign n302 = n5268;
/* FF 13 10  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1749 <= 1'b0; else if (n734) n1749 <= n5269;
/* FF 13  2  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1668 <= 1'b0; else if (n1670) n1668 <= n5270;
/* FF  2  9  3 */ assign n234 = n5271;
/* FF  3 13  5 */ assign n5272 = n5273;
/* FF  3  5  1 */ assign n374 = n5274;
/* FF 11 15  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1491 <= 1'b0; else if (1'b1) n1491 <= n5275;
/* FF 14 23  5 */ assign n2035 = n5276;
/* FF 11  7  0 */ always @(posedge io_13_31_1) if (n4) n1145 <= 1'b0 ? 1'b0 : n5277;
/* FF 15 19  3 */ assign n5278 = n5279;
/* FF 10  3  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1255 <= 1'b0; else if (n851) n1255 <= n5280;
/* FF 18  6  6 */ always @(posedge io_13_31_1) if (n2602) n2470 <= n1 ? 1'b0 : n5281;
/* FF 12  7  5 */ assign n1572 = n5282;
/* FF 22  9  3 */ always @(posedge io_13_31_1) if (n2686) n2950 <= 1'b0 ? 1'b0 : n5283;
/* FF 21 13  6 */ always @(posedge io_13_31_1) if (n2819) n2824 <= n2823 ? 1'b0 : n5284;
/* FF  4 21  6 */ assign n643 = n5285;
/* FF 21  5  2 */ always @(posedge io_13_31_1) if (n2902) n2778 <= n7 ? 1'b0 : n5286;
/* FF  8 16  5 */ assign n1047 = n5287;
/* FF 15  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2049 <= 1'b0; else if (n1547) n2049 <= n5288;
/* FF 17 22  6 */ assign n2160 = n5289;
/* FF 22  2  0 */ assign n2886 = n5290;
/* FF  7 17  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n465 <= 1'b1; else if (n916) n465 <= n5291;
/* FF 15  6  5 */ always @(posedge io_13_31_1) if (n2191) n1541 <= 1'b0 ? 1'b0 : n5292;
/* FF  5  9  4 */ assign n718 = n5293;
/* FF  4 13  7 */ assign n259 = n5294;
/* FF  4  5  3 */ assign n529 = n5295;
/* FF 16 19  5 */ assign n2287 = n5296;
/* FF 17 15  3 */ assign n2137 = n5297;
/* FF 11  3  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1407 <= 1'b0; else if (n979) n1407 <= n5298;
/* FF  7 18  2 */ assign n5299 = n5300;
/* FF 15  7  6 */ assign n2063 = n5301;
/* FF  9 21  0 */ assign n1221 = n5302;
/* FF  7 21  7 */ assign n929 = n5303;
/* FF 14  8  2 */ assign n1919 = n5304;
/* FF  8  9  1 */ assign n996 = n5305;
/* FF 20 23  3 */ assign n2754 = n5306;
/* FF 17  8  0 */ always @(posedge io_13_31_1) if (n2344) n2347 <= 1'b0 ? 1'b0 : n5307;
/* FF  5  2  0 */ assign n660 = n5308;
/* FF 23  2  2 */ always @(posedge io_13_31_1) if (1'b1) n3005 <= n2888 ? 1'b0 : n5309;
/* FF  4  6  3 */ assign n536 = n5310;
/* FF 17 11  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2377 <= 1'b0; else if (n1764) n2377 <= n5311;
/* FF  9 13  1 */ always @(posedge io_13_31_1) if (n4) n1173 <= 1'b0 ? 1'b0 : n5312;
/* FF 16 12  1 */ always @(posedge io_13_31_1) if (n2120) n2240 <= 1'b0 ? 1'b0 : n5313;
/* FF 13 17  0 */ assign n5314 = n5315;
/* FF  7  5  4 */ always @(posedge io_13_31_1) if (n4) n700 <= 1'b0 ? 1'b0 : n5317;
/* FF 14  4  4 */ assign n1880 = n5318;
/* FF  8  1  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n935 <= 1'b0; else if (n656) n935 <= n5319;
/* FF  1 19  4 */ assign n138 = n5320;
/* FF 23  3  3 */ assign n5321 = n5322;
/* FF  1 11  0 */ assign n76 = n5323;
/* FF  8  4  7 */ assign n957 = n5324;
/* FF 20  7  0 */ assign n5325 = n5326;
/* FF 12 21  1 */ assign n1655 = n5328;
/* FF 17  3  6 */ always @(posedge io_13_31_1) if (n2324) n2322 <= 1'b0 ? 1'b0 : n5329;
/* FF  7  6  5 */ assign n564 = n5330;
/* FF 10 13  4 */ always @(posedge io_13_31_1) if (n4) n1337 <= 1'b0 ? 1'b0 : n5331;
/* FF  9 17  7 */ assign n820 = n5332;
/* FF  9  9  3 */ always @(posedge io_13_31_1) if (n4) n1139 <= 1'b0 ? 1'b0 : n5333;
/* FF 13 21  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1834 <= 1'b0; else if (n1830) n1834 <= n5334;
/* FF  1 12  1 */ assign n83 = n5335;
/* FF 20  8  1 */ assign n5336 = n5337;
/* FF 12 22  2 */ assign n1660 = n5338;
/* FF 20 11  6 */ always @(posedge io_13_31_1) if (n2137) n2701 <= n3 ? 1'b0 : n5339;
/* FF 10 14  5 */ assign n1346 = n5340;
/* FF 10  6  1 */ assign n960 = n5341;
/* FF 18 16  4 */ always @(posedge io_13_31_1) if (n2011) n2554 <= 1'b0 ? 1'b0 : n5342;
/* FF  9 10  4 */ assign n1155 = n5343;
/* FF  9  2  0 */ assign n1084 = n5344;
/* FF 22 20  3 */ assign n2998 = n5345;
/* FF  7  2  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n659 <= 1'b0; else if (n509) n659 <= n5346;
/* FF 21 24  6 */ always @(posedge io_13_31_1) if (n2884) n2885 <= 1'b0 ? 1'b0 : n5347;
/* FF  2 19  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n323 <= 1'b0; else if (n322) n323 <= n5348;
/* FF 13 13  7 */ always @(posedge io_13_31_1) if (1'b1) n1777 <= 1'b0 ? 1'b0 : n5349;
/* FF  3 15  4 */ assign n434 = n5350;
/* FF 20  4  3 */ assign n2671 = n5351;
/* FF  3  7  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n396 <= 1'b0; else if (n224) n396 <= n5352;
/* FF 11 18  5 */ assign n1511 = n5353;
/* FF 18  9  1 */ assign n2492 = n5354;
/* FF  4 20  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n490 <= 1'b0; else if (n629) n490 <= n5355;
/* FF  2 20  7 */ assign n330 = n5356;
/* FF 12  9  4 */ assign n1587 = n5357;
/* FF 22 12  4 */ assign n2720 = n5358;
/* FF  2 12  3 */ assign n250 = n5359;
/* FF 13  5  2 */ assign n1280 = n5360;
/* FF  3  8  1 */ assign n403 = n5361;
/* FF 21  8  3 */ assign n5362 = n5363;
/* FF 14 18  1 */ always @(posedge io_13_31_1) if (n1513) n1993 <= n1 ? 1'b0 : n5364;
/* FF  3 11  6 */ assign n423 = n5365;
/* FF 11 14  7 */ assign n1485 = n5366;
/* FF 18  1  2 */ assign n2440 = n5367;
/* FF  2 13  4 */ assign n272 = n5368;
/* FF 13  6  3 */ assign n1710 = n5369;
/* FF  2  5  0 */ assign n202 = n5370;
/* FF  4 16  2 */ assign n607 = n5371;
/* FF 11 11  1 */ assign n5372 = n5373;
/* FF 14 19  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1982 <= 1'b0; else if (n1527) n1982 <= n5374;
/* FF 22  8  6 */ assign n2686 = n5375;
/* FF 15 15  0 */ assign n5376 = n5377;
/* FF  3  4  3 */ assign n366 = n5379;
/* FF 21  4  5 */ always @(posedge io_13_31_1) if (n2902) n2773 <= n7 ? 1'b0 : n5380;
/* FF 15 18  5 */ assign n5381 = n5382;
/* FF  8 19  5 */ assign n5383 = n5384;
/* FF 22  5  0 */ assign n2925 = n5385;
/* FF  7 20  1 */ assign n5386 = n5387;
/* FF  4  8  3 */ always @(posedge io_13_31_1) if (n4) n550 <= 1'b0 ? 1'b0 : n5388;
/* FF  8 20  6 */ assign n1063 = n5389;
/* FF 11  7  3 */ always @(posedge io_13_31_1) if (n4) n1032 <= 1'b0 ? 1'b0 : n5390;
/* FF 17 18  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2411 <= 1'b0; else if (n2011) n2411 <= n5391;
/* FF 15 10  6 */ always @(posedge io_13_31_1) if (n1591) n2090 <= 1'b0 ? 1'b0 : n5392;
/* FF 15  2  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1882 <= 1'b0; else if (n1552) n1882 <= n5393;
/* FF  5  5  1 */ assign n682 = n5394;
/* FF  4  1  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n492 <= 1'b0; else if (n656) n492 <= n5395;
/* FF 16 15  2 */ always @(posedge io_13_31_1) if (n2268) n2249 <= 1'b0 ? 1'b0 : n5396;
/* FF 15  3  3 */ assign n967 = n5397;
/* FF 23 13  6 */ always @(posedge io_13_31_1) if (n2842) n2962 <= 1'b0 ? 1'b0 : n5398;
/* FF 17 14  5 */ always @(posedge io_13_31_1) if (n2396) n2267 <= n1 ? 1'b0 : n5399;
/* FF  1 14  1 */ assign n106 = n5400;
/* FF  7 17  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n615 <= 1'b0; else if (n916) n615 <= n5401;
/* FF  7  9  0 */ assign n5402 = n5403;
/* FF  2  1  6 */ assign n165 = n5405;
/* FF 13 20  0 */ assign n5406 = n5407;
/* FF 14  7  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1909 <= 1'b0; else if (n1279) n1909 <= n5409;
/* FF 13 23  5 */ assign n1859 = n5410;
/* FF  3 18  0 */ assign n5411 = n5412;
/* FF 17  6  6 */ assign n5414 = n5415;
/* FF 10 16  4 */ always @(posedge io_13_31_1) if (n4) n1350 <= 1'b0 ? 1'b0 : n5416;
/* FF  7  1  1 */ assign n823 = n5417;
/* FF  9 20  7 */ assign n1219 = n5418;
/* FF  9 12  3 */ assign n1168 = n5419;
/* FF  7  4  6 */ assign n846 = n5420;
/* FF  3 19  1 */ assign n467 = n5421;
/* FF 20 14  6 */ always @(posedge io_13_31_1) if (n2137) n2718 <= n3 ? 1'b0 : n5422;
/* FF 10 17  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1360 <= 1'b0; else if (n1502) n1360 <= n5423;
/* FF 20  6  2 */ always @(posedge io_13_31_1) if (n2676) n2678 <= n1 ? 1'b0 : n5424;
/* FF 10  9  1 */ assign n1294 = n5425;
/* FF  9 13  4 */ always @(posedge io_13_31_1) if (n4) n1176 <= 1'b0 ? 1'b0 : n5426;
/* FF  9  5  0 */ assign n1108 = n5427;
/* FF  7  5  7 */ assign n524 = n5428;
/* FF 20  7  3 */ assign n5429 = n5430;
/* FF 13  8  3 */ assign n1734 = n5431;
/* FF 18 12  1 */ assign n2522 = n5432;
/* FF  3 14  7 */ assign n285 = n5433;
/* FF 10  1  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1236 <= 1'b0; else if (n1120) n1236 <= n5434;
/* FF 22 15  4 */ always @(posedge io_13_31_1) if (1'b1) n2974 <= n3025 ? 1'b0 : n5435;
/* FF  2 15  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n288 <= 1'b0; else if (1'b1) n288 <= n5436;
/* FF 10  4  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1262 <= 1'b0; else if (n979) n1262 <= n5437;
/* FF 21 11  3 */ always @(posedge io_13_31_1) if (n2213) n2629 <= 1'b0 ? 1'b0 : n5438;
/* FF 14 21  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2019 <= 1'b0; else if (1'b1) n2019 <= n5439;
/* FF  1  3  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n22 <= 1'b0; else if (n17) n22 <= n5440;
/* FF 13  4  5 */ assign n1685 = n5441;
/* FF 11 17  7 */ assign n1507 = n5442;
/* FF 11  9  3 */ assign n1445 = n5443;
/* FF 12 13  5 */ always @(posedge io_13_31_1) if (n4) n1613 <= 1'b0 ? 1'b0 : n5444;
/* FF 12  5  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1281 <= 1'b0; else if (n1426) n1281 <= n5445;
/* FF  2  8  0 */ assign n5446 = n5447;
/* FF  4 19  2 */ assign n625 = n5449;
/* FF  9  1  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1082 <= 1'b0; else if (n851) n1082 <= n5450;
/* FF  2 11  5 */ assign n255 = n5451;
/* FF 21  7  5 */ assign n5452 = n5453;
/* FF 11 10  4 */ assign n1459 = n5454;
/* FF 15 21  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2155 <= 1'b1; else if (n1526) n2155 <= n5455;
/* FF 12  6  2 */ assign n1558 = n5456;
/* FF 15 13  1 */ assign n2115 = n5457;
/* FF  5 16  0 */ assign n598 = n5458;
/* FF 12  9  7 */ assign n1590 = n5459;
/* FF 22 12  7 */ assign n2395 = n5460;
/* FF 22  4  3 */ assign n2902 = n5461;
/* FF  2  4  2 */ assign n190 = n5462;
/* FF 21  8  6 */ always @(posedge io_13_31_1) if (n2694) n2803 <= n1 ? 1'b0 : n5463;
/* FF  4 11  3 */ assign n104 = n5464;
/* FF  8 15  2 */ assign n5465 = n5466;
/* FF  2  3  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n186 <= 1'b0; else if (n17) n186 <= n5467;
/* FF  8 18  7 */ assign n1057 = n5468;
/* FF 18  1  5 */ assign n2313 = n5469;
/* FF 15  5  2 */ assign n2054 = n5470;
/* FF  5  8  1 */ always @(posedge io_13_31_1) if (n4) n703 <= 1'b0 ? 1'b0 : n5471;
/* FF  4  4  0 */ assign n519 = n5472;
/* FF 16 18  2 */ assign n1999 = n5473;
/* FF  4  7  5 */ assign n546 = n5474;
/* FF 14 10  5 */ assign n1935 = n5475;
/* FF  8 11  4 */ assign n1016 = n5476;
/* FF 14  2  1 */ assign n1549 = n5477;
/* FF 16 21  7 */ assign n2038 = n5478;
/* FF 23  8  2 */ always @(posedge io_13_31_1) if (1'b1) n3014 <= 1'b0 ? 1'b0 : n5479;
/* FF  7 20  4 */ assign n5480 = n5481;
/* FF 17  9  1 */ always @(posedge io_13_31_1) if (n1591) n2357 <= 1'b0 ? 1'b0 : n5482;
/* FF  5 12  7 */ assign n575 = n5483;
/* FF  5  4  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n41 <= 1'b0; else if (n217) n41 <= n5484;
/* FF  4  8  6 */ assign n553 = n5485;
/* FF 16 14  4 */ assign n2245 = n5486;
/* FF 17 10  2 */ assign n2366 = n5487;
/* FF 14  6  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1901 <= 1'b0; else if (n1279) n1901 <= n5488;
/* FF  3 21  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n482 <= 1'b0; else if (1'b1) n482 <= n5489;
/* FF  8  3  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n953 <= 1'b0; else if (n840) n953 <= n5490;
/* FF  1 21  7 */ assign n157 = n5491;
/* FF 15  2  5 */ assign n2046 = n5492;
/* FF 18 23  1 */ always @(posedge io_13_31_1) if (n2594) n2592 <= 1'b0 ? 1'b0 : n5493;
/* FF  1 13  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n96 <= 1'b0; else if (n105) n96 <= n5494;
/* FF 20 17  7 */ assign n2566 = n5495;
/* FF 14  3  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1704 <= 1'b0; else if (n1690) n1704 <= n5496;
/* FF 12 23  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1528 <= 1'b0; else if (n1666) n1528 <= n5497;
/* FF 13 19  2 */ assign n1817 = n5498;
/* FF  7  7  6 */ assign n859 = n5499;
/* FF  1 14  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n108 <= 1'b0; else if (1'b1) n108 <= n5500;
/* FF 16  6  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1692 <= 1'b0; else if (n1433) n1692 <= n5501;
/* FF  1  6  0 */ assign n5502 = n5503;
/* FF 10 20  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1380 <= 1'b0; else if (n1390) n1380 <= n5505;
/* FF 10 12  1 */ always @(posedge io_13_31_1) if (n1180) n1321 <= n1 ? 1'b0 : n5506;
/* FF  9  8  0 */ assign n1128 = n5507;
/* FF 13 20  3 */ assign n1827 = n5508;
/* FF  7  8  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n871 <= 1'b0; else if (1'b1) n871 <= n5509;
/* FF 18 18  7 */ assign n2565 = n5510;
/* FF 20 10  3 */ always @(posedge io_13_31_1) if (n2112) n2371 <= 1'b0 ? 1'b0 : n5511;
/* FF 16  2  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2169 <= 1'b0; else if (n1552) n2169 <= n5512;
/* FF 12 16  0 */ always @(posedge io_13_31_1) if (n4) n1633 <= 1'b0 ? 1'b0 : n5513;
/* FF  3 17  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n142 <= 1'b0; else if (1'b1) n142 <= n5514;
/* FF 10 16  7 */ always @(posedge io_13_31_1) if (n4) n1365 <= 1'b0 ? 1'b0 : n5515;
/* FF 22 19  0 */ assign n2868 = n5516;
/* FF  9 12  6 */ assign n1031 = n5517;
/* FF  5 18  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n642 <= 1'b0; else if (n474) n642 <= n5518;
/* FF 11 21  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n426 <= 1'b0; else if (1'b1) n426 <= n5519;
/* FF 12 11  7 */ assign n1600 = n5520;
/* FF 13  7  5 */ assign n1723 = n5521;
/* FF  3 10  4 */ assign n69 = n5522;
/* FF  3  2  0 */ assign n346 = n5523;
/* FF 18 11  3 */ assign n2515 = n5524;
/* FF  1  2  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n14 <= 1'b0; else if (n17) n14 <= n5525;
/* FF 12  8  1 */ assign n1578 = n5526;
/* FF 15 16  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2128 <= 1'b0; else if (n1811) n2128 <= n5527;
/* FF  9  4  7 */ assign n1100 = n5528;
/* FF 22 14  6 */ always @(posedge io_13_31_1) if (1'b1) n2969 <= n3025 ? 1'b0 : n5529;
/* FF  2 14  5 */ assign n283 = n5530;
/* FF 13  8  6 */ assign n1737 = n5531;
/* FF 21 10  5 */ always @(posedge io_13_31_1) if (n2137) n2808 <= n3 ? 1'b0 : n5532;
/* FF 21  2  1 */ always @(posedge io_13_31_1) if (1'b1) n7 <= n2761 ? 1'b0 : n5533;
/* FF 11 13  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n422 <= 1'b0; else if (n1461) n422 <= n5534;
/* FF 11  5  0 */ assign n979 = n5535;
/* FF  5 19  0 */ assign n782 = n5536;
/* FF 10  1  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1239 <= 1'b0; else if (n1120) n1239 <= n5537;
/* FF 12 12  7 */ assign n817 = n5538;
/* FF 22 15  7 */ assign n2977 = n5539;
/* FF  2 15  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n290 <= 1'b0; else if (1'b1) n290 <= n5540;
/* FF 12  4  3 */ assign n1544 = n5541;
/* FF 22  7  3 */ always @(posedge io_13_31_1) if (n2694) n2691 <= n1 ? 1'b0 : n5542;
/* FF  2  7  2 */ assign n219 = n5543;
/* FF 21 11  6 */ always @(posedge io_13_31_1) if (n2213) n2639 <= 1'b0 ? 1'b0 : n5544;
/* FF 21  3  2 */ always @(posedge io_13_31_1) if (n2902) n2762 <= n7 ? 1'b0 : n5545;
/* FF 11  6  1 */ assign n1106 = n5546;
/* FF  5 14  7 */ assign n756 = n5547;
/* FF  8 21  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1050 <= 1'b0; else if (n1068) n1050 <= n5548;
/* FF 17 20  6 */ assign n2298 = n5549;
/* FF 15  4  5 */ assign n2051 = n5550;
/* FF  5  6  2 */ assign n687 = n5551;
/* FF  4 10  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n64 <= 1'b0; else if (n576) n64 <= n5552;
/* FF 14 13  5 */ assign n1953 = n5553;
/* FF  4  2  1 */ assign n502 = n5554;
/* FF  8 14  4 */ assign n1039 = n5555;
/* FF 14  5  1 */ assign n1886 = n5556;
/* FF 16 24  7 */ always @(posedge io_13_31_1) if (n2301) n2302 <= 1'b0 ? 1'b0 : n5557;
/* FF 16 16  3 */ assign n2273 = n5558;
/* FF 11  1  7 */ assign n5559 = n5560;
/* FF  7 15  0 */ assign n5561 = n5562;
/* FF  5 15  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n761 <= 1'b0; else if (n451) n761 <= n5564;
/* FF  5  7  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n410 <= 1'b0; else if (n532) n410 <= n5565;
/* FF  9 19  0 */ assign n5566 = n5567;
/* FF  4 11  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n62 <= 1'b0; else if (1'b1) n62 <= n5568;
/* FF  4  3  2 */ assign n512 = n5569;
/* FF  8  7  1 */ assign n5570 = n5571;
/* FF 16  9  0 */ assign n2214 = n5572;
/* FF 20 21  3 */ assign n2749 = n5573;
/* FF 14  9  7 */ always @(posedge io_13_31_1) if (n1739) n1596 <= 1'b0 ? 1'b0 : n5574;
/* FF 17 13  2 */ always @(posedge io_13_31_1) if (n2536) n2385 <= n1 ? 1'b0 : n5575;
/* FF  8  6  5 */ assign n509 = n5576;
/* FF 15  5  5 */ assign n1115 = n5577;
/* FF 20 20  7 */ assign n2746 = n5578;
/* FF  7 11  2 */ always @(posedge io_13_31_1) if (n4) n883 <= 1'b0 ? 1'b0 : n5579;
/* FF 10 15  2 */ always @(posedge io_13_31_1) if (n4) n1351 <= 1'b0 ? 1'b0 : n5580;
/* FF 16 10  1 */ assign n2222 = n5581;
/* FF 13 22  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1843 <= 1'b0; else if (n1666) n1843 <= n5582;
/* FF 10 18  7 */ assign n5583 = n5584;
/* FF 14  2  4 */ assign n1865 = n5585;
/* FF  1 17  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n123 <= 1'b0; else if (n118) n123 <= n5586;
/* FF  1  9  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n53 <= 1'b0; else if (n70) n53 <= n5587;
/* FF  8  2  7 */ assign n946 = n5588;
/* FF 20  5  0 */ assign n5589 = n5590;
/* FF 12 19  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1553 <= 1'b0; else if (n1815) n1553 <= n5592;
/* FF  7  3  3 */ assign n178 = n5593;
/* FF 10 11  4 */ assign n1314 = n5594;
/* FF 18 21  7 */ always @(posedge io_13_31_1) if (n2584) n2585 <= 1'b0 ? 1'b0 : n5595;
/* FF  9 15  7 */ assign n1196 = n5596;
/* FF  1 10  1 */ assign n73 = n5597;
/* FF 13 18  4 */ assign n1813 = n5598;
/* FF  3 21  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n483 <= 1'b1; else if (1'b1) n483 <= n5599;
/* FF  1 13  6 */ assign n99 = n5600;
/* FF 16  5  7 */ assign n2181 = n5601;
/* FF 17  1  5 */ always @(posedge io_13_31_1) if (1'b1) n189 <= 1'b0 ? 1'b0 : n5602;
/* FF 20  9  6 */ always @(posedge io_13_31_1) if (n2093) n2624 <= 1'b0 ? 1'b0 : n5603;
/* FF 18 14  4 */ always @(posedge io_13_31_1) if (n2137) n2544 <= n3 ? 1'b0 : n5604;
/* FF  9  7  2 */ assign n811 = n5605;
/* FF 13 11  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1750 <= 1'b0; else if (n734) n1750 <= n5606;
/* FF 21 21  4 */ assign n2874 = n5607;
/* FF  2 17  6 */ assign n301 = n5608;
/* FF 13 10  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1732 <= 1'b0; else if (n734) n1732 <= n5609;
/* FF  3 13  4 */ assign n5610 = n5611;
/* FF  3  5  0 */ assign n373 = n5612;
/* FF 10  4  0 */ assign n1250 = n5613;
/* FF  1  5  7 */ always @(posedge io_13_31_1) if (n201) n40 <= n42 ? 1'b0 : n5614;
/* FF 15 19  2 */ assign n2145 = n5615;
/* FF 22 18  2 */ assign n2988 = n5616;
/* FF 10  3  4 */ assign n1254 = n5617;
/* FF 21 14  1 */ assign n2830 = n5618;
/* FF 12  7  4 */ assign n1571 = n5619;
/* FF 13  3  2 */ assign n1673 = n5620;
/* FF 21 13  5 */ assign n2823 = n5621;
/* FF  3  6  1 */ assign n385 = n5622;
/* FF  4 21  5 */ assign n647 = n5623;
/* FF 11  8  0 */ always @(posedge io_13_31_1) if (n4) n1436 <= 1'b0 ? 1'b0 : n5624;
/* FF 15 20  3 */ assign n2153 = n5625;
/* FF  3  9  6 */ assign n116 = n5626;
/* FF 17 23  1 */ always @(posedge io_13_31_1) if (n2437) n2436 <= 1'b0 ? 1'b0 : n5627;
/* FF 22 10  3 */ assign n2113 = n5628;
/* FF  2 10  2 */ assign n245 = n5629;
/* FF  5 18  3 */ assign n775 = n5630;
/* FF 21  6  2 */ always @(posedge io_13_31_1) if (n2686) n2195 <= 1'b0 ? 1'b0 : n5631;
/* FF 18  2  7 */ assign n2182 = n5632;
/* FF 21  9  7 */ always @(posedge io_13_31_1) if (1'b1) n188 <= 1'b0 ? 1'b0 : n5633;
/* FF 17 24  2 */ always @(posedge io_13_31_1) if (n2438) n2435 <= 1'b0 ? 1'b0 : n5634;
/* FF 11 12  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1474 <= 1'b0; else if (n102) n1474 <= n5635;
/* FF 12  8  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1575 <= 1'b0; else if (n1430) n1575 <= n5636;
/* FF 11  4  2 */ assign n1410 = n5637;
/* FF  3  1  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n345 <= 1'b0; else if (n500) n345 <= n5638;
/* FF 22  3  0 */ assign n2895 = n5639;
/* FF  4 14  1 */ assign n591 = n5640;
/* FF  7 18  1 */ assign n5641 = n5642;
/* FF 22  6  5 */ assign n2456 = n5643;
/* FF  5 10  4 */ always @(posedge io_13_31_1) if (n4) n727 <= 1'b0 ? 1'b0 : n5644;
/* FF 21  2  4 */ assign n2600 = n5645;
/* FF  7 21  6 */ assign n928 = n5646;
/* FF  8 17  4 */ assign n5647 = n5648;
/* FF  8  9  0 */ assign n5649 = n5650;
/* FF 18  3  7 */ always @(posedge io_13_31_1) if (n2191) n2178 <= 1'b0 ? 1'b0 : n5652;
/* FF 15  8  6 */ assign n2074 = n5653;
/* FF  9 22  0 */ assign n5654 = n5655;
/* FF  4  6  2 */ assign n538 = n5657;
/* FF  8 10  1 */ always @(posedge io_13_31_1) if (n4) n1007 <= 1'b0 ? 1'b0 : n5658;
/* FF 16 20  4 */ always @(posedge io_13_31_1) if (n2024) n2290 <= 1'b0 ? 1'b0 : n5659;
/* FF 16 12  0 */ assign n2238 = n5660;
/* FF 14 12  7 */ assign n1948 = n5661;
/* FF 14  4  3 */ assign n1879 = n5662;
/* FF  5  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n665 <= 1'b0; else if (n198) n665 <= n5663;
/* FF 23  3  2 */ assign n3013 = n5664;
/* FF 17 12  5 */ assign n2383 = n5665;
/* FF 17  4  1 */ always @(posedge io_13_31_1) if (n2316) n2326 <= 1'b0 ? 1'b0 : n5666;
/* FF  5  6  5 */ always @(posedge io_13_31_1) if (n4) n689 <= 1'b0 ? 1'b0 : n5667;
/* FF 16 13  1 */ assign n2247 = n5668;
/* FF  4  2  4 */ assign n505 = n5669;
/* FF  7  6  4 */ always @(posedge io_13_31_1) if (n4) n574 <= 1'b0 ? 1'b0 : n5670;
/* FF 14  5  4 */ assign n1443 = n5671;
/* FF 16 16  6 */ always @(posedge io_13_31_1) if (1'b1) n2274 <= 1'b0 ? 1'b0 : n5672;
/* FF  1 12  0 */ assign n82 = n5673;
/* FF  8  5  7 */ assign n971 = n5674;
/* FF 20  8  0 */ assign n2687 = n5675;
/* FF 12 22  1 */ assign n1659 = n5676;
/* FF 20 11  5 */ assign n2700 = n5677;
/* FF 10 14  4 */ always @(posedge io_13_31_1) if (n4) n1345 <= 1'b0 ? 1'b0 : n5678;
/* FF  9 18  7 */ assign n5679 = n5680;
/* FF  9 10  3 */ always @(posedge io_13_31_1) if (n4) n1154 <= 1'b0 ? 1'b0 : n5681;
/* FF 22 20  2 */ assign n2997 = n5682;
/* FF  7  2  6 */ assign n833 = n5683;
/* FF 21 16  1 */ assign n2844 = n5684;
/* FF 16  8  7 */ always @(posedge io_13_31_1) if (n2344) n2212 <= 1'b0 ? 1'b0 : n5685;
/* FF 20 12  6 */ assign n2705 = n5686;
/* FF 10 15  5 */ always @(posedge io_13_31_1) if (n4) n1340 <= 1'b0 ? 1'b0 : n5687;
/* FF 10  7  1 */ always @(posedge io_13_31_1) if (n4) n1273 <= 1'b0 ? 1'b0 : n5688;
/* FF 18  9  0 */ assign n2379 = n5689;
/* FF 22 21  3 */ always @(posedge io_13_31_1) if (n2882) n3000 <= 1'b0 ? 1'b0 : n5690;
/* FF  2 21  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n325 <= 1'b0; else if (n160) n325 <= n5691;
/* FF 20  5  3 */ always @(posedge io_13_31_1) if (n2472) n2674 <= n2471 ? 1'b0 : n5692;
/* FF  3  8  0 */ assign n5693 = n5694;
/* FF  1  8  7 */ assign n58 = n5696;
/* FF 18 10  1 */ assign n2504 = n5697;
/* FF 12 11  0 */ assign n1566 = n5698;
/* FF 21 17  1 */ assign n2735 = n5699;
/* FF 12 10  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1291 <= 1'b0; else if (n1430) n1291 <= n5700;
/* FF 13  6  2 */ assign n1709 = n5701;
/* FF 10  2  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1248 <= 1'b0; else if (n979) n1248 <= n5702;
/* FF 11 11  0 */ assign n5703 = n5704;
/* FF 13  9  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1741 <= 1'b0; else if (n734) n1741 <= n5706;
/* FF 14 19  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1956 <= 1'b0; else if (n1527) n1956 <= n5707;
/* FF  3 12  6 */ assign n429 = n5708;
/* FF  3  4  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n365 <= 1'b0; else if (n524) n365 <= n5709;
/* FF 15 18  4 */ assign n2140 = n5710;
/* FF 12  3  1 */ assign n5711 = n5712;
/* FF 24 17  3 */ always @(posedge io_13_31_1) if (n2736) n3054 <= 1'b0 ? 1'b0 : n5713;
/* FF  4 17  2 */ assign n613 = n5714;
/* FF 18  5  7 */ always @(posedge io_13_31_1) if (n2456) n2464 <= 1'b0 ? 1'b0 : n5715;
/* FF  2  9  5 */ assign n241 = n5716;
/* FF 13  2  4 */ assign n1670 = n5717;
/* FF  3  5  3 */ assign n376 = n5718;
/* FF 11 15  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1464 <= 1'b0; else if (1'b1) n1464 <= n5719;
/* FF 16 23  0 */ assign n2157 = n5720;
/* FF 11  7  2 */ always @(posedge io_13_31_1) if (n4) n893 <= 1'b0 ? 1'b0 : n5721;
/* FF  8 20  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1044 <= 1'b0; else if (n1062) n1044 <= n5722;
/* FF 15 19  5 */ always @(posedge io_13_31_1) if (n2287) n2010 <= 1'b0 ? 1'b0 : n5723;
/* FF 15 11  1 */ assign n2095 = n5724;
/* FF 10  3  7 */ assign n972 = n5725;
/* FF 23 21  4 */ always @(posedge io_13_31_1) if (n2751) n3041 <= 1'b0 ? 1'b0 : n5726;
/* FF  5 14  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n752 <= 1'b0; else if (1'b1) n752 <= n5727;
/* FF 12  7  7 */ assign n1444 = n5728;
/* FF 21  5  4 */ always @(posedge io_13_31_1) if (n2902) n2780 <= n7 ? 1'b0 : n5729;
/* FF 11  8  3 */ always @(posedge io_13_31_1) if (n4) n1438 <= 1'b0 ? 1'b0 : n5730;
/* FF 23 14  1 */ assign n3020 = n5731;
/* FF  8 16  7 */ assign n919 = n5732;
/* FF 15  3  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1890 <= 1'b0; else if (n1547) n1890 <= n5733;
/* FF 22  2  2 */ assign n2888 = n5734;
/* FF 17 14  4 */ always @(posedge io_13_31_1) if (n2396) n2265 <= n1 ? 1'b0 : n5735;
/* FF  7 17  3 */ assign n915 = n5736;
/* FF 15  6  7 */ assign n2058 = n5737;
/* FF  8 13  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n910 <= 1'b0; else if (n1166) n910 <= n5738;
/* FF  2  1  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n164 <= 1'b0; else if (n178) n164 <= n5739;
/* FF  5  9  6 */ assign n720 = n5740;
/* FF  4  5  5 */ assign n530 = n5741;
/* FF 14  7  3 */ assign n1908 = n5742;
/* FF 16 19  7 */ always @(posedge io_13_31_1) if (n1513) n1987 <= n1 ? 1'b0 : n5743;
/* FF 23  6  2 */ always @(posedge io_13_31_1) if (1'b1) n2693 <= n2916 ? 1'b0 : n5744;
/* FF 17  7  1 */ assign n2342 = n5745;
/* FF  7 18  4 */ assign n5746 = n5747;
/* FF  5 10  7 */ assign n728 = n5748;
/* FF  9 21  2 */ assign n1222 = n5749;
/* FF 20 20  0 */ assign n2740 = n5750;
/* FF 14  8  4 */ assign n1921 = n5751;
/* FF  8  9  3 */ assign n998 = n5752;
/* FF 13 16  1 */ assign n1803 = n5753;
/* FF  8  8  7 */ assign n986 = n5754;
/* FF  3 19  0 */ assign n5755 = n5756;
/* FF  5  2  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n657 <= 1'b0; else if (n509) n657 <= n5758;
/* FF 23  2  4 */ assign n5759 = n5760;
/* FF 10 17  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1370 <= 1'b0; else if (n1502) n1370 <= n5761;
/* FF  9 13  3 */ assign n1175 = n5762;
/* FF 16 12  3 */ assign n2241 = n5763;
/* FF 13 17  2 */ assign n1808 = n5764;
/* FF  7  5  6 */ always @(posedge io_13_31_1) if (n4) n701 <= 1'b0 ? 1'b0 : n5765;
/* FF  8  1  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n937 <= 1'b0; else if (n656) n937 <= n5766;
/* FF  1 19  6 */ assign n140 = n5767;
/* FF  1 11  2 */ assign n77 = n5768;
/* FF 20  7  2 */ assign n2684 = n5769;
/* FF 10 10  1 */ always @(posedge io_13_31_1) if (n4) n1303 <= 1'b0 ? 1'b0 : n5770;
/* FF 12 21  3 */ assign n1657 = n5771;
/* FF  7  6  7 */ always @(posedge io_13_31_1) if (n4) n722 <= 1'b0 ? 1'b0 : n5772;
/* FF 10 13  6 */ always @(posedge io_13_31_1) if (n4) n1338 <= 1'b0 ? 1'b0 : n5773;
/* FF  3 20  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n477 <= 1'b0; else if (n629) n477 <= n5774;
/* FF 21 20  2 */ assign n2863 = n5775;
/* FF  9  9  5 */ assign n1141 = n5776;
/* FF 20  8  3 */ assign n5777 = n5778;
/* FF 21 23  7 */ assign n2884 = n5779;
/* FF 12 22  4 */ assign n1662 = n5780;
/* FF 18 13  1 */ always @(posedge io_13_31_1) if (n2137) n2529 <= n3 ? 1'b0 : n5781;
/* FF 12 14  0 */ assign n5782 = n5783;
/* FF 10  6  3 */ assign n1268 = n5785;
/* FF 18 16  6 */ always @(posedge io_13_31_1) if (n2011) n2556 <= 1'b0 ? 1'b0 : n5786;
/* FF  9  2  2 */ assign n1085 = n5787;
/* FF 21 16  4 */ assign n2846 = n5788;
/* FF  3 15  6 */ assign n435 = n5789;
/* FF  3  7  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n398 <= 1'b0; else if (n224) n398 <= n5790;
/* FF 11 10  3 */ always @(posedge io_13_31_1) if (n4) n1458 <= 1'b0 ? 1'b0 : n5791;
/* FF 18  9  3 */ assign n2494 = n5792;
/* FF 12  6  1 */ assign n1557 = n5793;
/* FF 15 13  0 */ assign n2114 = n5794;
/* FF  4 20  2 */ assign n636 = n5795;
/* FF 12  9  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1589 <= 1'b0; else if (n1164) n1589 <= n5796;
/* FF  2 12  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n101 <= 1'b0; else if (1'b1) n101 <= n5797;
/* FF 13  5  4 */ assign n1695 = n5798;
/* FF 22  4  2 */ assign n2911 = n5799;
/* FF  3  8  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n405 <= 1'b0; else if (n71) n405 <= n5800;
/* FF  2  4  1 */ always @(posedge io_13_31_1) if (n201) n193 <= n42 ? 1'b0 : n5801;
/* FF 21  8  5 */ assign n2802 = n5802;
/* FF 14 18  3 */ always @(posedge io_13_31_1) if (n1513) n1995 <= n1 ? 1'b0 : n5803;
/* FF 15 14  1 */ assign n1180 = n5804;
/* FF  5 17  0 */ assign n768 = n5805;
/* FF 12 10  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1135 <= 1'b0; else if (n1430) n1135 <= n5806;
/* FF 18  1  4 */ assign n2442 = n5807;
/* FF 12  2  3 */ assign n1538 = n5808;
/* FF  2  5  2 */ assign n203 = n5809;
/* FF 24 16  5 */ always @(posedge io_13_31_1) if (n2980) n3053 <= 1'b0 ? 1'b0 : n5810;
/* FF  4 16  4 */ assign n609 = n5811;
/* FF 11 11  3 */ assign n5812 = n5813;
/* FF 14 19  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1984 <= 1'b0; else if (n1527) n1984 <= n5814;
/* FF 14 11  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1452 <= 1'b0; else if (n734) n1452 <= n5815;
/* FF 21  4  7 */ always @(posedge io_13_31_1) if (n2902) n2775 <= n7 ? 1'b0 : n5816;
/* FF  8 19  7 */ assign n5817 = n5818;
/* FF 20 22  0 */ always @(posedge io_13_31_1) if (n2740) n2752 <= 1'b0 ? 1'b0 : n5819;
/* FF  8 11  3 */ always @(posedge io_13_31_1) if (n4) n1015 <= 1'b0 ? 1'b0 : n5820;
/* FF 22  5  2 */ assign n2927 = n5821;
/* FF 21  1  1 */ always @(posedge io_13_31_1) if (n2600) n2314 <= n2757 ? 1'b1 : n5822;
/* FF  7 20  3 */ assign n5823 = n5824;
/* FF 15  9  7 */ assign n2084 = n5825;
/* FF  5 12  6 */ assign n734 = n5826;
/* FF  5  4  2 */ assign n674 = n5827;
/* FF  4  8  5 */ assign n552 = n5828;
/* FF 16 14  3 */ assign n1765 = n5829;
/* FF 17 18  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2413 <= 1'b0; else if (n2011) n2413 <= n5830;
/* FF 17 10  1 */ assign n2355 = n5831;
/* FF 14  6  6 */ assign n1900 = n5832;
/* FF  7 13  0 */ always @(posedge io_13_31_1) if (n4) n894 <= 1'b0 ? 1'b0 : n5833;
/* FF 15  2  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1691 <= 1'b0; else if (n1552) n1691 <= n5834;
/* FF  5  5  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n684 <= 1'b0; else if (n524) n684 <= n5835;
/* FF  4  1  2 */ assign n494 = n5836;
/* FF 14  3  0 */ assign n1870 = n5837;
/* FF 16 15  4 */ always @(posedge io_13_31_1) if (n2268) n2261 <= 1'b0 ? 1'b0 : n5838;
/* FF 16  7  0 */ assign n2198 = n5839;
/* FF 20 18  1 */ assign n2729 = n5840;
/* FF 15  3  5 */ assign n1547 = n5841;
/* FF 17 14  7 */ always @(posedge io_13_31_1) if (n2396) n2394 <= n1 ? 1'b0 : n5842;
/* FF  1 14  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n107 <= 1'b0; else if (1'b1) n107 <= n5843;
/* FF  7  9  2 */ assign n862 = n5844;
/* FF 13 20  2 */ assign n1824 = n5845;
/* FF  7  8  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n870 <= 1'b0; else if (1'b1) n870 <= n5846;
/* FF 14  7  6 */ assign n1911 = n5847;
/* FF 13 23  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1848 <= 1'b0; else if (n1666) n1848 <= n5848;
/* FF  3 18  2 */ assign n460 = n5849;
/* FF 10 16  6 */ assign n1364 = n5850;
/* FF  7  1  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n825 <= 1'b0; else if (n663) n825 <= n5851;
/* FF 18 19  7 */ assign n2575 = n5852;
/* FF  9 12  5 */ assign n1170 = n5853;
/* FF  1 15  3 */ assign n115 = n5854;
/* FF 13 16  4 */ always @(posedge io_13_31_1) if (1'b1) n1783 <= n1973 ? 1'b0 : n5855;
/* FF  3 19  3 */ assign n469 = n5856;
/* FF 11 21  2 */ assign n1522 = n5857;
/* FF 16  3  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1727 <= 1'b0; else if (n1690) n1727 <= n5858;
/* FF 12 17  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1635 <= 1'b0; else if (1'b1) n1635 <= n5859;
/* FF 10 17  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1328 <= 1'b0; else if (n1502) n1328 <= n5860;
/* FF 20  6  4 */ always @(posedge io_13_31_1) if (n2676) n2680 <= n1 ? 1'b0 : n5861;
/* FF 10  9  3 */ assign n1296 = n5862;
/* FF  9 13  6 */ always @(posedge io_13_31_1) if (n4) n1177 <= 1'b0 ? 1'b0 : n5863;
/* FF 18 11  2 */ assign n2514 = n5864;
/* FF  9  5  2 */ assign n1109 = n5865;
/* FF 21 19  4 */ always @(posedge io_13_31_1) if (n2861) n2860 <= 1'b0 ? 1'b0 : n5866;
/* FF 13  8  5 */ assign n1736 = n5867;
/* FF 18 20  7 */ assign n1837 = n5868;
/* FF 18 12  3 */ always @(posedge io_13_31_1) if (n2137) n2524 <= n3 ? 1'b0 : n5869;
/* FF 10  1  4 */ assign n1238 = n5870;
/* FF 12 12  6 */ assign n1607 = n5871;
/* FF 22 15  6 */ always @(posedge io_13_31_1) if (1'b1) n2976 <= n3025 ? 1'b0 : n5872;
/* FF  2  7  1 */ assign n218 = n5873;
/* FF 21 11  5 */ always @(posedge io_13_31_1) if (n2213) n2499 <= 1'b0 ? 1'b0 : n5874;
/* FF 21  3  1 */ assign n5875 = n5876;
/* FF  1  3  6 */ assign n24 = n5877;
/* FF 14 21  3 */ assign n2020 = n5878;
/* FF 11  6  0 */ assign n1426 = n5879;
/* FF 13  4  7 */ assign n1687 = n5880;
/* FF  5 20  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n621 <= 1'b0; else if (n629) n621 <= n5881;
/* FF 17 21  1 */ assign n2429 = n5882;
/* FF 11  9  5 */ always @(posedge io_13_31_1) if (n4) n1450 <= 1'b0 ? 1'b0 : n5883;
/* FF 12 13  7 */ always @(posedge io_13_31_1) if (n4) n1614 <= 1'b0 ? 1'b0 : n5884;
/* FF 12  5  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1301 <= 1'b0; else if (n1426) n1301 <= n5885;
/* FF  2  8  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n226 <= 1'b0; else if (n70) n226 <= n5886;
/* FF 13  1  1 */ assign n5887 = n5888;
/* FF  4 19  4 */ assign n626 = n5889;
/* FF 14 22  4 */ assign n2029 = n5890;
/* FF  2 11  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n91 <= 1'b0; else if (1'b1) n91 <= n5891;
/* FF 14 14  0 */ assign n1959 = n5892;
/* FF  3  7  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n400 <= 1'b0; else if (n224) n400 <= n5893;
/* FF 21  7  7 */ assign n5894 = n5895;
/* FF 11 10  6 */ assign n1461 = n5896;
/* FF  8 22  7 */ assign n1075 = n5897;
/* FF 15 13  3 */ assign n2117 = n5898;
/* FF  5 15  6 */ assign n451 = n5899;
/* FF 22  4  5 */ assign n2913 = n5900;
/* FF  4 11  5 */ assign n81 = n5901;
/* FF 11  2  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1398 <= 1'b0; else if (n1120) n1398 <= n5902;
/* FF  8 15  4 */ assign n5903 = n5904;
/* FF  8  7  0 */ assign n5905 = n5906;
/* FF 17 13  1 */ always @(posedge io_13_31_1) if (n2536) n2386 <= n1 ? 1'b0 : n5908;
/* FF 20 21  2 */ always @(posedge io_13_31_1) if (n2590) n2748 <= 1'b0 ? 1'b0 : n5909;
/* FF 14  9  6 */ always @(posedge io_13_31_1) if (n1739) n1930 <= 1'b0 ? 1'b0 : n5910;
/* FF 15  5  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1542 <= 1'b0; else if (n1869) n1542 <= n5911;
/* FF  5  8  3 */ assign n705 = n5912;
/* FF  4  4  2 */ assign n521 = n5913;
/* FF  7 11  1 */ always @(posedge io_13_31_1) if (n4) n882 <= 1'b0 ? 1'b0 : n5914;
/* FF 16 18  4 */ assign n2000 = n5915;
/* FF  4  7  7 */ assign n547 = n5916;
/* FF 16 10  0 */ always @(posedge io_13_31_1) if (n2112) n2221 <= 1'b0 ? 1'b0 : n5917;
/* FF 14 10  7 */ assign n1937 = n5918;
/* FF  8 11  6 */ always @(posedge io_13_31_1) if (n4) n1018 <= 1'b0 ? 1'b0 : n5919;
/* FF 14  2  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1864 <= 1'b0; else if (n1670) n1864 <= n5920;
/* FF  5  1  0 */ assign n649 = n5921;
/* FF  7 20  6 */ assign n5922 = n5923;
/* FF 17  9  3 */ assign n2359 = n5924;
/* FF  7 12  2 */ assign n886 = n5925;
/* FF  5  4  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n6 <= 1'b0; else if (n217) n6 <= n5926;
/* FF 16 11  1 */ always @(posedge io_13_31_1) if (n2076) n2230 <= 1'b0 ? 1'b0 : n5927;
/* FF 10 19  7 */ assign n1377 = n5928;
/* FF 16 14  6 */ assign n2254 = n5929;
/* FF  9 15  6 */ assign n1195 = n5930;
/* FF  1 10  0 */ assign n72 = n5931;
/* FF 17  2  0 */ assign n2170 = n5932;
/* FF  3 21  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n437 <= 1'b0; else if (1'b1) n437 <= n5933;
/* FF  8  3  7 */ assign n955 = n5934;
/* FF  1 13  5 */ assign n98 = n5935;
/* FF 12 20  1 */ assign n1654 = n5936;
/* FF 20  9  5 */ assign n2345 = n5937;
/* FF  9  7  1 */ assign n877 = n5938;
/* FF 13 19  4 */ assign n1819 = n5939;
/* FF 21 21  3 */ assign n2873 = n5940;
/* FF  1 14  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n110 <= 1'b0; else if (1'b1) n110 <= n5941;
/* FF 16  6  7 */ assign n2189 = n5942;
/* FF  1  6  2 */ assign n5943 = n5944;
/* FF 10 20  7 */ assign n909 = n5945;
/* FF 10 12  3 */ always @(posedge io_13_31_1) if (n1180) n1323 <= n1 ? 1'b0 : n5946;
/* FF  9  8  2 */ always @(posedge io_13_31_1) if (n4) n1129 <= 1'b0 ? 1'b0 : n5947;
/* FF 22 18  1 */ assign n2987 = n5948;
/* FF  2 18  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n309 <= 1'b0; else if (n310) n309 <= n5949;
/* FF 13 12  1 */ assign n1759 = n5950;
/* FF 21 14  0 */ always @(posedge io_13_31_1) if (n2842) n2829 <= 1'b0 ? 1'b0 : n5951;
/* FF 20 10  5 */ always @(posedge io_13_31_1) if (n2112) n2630 <= 1'b0 ? 1'b0 : n5952;
/* FF  3  6  0 */ assign n384 = n5953;
/* FF 10  5  0 */ assign n841 = n5954;
/* FF 12 16  2 */ assign n1033 = n5955;
/* FF 15 20  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1836 <= 1'b0; else if (n1815) n1836 <= n5956;
/* FF  3  9  5 */ assign n418 = n5957;
/* FF  2 10  1 */ assign n201 = n5958;
/* FF 18  8  0 */ always @(posedge io_13_31_1) if (n2120) n2488 <= 1'b0 ? 1'b0 : n5959;
/* FF 13  7  7 */ assign n1725 = n5960;
/* FF  3  2  2 */ assign n348 = n5961;
/* FF 11 12  5 */ assign n729 = n5962;
/* FF 18 11  5 */ always @(posedge io_13_31_1) if (n2137) n2517 <= n3 ? 1'b0 : n5963;
/* FF 12  8  3 */ assign n1580 = n5964;
/* FF 15 16  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1790 <= 1'b0; else if (n1811) n1790 <= n5965;
/* FF  4 14  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n297 <= 1'b0; else if (1'b1) n297 <= n5966;
/* FF  2 14  7 */ assign n284 = n5967;
/* FF 21  2  3 */ assign n2324 = n5968;
/* FF 11  5  2 */ assign n1419 = n5969;
/* FF 12  1  0 */ assign n5970 = n5971;
/* FF  5 19  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n777 <= 1'b0; else if (n474) n777 <= n5973;
/* FF 10  1  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1241 <= 1'b0; else if (n1120) n1241 <= n5974;
/* FF  4 15  1 */ assign n601 = n5975;
/* FF 12  4  5 */ assign n1546 = n5976;
/* FF 22  7  5 */ assign n2938 = n5977;
/* FF  2  7  4 */ assign n215 = n5978;
/* FF 21  3  4 */ always @(posedge io_13_31_1) if (n2902) n2764 <= n7 ? 1'b0 : n5979;
/* FF 14 21  6 */ assign n2012 = n5980;
/* FF 11  6  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1427 <= 1'b0; else if (n1426) n1427 <= n5981;
/* FF  8 10  0 */ always @(posedge io_13_31_1) if (n4) n1006 <= 1'b0 ? 1'b0 : n5982;
/* FF 15  9  0 */ assign n2077 = n5983;
/* FF 17 12  4 */ assign n2382 = n5984;
/* FF 17  4  0 */ always @(posedge io_13_31_1) if (n2316) n2325 <= 1'b0 ? 1'b0 : n5985;
/* FF 15  4  7 */ assign n2052 = n5986;
/* FF  5  6  4 */ assign n402 = n5987;
/* FF  4 10  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n567 <= 1'b0; else if (n576) n567 <= n5988;
/* FF 16 13  0 */ assign n2246 = n5989;
/* FF 14 13  7 */ assign n1955 = n5990;
/* FF  4  2  3 */ assign n504 = n5991;
/* FF  8 14  6 */ assign n1041 = n5992;
/* FF 14  5  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1887 <= 1'b0; else if (n1433) n1887 <= n5993;
/* FF 23 12  0 */ assign n5994 = n5995;
/* FF  7 15  2 */ assign n5997 = n5998;
/* FF  5  7  5 */ assign n694 = n5999;
/* FF  9 19  2 */ assign n1209 = n6000;
/* FF  4  3  4 */ assign n514 = n6001;
/* FF 16  9  2 */ assign n2216 = n6002;
/* FF 17 13  4 */ always @(posedge io_13_31_1) if (n2536) n2255 <= n1 ? 1'b0 : n6003;
/* FF 17  5  0 */ always @(posedge io_13_31_1) if (n2456) n2334 <= 1'b0 ? 1'b0 : n6004;
/* FF 20 13  1 */ assign n2707 = n6005;
/* FF  8  6  7 */ assign n224 = n6006;
/* FF 15  5  7 */ assign n1001 = n6007;
/* FF 10 15  4 */ assign n1355 = n6008;
/* FF 10  7  0 */ always @(posedge io_13_31_1) if (n4) n1272 <= 1'b0 ? 1'b0 : n6009;
/* FF 13 22  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1845 <= 1'b0; else if (n1666) n1845 <= n6010;
/* FF  2 21  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n324 <= 1'b0; else if (n160) n324 <= n6011;
/* FF 13 14  0 */ assign n1784 = n6012;
/* FF  1 17  6 */ assign n125 = n6013;
/* FF  1  9  2 */ assign n65 = n6014;
/* FF 20  5  2 */ always @(posedge io_13_31_1) if (n2472) n2673 <= n2471 ? 1'b0 : n6015;
/* FF  9 11  2 */ always @(posedge io_13_31_1) if (n4) n1160 <= 1'b0 ? 1'b0 : n6016;
/* FF 12 19  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1647 <= 1'b0; else if (n1815) n1647 <= n6017;
/* FF 18 10  0 */ assign n2503 = n6018;
/* FF 13 15  1 */ assign n1795 = n6019;
/* FF  7  3  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n836 <= 1'b0; else if (n663) n836 <= n6020;
/* FF 10 11  6 */ assign n1316 = n6021;
/* FF 13 18  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1780 <= 1'b0; else if (n1967) n1780 <= n6022;
/* FF 10  8  0 */ assign n1282 = n6023;
/* FF 21 21  6 */ assign n2848 = n6024;
/* FF  4 17  1 */ assign n612 = n6025;
/* FF 11 16  1 */ assign n1497 = n6026;
/* FF 13 10  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1728 <= 1'b0; else if (n734) n1728 <= n6027;
/* FF  2  9  4 */ assign n240 = n6028;
/* FF 13  2  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1669 <= 1'b0; else if (n1670) n1669 <= n6029;
/* FF  3 13  6 */ assign n278 = n6030;
/* FF  3  5  2 */ assign n375 = n6031;
/* FF 14 23  6 */ assign n2036 = n6032;
/* FF 15 19  4 */ assign n2146 = n6033;
/* FF 15 11  0 */ assign n2094 = n6034;
/* FF 10  3  6 */ assign n1256 = n6035;
/* FF 12  7  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1573 <= 1'b0; else if (n1279) n1573 <= n6036;
/* FF 14 20  0 */ always @(posedge io_13_31_1) if (n1838) n2006 <= n2155 ? 1'b0 : n6037;
/* FF 22  9  4 */ always @(posedge io_13_31_1) if (n2686) n2951 <= 1'b0 ? 1'b0 : n6038;
/* FF 13  3  4 */ assign n1675 = n6039;
/* FF 21 13  7 */ assign n2825 = n6040;
/* FF  3  6  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n382 <= 1'b0; else if (n224) n382 <= n6041;
/* FF 21  5  3 */ always @(posedge io_13_31_1) if (n2902) n2779 <= n7 ? 1'b0 : n6042;
/* FF  4 21  7 */ assign n644 = n6043;
/* FF 11  8  2 */ always @(posedge io_13_31_1) if (n4) n1437 <= 1'b0 ? 1'b0 : n6044;
/* FF 15 20  5 */ assign n2154 = n6045;
/* FF 15 12  1 */ assign n2106 = n6046;
/* FF 23 14  0 */ always @(posedge io_13_31_1) if (1'b1) n3019 <= 1'b0 ? 1'b0 : n6047;
/* FF  4 18  1 */ assign n6048 = n6049;
/* FF 22 10  5 */ always @(posedge io_13_31_1) if (n2113) n2196 <= 1'b0 ? 1'b0 : n6050;
/* FF  2 10  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n247 <= 1'b0; else if (1'b1) n247 <= n6051;
/* FF 22  2  1 */ always @(posedge io_13_31_1) if (1'b1) n2887 <= 1'b0 ? 1'b0 : n6052;
/* FF  2  2  0 */ assign n167 = n6053;
/* FF 21  6  4 */ always @(posedge io_13_31_1) if (n2686) n2455 <= 1'b0 ? 1'b0 : n6054;
/* FF  8 13  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1025 <= 1'b0; else if (n1166) n1025 <= n6055;
/* FF 11  4  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1409 <= 1'b0; else if (n979) n1409 <= n6056;
/* FF 22  3  2 */ always @(posedge io_13_31_1) if (1'b1) n2896 <= n2757 ? 1'b0 : n6057;
/* FF 17 15  4 */ always @(posedge io_13_31_1) if (1'b1) n2397 <= n2138 ? 1'b0 : n6058;
/* FF  7 18  3 */ assign n6059 = n6060;
/* FF 22  6  7 */ always @(posedge io_13_31_1) if (1'b1) n179 <= 1'b0 ? 1'b0 : n6061;
/* FF 15  7  7 */ assign n2064 = n6062;
/* FF  9 21  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1189 <= 1'b0; else if (n1068) n1189 <= n6063;
/* FF  8 17  6 */ assign n6064 = n6065;
/* FF 14  8  3 */ assign n1920 = n6066;
/* FF  8  9  2 */ assign n997 = n6067;
/* FF 23 11  3 */ always @(posedge io_13_31_1) if (n2826) n2500 <= n2395 ? 1'b1 : n6068;
/* FF 20 23  4 */ always @(posedge io_13_31_1) if (n2754) n2586 <= 1'b0 ? 1'b0 : n6069;
/* FF 17  8  1 */ always @(posedge io_13_31_1) if (n2344) n2348 <= 1'b0 ? 1'b0 : n6070;
/* FF  9 22  2 */ assign n1229 = n6071;
/* FF 17 11  6 */ assign n2111 = n6072;
/* FF  4  6  4 */ assign n534 = n6073;
/* FF  8 10  3 */ always @(posedge io_13_31_1) if (n4) n1008 <= 1'b0 ? 1'b0 : n6074;
/* FF 14  1  0 */ assign n1860 = n6075;
/* FF 16 20  6 */ assign n2024 = n6076;
/* FF  1 20  1 */ assign n143 = n6077;
/* FF 16 12  2 */ assign n2239 = n6078;
/* FF 14  4  5 */ assign n1433 = n6079;
/* FF 10 19  0 */ assign n1373 = n6080;
/* FF  1 19  5 */ assign n139 = n6081;
/* FF  5  3  2 */ assign n664 = n6082;
/* FF 23  3  4 */ assign n3009 = n6083;
/* FF 17  4  3 */ always @(posedge io_13_31_1) if (n2316) n2328 <= 1'b0 ? 1'b0 : n6084;
/* FF  5  6  7 */ assign n691 = n6085;
/* FF 16 13  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1757 <= 1'b0; else if (n735) n1757 <= n6086;
/* FF  4  2  6 */ assign n507 = n6087;
/* FF 14  5  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1888 <= 1'b0; else if (n1433) n1888 <= n6088;
/* FF  1 12  2 */ assign n84 = n6089;
/* FF 13 21  7 */ assign n1835 = n6090;
/* FF 20  8  2 */ assign n2688 = n6091;
/* FF 12 22  3 */ assign n1661 = n6092;
/* FF 20 11  7 */ assign n2702 = n6093;
/* FF 10 14  6 */ always @(posedge io_13_31_1) if (n4) n1347 <= 1'b0 ? 1'b0 : n6094;
/* FF 10  6  2 */ assign n1267 = n6095;
/* FF  9 10  5 */ always @(posedge io_13_31_1) if (n4) n1156 <= 1'b0 ? 1'b0 : n6096;
/* FF  9  2  1 */ assign n1083 = n6097;
/* FF 22 20  4 */ assign n2751 = n6098;
/* FF  3 16  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n446 <= 1'b0; else if (1'b1) n446 <= n6099;
/* FF 21 16  3 */ assign n2845 = n6100;
/* FF 12 15  0 */ always @(posedge io_13_31_1) if (n1180) n1628 <= n1 ? 1'b0 : n6101;
/* FF 20  4  4 */ assign n2316 = n6102;
/* FF 10 15  7 */ assign n1357 = n6103;
/* FF 10  7  3 */ assign n1275 = n6104;
/* FF 18 17  6 */ assign n2560 = n6105;
/* FF 18  9  2 */ assign n2493 = n6106;
/* FF  3  8  2 */ assign n404 = n6107;
/* FF 18 10  3 */ assign n2505 = n6108;
/* FF  9  3  1 */ assign n1092 = n6109;
/* FF 15 22  4 */ always @(posedge io_13_31_1) if (n2037) n2158 <= 1'b0 ? 1'b0 : n6110;
/* FF  3 11  7 */ assign n391 = n6111;
/* FF 15 14  0 */ assign n2124 = n6112;
/* FF 21 17  3 */ assign n2849 = n6113;
/* FF  2 13  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n113 <= 1'b0; else if (n432) n113 <= n6114;
/* FF 12  2  2 */ assign n1530 = n6115;
/* FF 13  6  4 */ assign n1711 = n6116;
/* FF  4 16  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n608 <= 1'b0; else if (1'b1) n608 <= n6117;
/* FF 11 11  2 */ assign n1466 = n6118;
/* FF 14 19  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1983 <= 1'b0; else if (n1527) n1983 <= n6119;
/* FF 22  8  7 */ assign n2947 = n6120;
/* FF 15 15  1 */ assign n6121 = n6122;
/* FF  3  4  4 */ assign n367 = n6123;
/* FF 21  4  6 */ always @(posedge io_13_31_1) if (n2902) n2774 <= n7 ? 1'b0 : n6124;
/* FF 15 18  6 */ assign n2141 = n6125;
/* FF 12  3  3 */ assign n6126 = n6127;
/* FF 22  5  1 */ assign n2926 = n6128;
/* FF  5 13  1 */ assign n444 = n6129;
/* FF  4 17  4 */ assign n258 = n6130;
/* FF 21  1  0 */ assign n2756 = n6131;
/* FF  2  9  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n235 <= 1'b0; else if (1'b1) n235 <= n6132;
/* FF 13  2  6 */ assign n1263 = n6133;
/* FF 17 19  0 */ assign n6134 = n6135;
/* FF 11  7  4 */ assign n1431 = n6137;
/* FF  8 20  7 */ assign n1064 = n6138;
/* FF 15 11  3 */ assign n2097 = n6139;
/* FF 14 20  3 */ always @(posedge io_13_31_1) if (n1838) n2008 <= n2155 ? 1'b0 : n6140;
/* FF 15 10  7 */ assign n2091 = n6141;
/* FF 22  9  7 */ always @(posedge io_13_31_1) if (n2686) n2953 <= 1'b0 ? 1'b0 : n6142;
/* FF 21  5  6 */ always @(posedge io_13_31_1) if (n2902) n2782 <= n7 ? 1'b0 : n6143;
/* FF  5  5  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n683 <= 1'b0; else if (n524) n683 <= n6144;
/* FF  4  1  1 */ assign n493 = n6145;
/* FF  8 12  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1021 <= 1'b0; else if (n1166) n1021 <= n6146;
/* FF 16 15  3 */ always @(posedge io_13_31_1) if (n2268) n2260 <= 1'b0 ? 1'b0 : n6147;
/* FF 20 18  0 */ assign n1518 = n6148;
/* FF 15  3  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1701 <= 1'b0; else if (n1547) n1701 <= n6149;
/* FF 17 14  6 */ always @(posedge io_13_31_1) if (n2396) n2393 <= n1 ? 1'b0 : n6150;
/* FF  7 17  5 */ assign n916 = n6151;
/* FF  7  9  1 */ assign n873 = n6152;
/* FF  2  1  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n166 <= 1'b0; else if (n178) n166 <= n6153;
/* FF  8 13  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1026 <= 1'b0; else if (n1166) n1026 <= n6154;
/* FF  4  5  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n390 <= 1'b0; else if (n524) n390 <= n6155;
/* FF 20 19  1 */ assign n2739 = n6156;
/* FF 14  7  5 */ assign n1910 = n6157;
/* FF 17 15  7 */ assign n2275 = n6158;
/* FF 17  7  3 */ assign n2343 = n6159;
/* FF  9 21  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n907 <= 1'b0; else if (n1068) n907 <= n6160;
/* FF 14  8  6 */ assign n1916 = n6161;
/* FF  1 15  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n114 <= 1'b0; else if (n115) n114 <= n6162;
/* FF 13 16  3 */ assign n1804 = n6163;
/* FF  3 19  2 */ assign n468 = n6164;
/* FF 23  2  6 */ assign n6165 = n6166;
/* FF 20 14  7 */ assign n2719 = n6167;
/* FF 10  9  2 */ assign n1295 = n6168;
/* FF  9 13  5 */ always @(posedge io_13_31_1) if (n4) n908 <= 1'b0 ? 1'b0 : n6169;
/* FF  9  5  1 */ assign n362 = n6170;
/* FF 13 17  4 */ assign n1809 = n6171;
/* FF 16  4  1 */ assign n2173 = n6172;
/* FF  8  1  6 */ assign n939 = n6173;
/* FF 21 19  3 */ assign n2855 = n6174;
/* FF 12 18  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1640 <= 1'b0; else if (1'b1) n1640 <= n6175;
/* FF 20  7  4 */ assign n2685 = n6176;
/* FF 10 10  3 */ assign n1305 = n6177;
/* FF 12 21  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1391 <= 1'b0; else if (n1658) n1391 <= n6178;
/* FF 18 12  2 */ always @(posedge io_13_31_1) if (n2137) n2523 <= n3 ? 1'b0 : n6179;
/* FF  9  6  2 */ assign n861 = n6180;
/* FF  2 16  0 */ assign n292 = n6181;
/* FF 21 20  4 */ assign n2864 = n6182;
/* FF  9  9  7 */ always @(posedge io_13_31_1) if (n4) n1143 <= 1'b0 ? 1'b0 : n6183;
/* FF 21 12  0 */ always @(posedge io_13_31_1) if (n2663) n2811 <= 1'b0 ? 1'b0 : n6184;
/* FF  1  4  1 */ assign n28 = n6185;
/* FF 20  8  5 */ assign n2683 = n6186;
/* FF 18 13  3 */ always @(posedge io_13_31_1) if (n2137) n2531 <= n3 ? 1'b0 : n6187;
/* FF  1  3  5 */ assign n23 = n6188;
/* FF 12 14  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1618 <= 1'b0; else if (n1630) n1618 <= n6189;
/* FF 12 13  6 */ always @(posedge io_13_31_1) if (n4) n1182 <= 1'b0 ? 1'b0 : n6190;
/* FF 22 20  7 */ assign n2995 = n6191;
/* FF  2  8  1 */ assign n6192 = n6193;
/* FF 13  1  0 */ assign n6194 = n6195;
/* FF  4 19  3 */ assign n6197 = n6198;
/* FF 14 22  3 */ assign n2028 = n6199;
/* FF 18  6  0 */ assign n6200 = n6201;
/* FF  2 11  6 */ assign n256 = n6203;
/* FF  3  7  4 */ assign n399 = n6204;
/* FF 11 10  5 */ assign n1460 = n6205;
/* FF 18  9  5 */ always @(posedge io_13_31_1) if (n2076) n2496 <= 1'b0 ? 1'b0 : n6206;
/* FF 12  6  3 */ assign n1559 = n6207;
/* FF 15 13  2 */ assign n2116 = n6208;
/* FF  4 20  4 */ assign n638 = n6209;
/* FF  4 12  0 */ assign n6210 = n6211;
/* FF  2 12  7 */ assign n263 = n6213;
/* FF 13  5  6 */ assign n1697 = n6214;
/* FF 14 15  0 */ assign n1968 = n6215;
/* FF  2  4  3 */ always @(posedge io_13_31_1) if (n201) n194 <= n42 ? 1'b0 : n6216;
/* FF  3  8  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n407 <= 1'b0; else if (n71) n407 <= n6217;
/* FF 21  8  7 */ always @(posedge io_13_31_1) if (n2694) n2804 <= n1 ? 1'b0 : n6218;
/* FF 22  4  4 */ assign n2912 = n6219;
/* FF 14 18  5 */ assign n1996 = n6220;
/* FF 11  2  0 */ assign n1397 = n6221;
/* FF 15 14  3 */ assign n2126 = n6222;
/* FF  4 13  1 */ assign n6223 = n6224;
/* FF  4 16  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n452 <= 1'b0; else if (1'b1) n452 <= n6225;
/* FF 11 11  5 */ always @(posedge io_13_31_1) if (n4) n1468 <= 1'b0 ? 1'b0 : n6226;
/* FF 11  3  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1403 <= 1'b0; else if (n979) n1403 <= n6227;
/* FF 14 11  2 */ assign n1939 = n6228;
/* FF  8 11  5 */ assign n1017 = n6229;
/* FF  7 20  5 */ assign n6230 = n6231;
/* FF  7 12  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n885 <= 1'b0; else if (n818) n885 <= n6232;
/* FF  5  4  4 */ assign n675 = n6233;
/* FF  4  8  7 */ assign n554 = n6234;
/* FF 16 11  0 */ assign n2110 = n6235;
/* FF 16 14  5 */ assign n2251 = n6236;
/* FF 17 18  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2415 <= 1'b0; else if (n2011) n2415 <= n6237;
/* FF 17 10  3 */ always @(posedge io_13_31_1) if (n2213) n2367 <= 1'b0 ? 1'b0 : n6238;
/* FF  7 13  2 */ always @(posedge io_13_31_1) if (n4) n896 <= 1'b0 ? 1'b0 : n6239;
/* FF 15  2  6 */ assign n2047 = n6240;
/* FF  5  5  5 */ assign n685 = n6241;
/* FF  9 16  0 */ assign n6242 = n6243;
/* FF  7 16  7 */ assign n821 = n6245;
/* FF  4  1  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n496 <= 1'b0; else if (n656) n496 <= n6246;
/* FF 14  3  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1871 <= 1'b0; else if (n1690) n1871 <= n6247;
/* FF  8  4  1 */ assign n962 = n6248;
/* FF 16 15  6 */ always @(posedge io_13_31_1) if (n2268) n2263 <= 1'b0 ? 1'b0 : n6249;
/* FF 16  7  2 */ always @(posedge io_13_31_1) if (n2093) n2199 <= 1'b0 ? 1'b0 : n6250;
/* FF 13 19  3 */ assign n1818 = n6251;
/* FF 20 18  3 */ assign n2730 = n6252;
/* FF 17  3  0 */ always @(posedge io_13_31_1) if (n2324) n2317 <= 1'b0 ? 1'b0 : n6253;
/* FF 23  5  6 */ always @(posedge io_13_31_1) if (1'b1) n1 <= n2927 ? 1'b0 : n6254;
/* FF  1 14  5 */ assign n109 = n6255;
/* FF  1  6  1 */ assign n6256 = n6257;
/* FF 10 20  6 */ assign n1381 = n6258;
/* FF  9  8  1 */ always @(posedge io_13_31_1) if (n4) n1121 <= 1'b0 ? 1'b0 : n6259;
/* FF 13 20  4 */ assign n1828 = n6260;
/* FF 13 12  0 */ assign n1758 = n6261;
/* FF  3 18  4 */ assign n457 = n6262;
/* FF 20  2  0 */ always @(posedge io_13_31_1) if (n2324) n2668 <= 1'b0 ? 1'b0 : n6263;
/* FF 12 16  1 */ always @(posedge io_13_31_1) if (n4) n1634 <= 1'b0 ? 1'b0 : n6264;
/* FF 22 19  1 */ always @(posedge io_13_31_1) if (n2747) n2728 <= 1'b0 ? 1'b0 : n6265;
/* FF  2 19  0 */ assign n6266 = n6267;
/* FF  7  1  5 */ assign n826 = n6269;
/* FF 13 13  1 */ always @(posedge io_13_31_1) if (1'b1) n1771 <= 1'b0 ? 1'b0 : n6270;
/* FF  9 12  7 */ assign n1166 = n6271;
/* FF 21 15  0 */ assign n2827 = n6272;
/* FF  1  7  1 */ assign n46 = n6273;
/* FF 13 16  6 */ assign n1806 = n6274;
/* FF 20  3  1 */ always @(posedge io_13_31_1) if (1'b1) n177 <= 1'b0 ? 1'b0 : n6275;
/* FF 11 21  4 */ assign n1523 = n6276;
/* FF 12 17  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1636 <= 1'b1; else if (1'b1) n1636 <= n6277;
/* FF 20  6  6 */ always @(posedge io_13_31_1) if (n2676) n2682 <= n1 ? 1'b0 : n6278;
/* FF 10  9  5 */ always @(posedge io_13_31_1) if (n4) n1298 <= 1'b0 ? 1'b0 : n6279;
/* FF 18 11  4 */ always @(posedge io_13_31_1) if (n2137) n2516 <= n3 ? 1'b0 : n6280;
/* FF  9  5  4 */ assign n1111 = n6281;
/* FF 11 14  1 */ always @(posedge io_13_31_1) if (n1180) n1480 <= n1 ? 1'b0 : n6282;
/* FF  2 14  6 */ assign n117 = n6283;
/* FF 13  8  7 */ assign n1717 = n6284;
/* FF 11 13  5 */ assign n1476 = n6285;
/* FF 18 12  5 */ always @(posedge io_13_31_1) if (n2137) n2526 <= n3 ? 1'b0 : n6286;
/* FF 18  4  1 */ always @(posedge io_13_31_1) if (n2603) n2451 <= 1'b0 ? 1'b0 : n6287;
/* FF  5 19  1 */ assign n783 = n6288;
/* FF 10  1  6 */ assign n1240 = n6289;
/* FF 24 15  1 */ always @(posedge io_13_31_1) if (n2981) n2983 <= 1'b0 ? 1'b0 : n6290;
/* FF  4 15  0 */ assign n600 = n6291;
/* FF  2 15  7 */ assign n121 = n6292;
/* FF 12  4  4 */ assign n1545 = n6293;
/* FF 22  7  4 */ assign n2937 = n6294;
/* FF  2  7  3 */ assign n220 = n6295;
/* FF  3  3  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n356 <= 1'b0; else if (n198) n356 <= n6296;
/* FF 21  3  3 */ always @(posedge io_13_31_1) if (n2902) n2763 <= n7 ? 1'b0 : n6297;
/* FF 14 21  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2021 <= 1'b0; else if (1'b1) n2021 <= n6298;
/* FF 11  6  2 */ assign n1424 = n6299;
/* FF  5 20  2 */ assign n792 = n6300;
/* FF 17 21  3 */ always @(posedge io_13_31_1) if (n2423) n2430 <= 1'b0 ? 1'b0 : n6301;
/* FF 11  9  7 */ assign n1451 = n6302;
/* FF 12  5  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1270 <= 1'b0; else if (n1426) n1270 <= n6303;
/* FF  2  8  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n230 <= 1'b0; else if (n70) n230 <= n6304;
/* FF 13  1  3 */ assign n6305 = n6306;
/* FF  4 19  6 */ assign n628 = n6307;
/* FF 14 22  6 */ assign n2030 = n6308;
/* FF 14 14  2 */ assign n1958 = n6309;
/* FF 15 10  0 */ always @(posedge io_13_31_1) if (n1591) n2085 <= 1'b0 ? 1'b0 : n6310;
/* FF  8 14  5 */ assign n1040 = n6311;
/* FF 15 13  5 */ assign n2118 = n6312;
/* FF 23 16  6 */ always @(posedge io_13_31_1) if (n2859) n2854 <= 1'b0 ? 1'b0 : n6313;
/* FF  7 15  1 */ assign n6314 = n6315;
/* FF  5  7  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n693 <= 1'b0; else if (n532) n693 <= n6316;
/* FF  9 19  1 */ assign n797 = n6317;
/* FF  4 11  7 */ assign n265 = n6318;
/* FF 23 13  0 */ always @(posedge io_13_31_1) if (n2842) n3016 <= 1'b0 ? 1'b0 : n6319;
/* FF 11  2  3 */ assign n1400 = n6320;
/* FF  4  3  3 */ assign n513 = n6321;
/* FF  8 15  6 */ assign n6322 = n6323;
/* FF  8  7  2 */ assign n6324 = n6325;
/* FF 16 17  5 */ assign n1513 = n6326;
/* FF 17 13  3 */ always @(posedge io_13_31_1) if (n2536) n2387 <= n1 ? 1'b0 : n6327;
/* FF 20 13  0 */ always @(posedge io_13_31_1) if (n2663) n2706 <= 1'b0 ? 1'b0 : n6328;
/* FF 15  5  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1714 <= 1'b0; else if (n1869) n1714 <= n6329;
/* FF  5  8  5 */ assign n707 = n6330;
/* FF  7 19  7 */ assign n648 = n6331;
/* FF 16 18  6 */ assign n2143 = n6332;
/* FF 16 10  2 */ assign n2223 = n6333;
/* FF 17  6  0 */ assign n6334 = n6335;
/* FF 14  2  5 */ assign n1866 = n6337;
/* FF  9 20  1 */ assign n6338 = n6339;
/* FF  1 17  5 */ assign n124 = n6340;
/* FF 17  9  5 */ assign n2361 = n6341;
/* FF  7 12  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n888 <= 1'b0; else if (n818) n888 <= n6342;
/* FF  7  4  0 */ assign n500 = n6343;
/* FF 13 15  0 */ assign n6344 = n6345;
/* FF 10 11  5 */ always @(posedge io_13_31_1) if (n4) n1315 <= 1'b0 ? 1'b0 : n6347;
/* FF 13 18  5 */ assign n1814 = n6348;
/* FF  3 21  4 */ assign n484 = n6349;
/* FF  1 13  7 */ assign n100 = n6350;
/* FF 20  9  7 */ always @(posedge io_13_31_1) if (n2093) n2502 <= 1'b0 ? 1'b0 : n6351;
/* FF 21 18  0 */ always @(posedge io_13_31_1) if (n2666) n2857 <= 1'b0 ? 1'b0 : n6352;
/* FF 13 19  6 */ assign n1821 = n6353;
/* FF 13 11  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1740 <= 1'b0; else if (n734) n1740 <= n6354;
/* FF 21 21  5 */ assign n2869 = n6355;
/* FF  3 14  1 */ assign n6356 = n6357;
/* FF 11 16  0 */ always @(posedge io_13_31_1) if (n4) n1496 <= 1'b0 ? 1'b0 : n6358;
/* FF  1  6  4 */ assign n6359 = n6360;
/* FF 10 12  5 */ always @(posedge io_13_31_1) if (n1180) n1325 <= n1 ? 1'b0 : n6361;
/* FF 10  4  1 */ assign n1107 = n6362;
/* FF  9  8  4 */ always @(posedge io_13_31_1) if (n4) n1131 <= 1'b0 ? 1'b0 : n6363;
/* FF 22 18  3 */ assign n2989 = n6364;
/* FF  2 18  2 */ assign n311 = n6365;
/* FF 21 14  2 */ always @(posedge io_13_31_1) if (n2842) n2831 <= 1'b0 ? 1'b0 : n6366;
/* FF 13  3  3 */ assign n1674 = n6367;
/* FF  3  6  2 */ assign n386 = n6368;
/* FF 18 15  5 */ assign n2402 = n6369;
/* FF  3  9  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n419 <= 1'b1; else if (n70) n419 <= n6370;
/* FF 15 12  0 */ assign n2105 = n6371;
/* FF 17 23  2 */ assign n2437 = n6372;
/* FF  4 18  0 */ assign n6373 = n6374;
/* FF 22 10  4 */ assign n2954 = n6376;
/* FF  2 10  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n246 <= 1'b0; else if (1'b1) n246 <= n6377;
/* FF  5 18  4 */ assign n776 = n6378;
/* FF 21  6  3 */ always @(posedge io_13_31_1) if (n2686) n2484 <= 1'b0 ? 1'b0 : n6379;
/* FF 14 16  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1978 <= 1'b0; else if (n1967) n1978 <= n6380;
/* FF  3  2  4 */ assign n350 = n6381;
/* FF 11 12  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1330 <= 1'b0; else if (n102) n1330 <= n6382;
/* FF 23 15  0 */ assign n3025 = n6383;
/* FF 11  4  3 */ assign n1412 = n6384;
/* FF 12  8  5 */ assign n1581 = n6385;
/* FF 15 16  6 */ assign n1811 = n6386;
/* FF  2  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n180 <= 1'b0; else if (n17) n180 <= n6387;
/* FF  4 14  2 */ assign n592 = n6388;
/* FF  8 18  1 */ assign n1052 = n6389;
/* FF 21  2  5 */ assign n2758 = n6390;
/* FF 11  5  4 */ assign n1120 = n6391;
/* FF  8 17  5 */ assign n6392 = n6393;
/* FF 12  1  2 */ assign n6394 = n6395;
/* FF  5 11  0 */ assign n6396 = n6397;
/* FF 12  4  7 */ assign n973 = n6399;
/* FF 15  8  7 */ assign n2075 = n6400;
/* FF 22  7  7 */ assign n2939 = n6401;
/* FF  9 22  1 */ assign n1228 = n6402;
/* FF 21  3  6 */ always @(posedge io_13_31_1) if (n2902) n2766 <= n7 ? 1'b0 : n6403;
/* FF 16 21  1 */ assign n2037 = n6404;
/* FF  7 14  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n905 <= 1'b0; else if (1'b1) n905 <= n6405;
/* FF  8 10  2 */ assign n711 = n6406;
/* FF  1 20  0 */ assign n6407 = n6408;
/* FF  5  3  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n666 <= 1'b0; else if (n198) n666 <= n6410;
/* FF 17  4  2 */ always @(posedge io_13_31_1) if (n2316) n2327 <= 1'b0 ? 1'b0 : n6411;
/* FF  5  6  6 */ always @(posedge io_13_31_1) if (n4) n690 <= 1'b0 ? 1'b0 : n6412;
/* FF  1 21  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n152 <= 1'b0; else if (n80) n152 <= n6413;
/* FF 16 13  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1755 <= 1'b0; else if (n735) n1755 <= n6414;
/* FF  4  2  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n506 <= 1'b0; else if (n509) n506 <= n6415;
/* FF 14  5  5 */ assign n807 = n6416;
/* FF 16 16  7 */ assign n2268 = n6417;
/* FF  7 15  4 */ assign n6418 = n6419;
/* FF  7  7  0 */ assign n853 = n6420;
/* FF  5  7  7 */ assign n697 = n6421;
/* FF  9 19  4 */ assign n1207 = n6422;
/* FF  4  3  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n516 <= 1'b0; else if (n509) n516 <= n6423;
/* FF 16  9  4 */ always @(posedge io_13_31_1) if (n2093) n2092 <= 1'b0 ? 1'b0 : n6424;
/* FF 17  5  2 */ always @(posedge io_13_31_1) if (n2456) n2336 <= 1'b0 ? 1'b0 : n6425;
/* FF  3 16  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n445 <= 1'b0; else if (1'b1) n445 <= n6426;
/* FF 18 18  1 */ assign n2562 = n6427;
/* FF 20 12  7 */ always @(posedge io_13_31_1) if (n2112) n2373 <= 1'b0 ? 1'b0 : n6428;
/* FF 10 15  6 */ always @(posedge io_13_31_1) if (n4) n1356 <= 1'b0 ? 1'b0 : n6429;
/* FF 10  7  2 */ assign n1274 = n6430;
/* FF 13 22  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1847 <= 1'b0; else if (n1666) n1847 <= n6431;
/* FF 22 21  4 */ assign n3001 = n6432;
/* FF  2 21  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n331 <= 1'b0; else if (n160) n331 <= n6433;
/* FF 13 14  2 */ assign n1494 = n6434;
/* FF 22 13  0 */ always @(posedge io_13_31_1) if (n2663) n2958 <= 1'b0 ? 1'b0 : n6435;
/* FF  3 17  1 */ assign n131 = n6436;
/* FF 16  1  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2167 <= 1'b1; else if (1'b1) n2167 <= n6437;
/* FF  9 11  4 */ always @(posedge io_13_31_1) if (n4) n1162 <= 1'b0 ? 1'b0 : n6438;
/* FF 18 10  2 */ assign n2384 = n6439;
/* FF  9  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1091 <= 1'b0; else if (n851) n1091 <= n6440;
/* FF 12 11  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1592 <= 1'b0; else if (n734) n1592 <= n6441;
/* FF  7  3  7 */ assign n839 = n6442;
/* FF 13 15  3 */ assign n1792 = n6443;
/* FF 11 20  1 */ assign n1519 = n6444;
/* FF 10  8  2 */ always @(posedge io_13_31_1) if (n4) n1284 <= 1'b0 ? 1'b0 : n6445;
/* FF  9  4  1 */ assign n1101 = n6446;
/* FF 22 22  4 */ always @(posedge io_13_31_1) if (n2593) n2883 <= 1'b0 ? 1'b0 : n6447;
/* FF 22 14  0 */ assign n6448 = n6449;
/* FF 21 18  3 */ assign n2858 = n6451;
/* FF  9  7  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n209 <= 1'b0; else if (n877) n209 <= n6452;
/* FF 12  3  2 */ assign n6453 = n6454;
/* FF  5 13  0 */ assign n606 = n6455;
/* FF  4 17  3 */ assign n597 = n6456;
/* FF 11 16  3 */ always @(posedge io_13_31_1) if (n4) n1486 <= 1'b0 ? 1'b0 : n6457;
/* FF  2  9  6 */ assign n242 = n6458;
/* FF 13  2  5 */ assign n1417 = n6459;
/* FF  3  5  4 */ assign n377 = n6460;
/* FF 11 15  7 */ assign n1493 = n6461;
/* FF 15 11  2 */ assign n2096 = n6462;
/* FF  2  6  0 */ assign n6463 = n6464;
/* FF  5 14  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n753 <= 1'b0; else if (1'b1) n753 <= n6466;
/* FF 14 20  2 */ always @(posedge io_13_31_1) if (n1838) n2007 <= n2155 ? 1'b0 : n6467;
/* FF  8 21  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n931 <= 1'b0; else if (n1068) n931 <= n6468;
/* FF 13  3  6 */ assign n1676 = n6469;
/* FF 22  9  6 */ always @(posedge io_13_31_1) if (n2686) n2952 <= 1'b0 ? 1'b0 : n6470;
/* FF 21  5  5 */ always @(posedge io_13_31_1) if (n2902) n2781 <= n7 ? 1'b0 : n6471;
/* FF 17 20  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n2297 <= 1'b0; else if (n2023) n2297 <= n6472;
/* FF 11  8  4 */ always @(posedge io_13_31_1) if (n4) n1439 <= 1'b0 ? 1'b0 : n6473;
/* FF 15 12  3 */ assign n2103 = n6474;
/* FF 23 14  2 */ always @(posedge io_13_31_1) if (1'b1) n3021 <= 1'b0 ? 1'b0 : n6475;
/* FF  4 18  3 */ assign n6476 = n6477;
/* FF  2 10  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n93 <= 1'b0; else if (1'b1) n93 <= n6478;
/* FF 22  2  3 */ assign n2889 = n6479;
/* FF  2  2  2 */ assign n169 = n6480;
/* FF 21  6  6 */ always @(posedge io_13_31_1) if (n2686) n2454 <= 1'b0 ? 1'b0 : n6481;
/* FF 11  1  1 */ assign n6482 = n6483;
/* FF  8 13  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1023 <= 1'b1; else if (n1166) n1023 <= n6484;
/* FF  5  9  7 */ assign n721 = n6485;
/* FF  4  5  6 */ assign n531 = n6486;
/* FF 11  4  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1414 <= 1'b0; else if (n979) n1414 <= n6487;
/* FF  7 18  5 */ assign n6488 = n6489;
/* FF 17  7  2 */ assign n6490 = n6491;
/* FF  7 10  1 */ always @(posedge io_13_31_1) if (n4) n872 <= 1'b0 ? 1'b0 : n6492;
/* FF  9 21  3 */ assign n1223 = n6493;
/* FF 20 20  1 */ assign n2741 = n6494;
/* FF 14  8  5 */ always @(posedge io_13_31_1) if (n2076) n1748 <= 1'b0 ? 1'b0 : n6495;
/* FF  8  9  4 */ assign n999 = n6496;
/* FF 11 30  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n5 <= 1'b1; else if (1'b1) n5 <= n6497;
/* FF 17  8  3 */ always @(posedge io_13_31_1) if (n2344) n2350 <= 1'b0 ? 1'b0 : n6498;
/* FF 10 18  1 */ assign n6499 = n6500;
/* FF  9 22  4 */ assign n1231 = n6501;
/* FF 23  2  5 */ assign n3007 = n6502;
/* FF  4  6  6 */ assign n540 = n6503;
/* FF 14  1  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1861 <= 1'b0; else if (n1860) n1861 <= n6504;
/* FF  8  2  1 */ assign n941 = n6505;
/* FF 16 12  4 */ assign n2242 = n6506;
/* FF 16  4  0 */ assign n2172 = n6507;
/* FF 13 17  3 */ assign n6508 = n6509;
/* FF 14  4  7 */ assign n1881 = n6510;
/* FF 20 16  3 */ always @(posedge io_13_31_1) if (n2568) n2723 <= 1'b0 ? 1'b0 : n6511;
/* FF  8  1  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n938 <= 1'b0; else if (n656) n938 <= n6512;
/* FF  1 19  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n141 <= 1'b0; else if (n140) n141 <= n6513;
/* FF 18 21  1 */ assign n2583 = n6514;
/* FF  1 11  3 */ assign n42 = n6515;
/* FF 20 15  7 */ assign io_19_31_1 = n6516;
/* FF 17  4  5 */ always @(posedge io_13_31_1) if (n2316) n2330 <= 1'b0 ? 1'b0 : n6517;
/* FF 10 10  2 */ always @(posedge io_13_31_1) if (n4) n1304 <= 1'b0 ? 1'b0 : n6518;
/* FF  9  6  1 */ always @(posedge io_13_31_1) if (n4) n1117 <= 1'b0 ? 1'b0 : n6519;
/* FF 16  5  1 */ assign n1924 = n6520;
/* FF 10 13  7 */ always @(posedge io_13_31_1) if (n4) n1339 <= 1'b0 ? 1'b0 : n6521;
/* FF  3 20  1 */ assign n475 = n6522;
/* FF  9  9  6 */ always @(posedge io_13_31_1) if (n4) n1142 <= 1'b0 ? 1'b0 : n6523;
/* FF  1 12  4 */ assign n86 = n6524;
/* FF  1  4  0 */ always @(posedge io_13_31_1) if (n201) n27 <= n42 ? 1'b0 : n6525;
/* FF 20  8  4 */ assign n2689 = n6526;
/* FF 12 22  5 */ assign n1663 = n6527;
/* FF 18 13  2 */ always @(posedge io_13_31_1) if (n2137) n2530 <= n3 ? 1'b0 : n6528;
/* FF 12 14  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1617 <= 1'b0; else if (n1630) n1617 <= n6529;
/* FF 22 17  1 */ assign n2859 = n6530;
/* FF  2 17  0 */ assign n6531 = n6532;
/* FF 10  6  4 */ always @(posedge io_13_31_1) if (n4) n1269 <= 1'b0 ? 1'b0 : n6534;
/* FF  9 10  7 */ assign n1158 = n6535;
/* FF  9  2  3 */ assign n1086 = n6536;
/* FF 22 20  6 */ assign n2876 = n6537;
/* FF  3 16  3 */ assign n128 = n6538;
/* FF 21 16  5 */ assign n2828 = n6539;
/* FF 20  1  1 */ assign n6540 = n6541;
/* FF  3 15  7 */ assign n443 = n6542;
/* FF 10  7  5 */ always @(posedge io_13_31_1) if (n4) n1276 <= 1'b0 ? 1'b0 : n6543;
/* FF 18  9  4 */ assign n2495 = n6544;
/* FF 22 21  7 */ assign n2882 = n6545;
/* FF 22 13  3 */ always @(posedge io_13_31_1) if (n2663) n2960 <= 1'b0 ? 1'b0 : n6546;
/* FF  4 20  3 */ assign n637 = n6547;
/* FF  2 12  6 */ always @(posedge io_13_31_1, posedge n1) if (n1) n103 <= 1'b0; else if (1'b1) n103 <= n6548;
/* FF 13  5  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1696 <= 1'b0; else if (n1279) n1696 <= n6549;
/* FF  3  8  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n406 <= 1'b0; else if (n71) n406 <= n6550;
/* FF 18 10  5 */ assign n2506 = n6551;
/* FF 18  2  1 */ always @(posedge io_13_31_1) if (n2456) n2444 <= 1'b0 ? 1'b0 : n6552;
/* FF 15 14  2 */ always @(posedge io_13_31_1) if (1'b1) n2125 <= n1970 ? 1'b1 : n6553;
/* FF  5 17  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n769 <= 1'b0; else if (1'b1) n769 <= n6554;
/* FF  4 13  0 */ assign n6555 = n6556;
/* FF  2 13  7 */ assign n268 = n6558;
/* FF 12  2  4 */ assign n1531 = n6559;
/* FF 13  6  6 */ assign n1713 = n6560;
/* FF  2  5  3 */ assign n204 = n6561;
/* FF  3  1  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n339 <= 1'b0; else if (n500) n339 <= n6562;
/* FF  4 16  5 */ assign n249 = n6563;
/* FF 11 11  4 */ assign n1467 = n6564;
/* FF 14 19  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1503 <= 1'b0; else if (n1527) n1503 <= n6565;
/* FF 11  3  0 */ assign n1249 = n6566;
/* FF 14 11  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1556 <= 1'b0; else if (n734) n1556 <= n6567;
/* FF 15 15  3 */ assign n2129 = n6568;
/* FF  3  4  6 */ assign n369 = n6569;
/* FF  7 21  0 */ assign n6570 = n6571;
/* FF 12  3  5 */ assign n6572 = n6573;
/* FF 22  5  3 */ assign n2928 = n6574;
/* FF  5 13  3 */ assign n744 = n6575;
/* FF  4 17  6 */ assign n317 = n6576;
/* FF  4  9  2 */ always @(posedge io_13_31_1) if (n4) n558 <= 1'b0 ? 1'b0 : n6577;
/* FF 17 19  2 */ assign n2420 = n6578;
/* FF 11  7  6 */ assign n1146 = n6579;
/* FF 17 18  6 */ assign n2414 = n6580;
/* FF  7 13  1 */ always @(posedge io_13_31_1) if (n4) n895 <= 1'b0 ? 1'b0 : n6581;
/* FF 14 12  1 */ assign n1942 = n6582;
/* FF  5  5  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n541 <= 1'b0; else if (n524) n541 <= n6583;
/* FF  4  1  3 */ assign n495 = n6584;
/* FF  8 12  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1020 <= 1'b0; else if (n1166) n1020 <= n6585;
/* FF  8  4  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n961 <= 1'b0; else if (n663) n961 <= n6586;
/* FF 16 15  5 */ always @(posedge io_13_31_1) if (n2268) n2262 <= 1'b0 ? 1'b0 : n6587;
/* FF 23 14  5 */ always @(posedge io_13_31_1) if (1'b1) n3023 <= 1'b0 ? 1'b0 : n6588;
/* FF 20 18  2 */ always @(posedge io_13_31_1) if (n2732) n2576 <= 1'b0 ? 1'b0 : n6589;
/* FF 15  3  6 */ assign n1690 = n6590;
/* FF  9 17  0 */ assign n6591 = n6592;
/* FF  7 17  7 */ assign n918 = n6593;
/* FF  7  9  3 */ assign n863 = n6594;
/* FF  8 13  5 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1028 <= 1'b0; else if (n1166) n1028 <= n6595;
/* FF  8  5  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n969 <= 1'b0; else if (n663) n969 <= n6596;
/* FF 14  7  7 */ assign n1912 = n6597;
/* FF 17  7  5 */ always @(posedge io_13_31_1) if (n2191) n2315 <= 1'b0 ? 1'b0 : n6598;
/* FF  3 18  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n461 <= 1'b0; else if (n310) n461 <= n6599;
/* FF  7  2  0 */ assign n829 = n6600;
/* FF  9 21  6 */ assign n1225 = n6601;
/* FF 16  8  1 */ assign n2206 = n6602;
/* FF 13 13  0 */ assign n1770 = n6603;
/* FF  1  7  0 */ assign n6604 = n6605;
/* FF 13 16  5 */ assign n1805 = n6607;
/* FF  3 19  4 */ assign n470 = n6608;
/* FF 12 17  1 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1358 <= 1'b0; else if (1'b1) n1358 <= n6609;
/* FF 20  6  5 */ always @(posedge io_13_31_1) if (n2676) n2681 <= n1 ? 1'b0 : n6610;
/* FF  2 20  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n327 <= 1'b0; else if (1'b1) n327 <= n6611;
/* FF 10  9  4 */ always @(posedge io_13_31_1) if (n4) n1297 <= 1'b0 ? 1'b0 : n6612;
/* FF  9 13  7 */ always @(posedge io_13_31_1) if (n4) n1178 <= 1'b0 ? 1'b0 : n6613;
/* FF  9  5  3 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1110 <= 1'b0; else if (n840) n1110 <= n6614;
/* FF 13 17  6 */ assign n1810 = n6615;
/* FF  1  8  1 */ assign n6616 = n6617;
/* FF 22 23  6 */ always @(posedge io_13_31_1) if (n3004) n3002 <= 1'b0 ? 1'b0 : n6618;
/* FF  1 11  6 */ assign n75 = n6619;
/* FF 12 18  2 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1188 <= 1'b0; else if (1'b1) n1188 <= n6620;
/* FF 20  7  6 */ assign n2622 = n6621;
/* FF 10 10  5 */ assign n1307 = n6622;
/* FF 10  2  1 */ assign n1242 = n6623;
/* FF 12 21  7 */ assign n1658 = n6624;
/* FF  9  6  4 */ assign n806 = n6625;
/* FF 18 12  4 */ always @(posedge io_13_31_1) if (n2137) n2525 <= n3 ? 1'b0 : n6626;
/* FF 18  4  0 */ always @(posedge io_13_31_1) if (n2603) n2450 <= 1'b0 ? 1'b0 : n6627;
/* FF 22 16  3 */ always @(posedge io_13_31_1) if (n2971) n2979 <= 1'b0 ? 1'b0 : n6628;
/* FF 13  9  1 */ assign n1743 = n6629;
/* FF 21 20  6 */ always @(posedge io_13_31_1) if (n2865) n2866 <= 1'b0 ? 1'b0 : n6630;
/* FF 21 12  2 */ always @(posedge io_13_31_1) if (n2663) n2813 <= 1'b0 ? 1'b0 : n6631;
/* FF  3  3  0 */ always @(posedge io_13_31_1, posedge n1) if (n1) n355 <= 1'b0; else if (n198) n355 <= n6632;
/* FF 18 13  5 */ always @(posedge io_13_31_1) if (n2137) n2533 <= n3 ? 1'b0 : n6633;
/* FF  1  3  7 */ always @(posedge io_13_31_1, posedge n1) if (n1) n25 <= 1'b0; else if (n17) n25 <= n6634;
/* FF 18  5  1 */ always @(posedge io_13_31_1) if (n2456) n2458 <= 1'b0 ? 1'b0 : n6635;
/* FF  5 20  1 */ assign n791 = n6636;
/* FF 17 21  2 */ assign n1526 = n6637;
/* FF 12  5  4 */ always @(posedge io_13_31_1, posedge n1) if (n1) n1290 <= 1'b0; else if (n1426) n1290 <= n6638;

endmodule

